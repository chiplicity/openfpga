magic
tech sky130A
magscale 1 2
timestamp 1606929812
<< locali >>
rect 12265 19015 12299 19117
rect 20453 18675 20487 18777
rect 12633 16839 12667 17145
rect 21741 16635 21775 17281
rect 15301 14187 15335 14289
rect 13461 13575 13495 13881
rect 12265 13099 12299 13337
rect 15761 10923 15795 11025
rect 11253 7047 11287 7217
<< viali >>
rect 5089 19865 5123 19899
rect 17877 19865 17911 19899
rect 18613 19865 18647 19899
rect 20729 19865 20763 19899
rect 4997 19729 5031 19763
rect 17693 19729 17727 19763
rect 18429 19729 18463 19763
rect 19533 19729 19567 19763
rect 20545 19729 20579 19763
rect 5181 19661 5215 19695
rect 19809 19661 19843 19695
rect 4629 19525 4663 19559
rect 11069 19321 11103 19355
rect 9689 19185 9723 19219
rect 11897 19185 11931 19219
rect 15853 19185 15887 19219
rect 17233 19185 17267 19219
rect 4077 19117 4111 19151
rect 4344 19117 4378 19151
rect 7757 19117 7791 19151
rect 12265 19117 12299 19151
rect 12357 19117 12391 19151
rect 15761 19117 15795 19151
rect 16957 19117 16991 19151
rect 18153 19117 18187 19151
rect 19533 19117 19567 19151
rect 19809 19117 19843 19151
rect 20269 19117 20303 19151
rect 8024 19049 8058 19083
rect 9956 19049 9990 19083
rect 12624 19049 12658 19083
rect 18797 19049 18831 19083
rect 5457 18981 5491 19015
rect 9137 18981 9171 19015
rect 11345 18981 11379 19015
rect 11713 18981 11747 19015
rect 11805 18981 11839 19015
rect 12265 18981 12299 19015
rect 13737 18981 13771 19015
rect 14013 18981 14047 19015
rect 15301 18981 15335 19015
rect 15669 18981 15703 19015
rect 20453 18981 20487 19015
rect 3801 18777 3835 18811
rect 5273 18777 5307 18811
rect 8217 18777 8251 18811
rect 9689 18777 9723 18811
rect 14841 18777 14875 18811
rect 16773 18777 16807 18811
rect 20453 18777 20487 18811
rect 20729 18777 20763 18811
rect 2688 18709 2722 18743
rect 10968 18709 11002 18743
rect 12909 18709 12943 18743
rect 13728 18709 13762 18743
rect 15384 18709 15418 18743
rect 17233 18709 17267 18743
rect 18337 18709 18371 18743
rect 2421 18641 2455 18675
rect 5181 18641 5215 18675
rect 5825 18641 5859 18675
rect 7104 18641 7138 18675
rect 9597 18641 9631 18675
rect 10701 18641 10735 18675
rect 12817 18641 12851 18675
rect 17141 18641 17175 18675
rect 18061 18641 18095 18675
rect 19533 18641 19567 18675
rect 20453 18641 20487 18675
rect 20545 18641 20579 18675
rect 5457 18573 5491 18607
rect 6837 18573 6871 18607
rect 8493 18573 8527 18607
rect 9781 18573 9815 18607
rect 13001 18573 13035 18607
rect 13461 18573 13495 18607
rect 15117 18573 15151 18607
rect 17325 18573 17359 18607
rect 19717 18573 19751 18607
rect 12081 18505 12115 18539
rect 4813 18437 4847 18471
rect 9229 18437 9263 18471
rect 12449 18437 12483 18471
rect 16497 18437 16531 18471
rect 19717 18233 19751 18267
rect 13369 18165 13403 18199
rect 8033 18097 8067 18131
rect 8861 18097 8895 18131
rect 8953 18097 8987 18131
rect 10793 18097 10827 18131
rect 14013 18097 14047 18131
rect 16589 18097 16623 18131
rect 5273 18029 5307 18063
rect 7757 18029 7791 18063
rect 8769 18029 8803 18063
rect 13829 18029 13863 18063
rect 19533 18029 19567 18063
rect 5549 17961 5583 17995
rect 13737 17961 13771 17995
rect 7389 17893 7423 17927
rect 7849 17893 7883 17927
rect 8401 17893 8435 17927
rect 2881 17689 2915 17723
rect 20453 17689 20487 17723
rect 21005 17689 21039 17723
rect 5264 17621 5298 17655
rect 1501 17553 1535 17587
rect 1768 17553 1802 17587
rect 19717 17553 19751 17587
rect 20269 17553 20303 17587
rect 20821 17553 20855 17587
rect 3341 17485 3375 17519
rect 4997 17485 5031 17519
rect 6377 17349 6411 17383
rect 19901 17349 19935 17383
rect 21741 17281 21775 17315
rect 7941 17145 7975 17179
rect 12633 17145 12667 17179
rect 17877 17145 17911 17179
rect 18153 17145 18187 17179
rect 9781 17077 9815 17111
rect 3525 17009 3559 17043
rect 4537 17009 4571 17043
rect 4629 17009 4663 17043
rect 9137 17009 9171 17043
rect 10425 17009 10459 17043
rect 12357 17009 12391 17043
rect 3341 16941 3375 16975
rect 6561 16941 6595 16975
rect 9045 16941 9079 16975
rect 12265 16941 12299 16975
rect 6828 16873 6862 16907
rect 10241 16873 10275 16907
rect 13369 17009 13403 17043
rect 18705 17009 18739 17043
rect 20269 17009 20303 17043
rect 16497 16941 16531 16975
rect 19257 16941 19291 16975
rect 19993 16941 20027 16975
rect 13277 16873 13311 16907
rect 16764 16873 16798 16907
rect 18613 16873 18647 16907
rect 19533 16873 19567 16907
rect 2973 16805 3007 16839
rect 3433 16805 3467 16839
rect 4077 16805 4111 16839
rect 4445 16805 4479 16839
rect 8585 16805 8619 16839
rect 8953 16805 8987 16839
rect 10149 16805 10183 16839
rect 11805 16805 11839 16839
rect 12173 16805 12207 16839
rect 12633 16805 12667 16839
rect 12817 16805 12851 16839
rect 13185 16805 13219 16839
rect 18521 16805 18555 16839
rect 6929 16601 6963 16635
rect 10149 16601 10183 16635
rect 11805 16601 11839 16635
rect 16957 16601 16991 16635
rect 18061 16601 18095 16635
rect 20729 16601 20763 16635
rect 21741 16601 21775 16635
rect 9036 16533 9070 16567
rect 10670 16533 10704 16567
rect 15844 16533 15878 16567
rect 18981 16533 19015 16567
rect 19717 16533 19751 16567
rect 3893 16465 3927 16499
rect 7297 16465 7331 16499
rect 7941 16465 7975 16499
rect 8769 16465 8803 16499
rect 13257 16465 13291 16499
rect 15025 16465 15059 16499
rect 18705 16465 18739 16499
rect 19441 16465 19475 16499
rect 20545 16465 20579 16499
rect 4169 16397 4203 16431
rect 7389 16397 7423 16431
rect 7481 16397 7515 16431
rect 10425 16397 10459 16431
rect 13001 16397 13035 16431
rect 15577 16397 15611 16431
rect 14381 16261 14415 16295
rect 3157 16057 3191 16091
rect 7113 16057 7147 16091
rect 7389 16057 7423 16091
rect 12909 16057 12943 16091
rect 16589 16057 16623 16091
rect 20453 16057 20487 16091
rect 1777 15921 1811 15955
rect 7849 15921 7883 15955
rect 7941 15921 7975 15955
rect 10149 15921 10183 15955
rect 13185 15921 13219 15955
rect 14657 15921 14691 15955
rect 15853 15921 15887 15955
rect 17141 15921 17175 15955
rect 5733 15853 5767 15887
rect 6000 15853 6034 15887
rect 11529 15853 11563 15887
rect 11796 15853 11830 15887
rect 14565 15853 14599 15887
rect 15669 15853 15703 15887
rect 17049 15853 17083 15887
rect 18889 15853 18923 15887
rect 20269 15853 20303 15887
rect 2044 15785 2078 15819
rect 15761 15785 15795 15819
rect 19165 15785 19199 15819
rect 7757 15717 7791 15751
rect 14105 15717 14139 15751
rect 14473 15717 14507 15751
rect 15301 15717 15335 15751
rect 16957 15717 16991 15751
rect 2973 15513 3007 15547
rect 3249 15513 3283 15547
rect 6193 15513 6227 15547
rect 20177 15513 20211 15547
rect 20729 15513 20763 15547
rect 1593 15377 1627 15411
rect 1860 15377 1894 15411
rect 3617 15377 3651 15411
rect 4261 15377 4295 15411
rect 5080 15377 5114 15411
rect 7389 15377 7423 15411
rect 18981 15377 19015 15411
rect 19993 15377 20027 15411
rect 20545 15377 20579 15411
rect 3709 15309 3743 15343
rect 3801 15309 3835 15343
rect 4813 15309 4847 15343
rect 19257 15309 19291 15343
rect 7205 15173 7239 15207
rect 4077 14969 4111 15003
rect 9689 14969 9723 15003
rect 19901 14969 19935 15003
rect 20453 14969 20487 15003
rect 8033 14901 8067 14935
rect 13185 14901 13219 14935
rect 14933 14901 14967 14935
rect 4629 14833 4663 14867
rect 8493 14833 8527 14867
rect 8677 14833 8711 14867
rect 10149 14833 10183 14867
rect 10241 14833 10275 14867
rect 12449 14833 12483 14867
rect 12541 14833 12575 14867
rect 13553 14833 13587 14867
rect 17049 14833 17083 14867
rect 19073 14833 19107 14867
rect 4537 14765 4571 14799
rect 13369 14765 13403 14799
rect 13820 14765 13854 14799
rect 18797 14765 18831 14799
rect 19717 14765 19751 14799
rect 20269 14765 20303 14799
rect 4445 14697 4479 14731
rect 10057 14697 10091 14731
rect 10701 14697 10735 14731
rect 16865 14697 16899 14731
rect 8401 14629 8435 14663
rect 11989 14629 12023 14663
rect 12357 14629 12391 14663
rect 16497 14629 16531 14663
rect 16957 14629 16991 14663
rect 9781 14425 9815 14459
rect 12909 14425 12943 14459
rect 16865 14425 16899 14459
rect 20913 14425 20947 14459
rect 4160 14357 4194 14391
rect 14096 14357 14130 14391
rect 19533 14357 19567 14391
rect 3893 14289 3927 14323
rect 6101 14289 6135 14323
rect 8668 14289 8702 14323
rect 12817 14289 12851 14323
rect 13829 14289 13863 14323
rect 15301 14289 15335 14323
rect 15752 14289 15786 14323
rect 19257 14289 19291 14323
rect 19993 14289 20027 14323
rect 20729 14289 20763 14323
rect 6193 14221 6227 14255
rect 6285 14221 6319 14255
rect 8401 14221 8435 14255
rect 13001 14221 13035 14255
rect 15485 14221 15519 14255
rect 17325 14221 17359 14255
rect 20177 14221 20211 14255
rect 15209 14153 15243 14187
rect 15301 14153 15335 14187
rect 5273 14085 5307 14119
rect 5733 14085 5767 14119
rect 12449 14085 12483 14119
rect 6285 13881 6319 13915
rect 8677 13881 8711 13915
rect 8953 13881 8987 13915
rect 12357 13881 12391 13915
rect 12633 13881 12667 13915
rect 13461 13881 13495 13915
rect 17417 13881 17451 13915
rect 18613 13881 18647 13915
rect 20453 13881 20487 13915
rect 3617 13813 3651 13847
rect 6561 13745 6595 13779
rect 13185 13745 13219 13779
rect 2237 13677 2271 13711
rect 4905 13677 4939 13711
rect 5172 13677 5206 13711
rect 7297 13677 7331 13711
rect 7564 13677 7598 13711
rect 9137 13677 9171 13711
rect 10977 13677 11011 13711
rect 2504 13609 2538 13643
rect 11222 13609 11256 13643
rect 13001 13609 13035 13643
rect 16405 13813 16439 13847
rect 16865 13745 16899 13779
rect 17049 13745 17083 13779
rect 17969 13745 18003 13779
rect 17877 13677 17911 13711
rect 18429 13677 18463 13711
rect 20269 13677 20303 13711
rect 13645 13609 13679 13643
rect 17785 13609 17819 13643
rect 13093 13541 13127 13575
rect 13461 13541 13495 13575
rect 16773 13541 16807 13575
rect 5641 13337 5675 13371
rect 11345 13337 11379 13371
rect 12265 13337 12299 13371
rect 19625 13337 19659 13371
rect 20177 13337 20211 13371
rect 20729 13337 20763 13371
rect 6101 13269 6135 13303
rect 10059 13269 10093 13303
rect 6009 13201 6043 13235
rect 6285 13133 6319 13167
rect 18981 13269 19015 13303
rect 18705 13201 18739 13235
rect 19441 13201 19475 13235
rect 19993 13201 20027 13235
rect 20545 13201 20579 13235
rect 12265 13065 12299 13099
rect 7573 12793 7607 12827
rect 11345 12793 11379 12827
rect 12449 12793 12483 12827
rect 20177 12793 20211 12827
rect 13001 12725 13035 12759
rect 9965 12657 9999 12691
rect 11713 12657 11747 12691
rect 13461 12657 13495 12691
rect 13645 12657 13679 12691
rect 14657 12657 14691 12691
rect 16589 12657 16623 12691
rect 7757 12589 7791 12623
rect 11437 12589 11471 12623
rect 12641 12589 12675 12623
rect 15301 12589 15335 12623
rect 15577 12589 15611 12623
rect 19165 12589 19199 12623
rect 19441 12589 19475 12623
rect 19993 12589 20027 12623
rect 10232 12521 10266 12555
rect 14473 12521 14507 12555
rect 16856 12521 16890 12555
rect 13369 12453 13403 12487
rect 14013 12453 14047 12487
rect 14381 12453 14415 12487
rect 17969 12453 18003 12487
rect 10425 12249 10459 12283
rect 14565 12249 14599 12283
rect 16589 12249 16623 12283
rect 18061 12249 18095 12283
rect 20177 12249 20211 12283
rect 12716 12181 12750 12215
rect 14473 12181 14507 12215
rect 15476 12181 15510 12215
rect 7021 12113 7055 12147
rect 7288 12113 7322 12147
rect 8769 12113 8803 12147
rect 9025 12113 9059 12147
rect 10793 12113 10827 12147
rect 15209 12113 15243 12147
rect 18429 12113 18463 12147
rect 19993 12113 20027 12147
rect 20545 12113 20579 12147
rect 10885 12045 10919 12079
rect 10977 12045 11011 12079
rect 12449 12045 12483 12079
rect 14657 12045 14691 12079
rect 18521 12045 18555 12079
rect 18613 12045 18647 12079
rect 10149 11977 10183 12011
rect 13829 11977 13863 12011
rect 20729 11977 20763 12011
rect 8401 11909 8435 11943
rect 14105 11909 14139 11943
rect 8033 11705 8067 11739
rect 10425 11705 10459 11739
rect 13277 11705 13311 11739
rect 13553 11705 13587 11739
rect 18061 11705 18095 11739
rect 20453 11705 20487 11739
rect 7205 11569 7239 11603
rect 7297 11569 7331 11603
rect 8677 11569 8711 11603
rect 10885 11569 10919 11603
rect 10977 11569 11011 11603
rect 14013 11569 14047 11603
rect 14105 11569 14139 11603
rect 18613 11569 18647 11603
rect 7113 11501 7147 11535
rect 13461 11501 13495 11535
rect 20269 11501 20303 11535
rect 8493 11433 8527 11467
rect 10793 11433 10827 11467
rect 11437 11433 11471 11467
rect 18429 11433 18463 11467
rect 19073 11433 19107 11467
rect 6745 11365 6779 11399
rect 8401 11365 8435 11399
rect 13921 11365 13955 11399
rect 18521 11365 18555 11399
rect 8309 11161 8343 11195
rect 8769 11161 8803 11195
rect 13737 11161 13771 11195
rect 15945 11161 15979 11195
rect 17417 11161 17451 11195
rect 18797 11161 18831 11195
rect 20177 11161 20211 11195
rect 20729 11161 20763 11195
rect 8677 11093 8711 11127
rect 10977 11093 11011 11127
rect 10701 11025 10735 11059
rect 14105 11025 14139 11059
rect 14749 11025 14783 11059
rect 15761 11025 15795 11059
rect 16313 11025 16347 11059
rect 17325 11025 17359 11059
rect 19165 11025 19199 11059
rect 19993 11025 20027 11059
rect 20545 11025 20579 11059
rect 8861 10957 8895 10991
rect 14197 10957 14231 10991
rect 14289 10957 14323 10991
rect 16405 10957 16439 10991
rect 16589 10957 16623 10991
rect 17509 10957 17543 10991
rect 19257 10957 19291 10991
rect 19349 10957 19383 10991
rect 15761 10889 15795 10923
rect 16957 10889 16991 10923
rect 14105 10617 14139 10651
rect 16589 10617 16623 10651
rect 18429 10617 18463 10651
rect 20453 10617 20487 10651
rect 8585 10549 8619 10583
rect 11529 10481 11563 10515
rect 11713 10481 11747 10515
rect 12725 10481 12759 10515
rect 17233 10481 17267 10515
rect 19073 10481 19107 10515
rect 7205 10413 7239 10447
rect 11437 10413 11471 10447
rect 12992 10413 13026 10447
rect 16957 10413 16991 10447
rect 20269 10413 20303 10447
rect 7472 10345 7506 10379
rect 18797 10345 18831 10379
rect 11069 10277 11103 10311
rect 17049 10277 17083 10311
rect 18889 10277 18923 10311
rect 10057 10073 10091 10107
rect 10425 10073 10459 10107
rect 11069 10073 11103 10107
rect 17325 10073 17359 10107
rect 19901 10073 19935 10107
rect 20729 10073 20763 10107
rect 11437 10005 11471 10039
rect 16212 10005 16246 10039
rect 11529 9937 11563 9971
rect 15945 9937 15979 9971
rect 18788 9937 18822 9971
rect 20545 9937 20579 9971
rect 10517 9869 10551 9903
rect 10609 9869 10643 9903
rect 11621 9869 11655 9903
rect 18521 9869 18555 9903
rect 10517 9529 10551 9563
rect 12357 9529 12391 9563
rect 18705 9529 18739 9563
rect 9321 9461 9355 9495
rect 14933 9461 14967 9495
rect 15485 9461 15519 9495
rect 11161 9393 11195 9427
rect 11529 9393 11563 9427
rect 13001 9393 13035 9427
rect 13553 9393 13587 9427
rect 19257 9393 19291 9427
rect 19717 9393 19751 9427
rect 7941 9325 7975 9359
rect 8208 9325 8242 9359
rect 13820 9325 13854 9359
rect 15301 9325 15335 9359
rect 19073 9325 19107 9359
rect 10977 9257 11011 9291
rect 12725 9257 12759 9291
rect 10885 9189 10919 9223
rect 12817 9189 12851 9223
rect 19165 9189 19199 9223
rect 10977 8985 11011 9019
rect 11437 8985 11471 9019
rect 13461 8985 13495 9019
rect 19717 8985 19751 9019
rect 20177 8985 20211 9019
rect 20729 8985 20763 9019
rect 11345 8917 11379 8951
rect 15761 8917 15795 8951
rect 8484 8849 8518 8883
rect 13277 8849 13311 8883
rect 15485 8849 15519 8883
rect 18604 8849 18638 8883
rect 19993 8849 20027 8883
rect 20545 8849 20579 8883
rect 8217 8781 8251 8815
rect 11529 8781 11563 8815
rect 18337 8781 18371 8815
rect 9597 8713 9631 8747
rect 11529 8441 11563 8475
rect 16313 8441 16347 8475
rect 20453 8441 20487 8475
rect 13553 8305 13587 8339
rect 16957 8305 16991 8339
rect 11345 8237 11379 8271
rect 13369 8237 13403 8271
rect 20269 8237 20303 8271
rect 16681 8169 16715 8203
rect 17325 8169 17359 8203
rect 10701 8101 10735 8135
rect 16773 8101 16807 8135
rect 10793 7897 10827 7931
rect 13737 7897 13771 7931
rect 17693 7897 17727 7931
rect 19441 7897 19475 7931
rect 11713 7829 11747 7863
rect 16580 7829 16614 7863
rect 18306 7829 18340 7863
rect 11437 7761 11471 7795
rect 14105 7761 14139 7795
rect 16313 7761 16347 7795
rect 19993 7761 20027 7795
rect 20545 7761 20579 7795
rect 10885 7693 10919 7727
rect 11069 7693 11103 7727
rect 14197 7693 14231 7727
rect 14381 7693 14415 7727
rect 18061 7693 18095 7727
rect 10425 7625 10459 7659
rect 20729 7625 20763 7659
rect 20177 7557 20211 7591
rect 11069 7353 11103 7387
rect 16681 7353 16715 7387
rect 16957 7353 16991 7387
rect 14381 7285 14415 7319
rect 11253 7217 11287 7251
rect 11345 7217 11379 7251
rect 14657 7217 14691 7251
rect 17509 7217 17543 7251
rect 9689 7149 9723 7183
rect 9934 7081 9968 7115
rect 13001 7149 13035 7183
rect 13268 7149 13302 7183
rect 15301 7149 15335 7183
rect 17417 7149 17451 7183
rect 11590 7081 11624 7115
rect 15546 7081 15580 7115
rect 17325 7081 17359 7115
rect 11253 7013 11287 7047
rect 12725 7013 12759 7047
rect 10609 6809 10643 6843
rect 14105 6809 14139 6843
rect 10977 6741 11011 6775
rect 14473 6741 14507 6775
rect 7645 6673 7679 6707
rect 11069 6673 11103 6707
rect 14565 6673 14599 6707
rect 20545 6673 20579 6707
rect 7389 6605 7423 6639
rect 11161 6605 11195 6639
rect 14657 6605 14691 6639
rect 8769 6537 8803 6571
rect 20729 6537 20763 6571
rect 20729 5721 20763 5755
rect 20545 5585 20579 5619
rect 20729 4633 20763 4667
rect 20545 4497 20579 4531
<< metal1 >>
rect 1104 20010 21620 20032
rect 1104 19958 7846 20010
rect 7898 19958 7910 20010
rect 7962 19958 7974 20010
rect 8026 19958 8038 20010
rect 8090 19958 14710 20010
rect 14762 19958 14774 20010
rect 14826 19958 14838 20010
rect 14890 19958 14902 20010
rect 14954 19958 21620 20010
rect 1104 19936 21620 19958
rect 4706 19856 4712 19908
rect 4764 19896 4770 19908
rect 5077 19899 5135 19905
rect 5077 19896 5089 19899
rect 4764 19868 5089 19896
rect 4764 19856 4770 19868
rect 5077 19865 5089 19868
rect 5123 19865 5135 19899
rect 5077 19859 5135 19865
rect 17865 19899 17923 19905
rect 17865 19865 17877 19899
rect 17911 19896 17923 19899
rect 17954 19896 17960 19908
rect 17911 19868 17960 19896
rect 17911 19865 17923 19868
rect 17865 19859 17923 19865
rect 17954 19856 17960 19868
rect 18012 19856 18018 19908
rect 18601 19899 18659 19905
rect 18601 19865 18613 19899
rect 18647 19896 18659 19899
rect 18690 19896 18696 19908
rect 18647 19868 18696 19896
rect 18647 19865 18659 19868
rect 18601 19859 18659 19865
rect 18690 19856 18696 19868
rect 18748 19856 18754 19908
rect 20622 19856 20628 19908
rect 20680 19896 20686 19908
rect 20717 19899 20775 19905
rect 20717 19896 20729 19899
rect 20680 19868 20729 19896
rect 20680 19856 20686 19868
rect 20717 19865 20729 19868
rect 20763 19865 20775 19899
rect 20717 19859 20775 19865
rect 4985 19763 5043 19769
rect 4985 19729 4997 19763
rect 5031 19760 5043 19763
rect 9582 19760 9588 19772
rect 5031 19732 9588 19760
rect 5031 19729 5043 19732
rect 4985 19723 5043 19729
rect 9582 19720 9588 19732
rect 9640 19720 9646 19772
rect 17678 19760 17684 19772
rect 17639 19732 17684 19760
rect 17678 19720 17684 19732
rect 17736 19720 17742 19772
rect 18417 19763 18475 19769
rect 18417 19729 18429 19763
rect 18463 19760 18475 19763
rect 18506 19760 18512 19772
rect 18463 19732 18512 19760
rect 18463 19729 18475 19732
rect 18417 19723 18475 19729
rect 18506 19720 18512 19732
rect 18564 19720 18570 19772
rect 19426 19720 19432 19772
rect 19484 19760 19490 19772
rect 19521 19763 19579 19769
rect 19521 19760 19533 19763
rect 19484 19732 19533 19760
rect 19484 19720 19490 19732
rect 19521 19729 19533 19732
rect 19567 19729 19579 19763
rect 19521 19723 19579 19729
rect 19702 19720 19708 19772
rect 19760 19760 19766 19772
rect 20533 19763 20591 19769
rect 20533 19760 20545 19763
rect 19760 19732 20545 19760
rect 19760 19720 19766 19732
rect 20533 19729 20545 19732
rect 20579 19729 20591 19763
rect 20533 19723 20591 19729
rect 5166 19692 5172 19704
rect 5127 19664 5172 19692
rect 5166 19652 5172 19664
rect 5224 19652 5230 19704
rect 19794 19692 19800 19704
rect 19755 19664 19800 19692
rect 19794 19652 19800 19664
rect 19852 19652 19858 19704
rect 4617 19559 4675 19565
rect 4617 19525 4629 19559
rect 4663 19556 4675 19559
rect 5258 19556 5264 19568
rect 4663 19528 5264 19556
rect 4663 19525 4675 19528
rect 4617 19519 4675 19525
rect 5258 19516 5264 19528
rect 5316 19516 5322 19568
rect 1104 19466 21620 19488
rect 1104 19414 4414 19466
rect 4466 19414 4478 19466
rect 4530 19414 4542 19466
rect 4594 19414 4606 19466
rect 4658 19414 11278 19466
rect 11330 19414 11342 19466
rect 11394 19414 11406 19466
rect 11458 19414 11470 19466
rect 11522 19414 18142 19466
rect 18194 19414 18206 19466
rect 18258 19414 18270 19466
rect 18322 19414 18334 19466
rect 18386 19414 21620 19466
rect 1104 19392 21620 19414
rect 11054 19352 11060 19364
rect 10967 19324 11060 19352
rect 11054 19312 11060 19324
rect 11112 19352 11118 19364
rect 11112 19324 11928 19352
rect 11112 19312 11118 19324
rect 11900 19225 11928 19324
rect 9677 19219 9735 19225
rect 9677 19185 9689 19219
rect 9723 19185 9735 19219
rect 9677 19179 9735 19185
rect 11885 19219 11943 19225
rect 11885 19185 11897 19219
rect 11931 19185 11943 19219
rect 11885 19179 11943 19185
rect 2406 19108 2412 19160
rect 2464 19148 2470 19160
rect 4338 19157 4344 19160
rect 4065 19151 4123 19157
rect 4065 19148 4077 19151
rect 2464 19120 4077 19148
rect 2464 19108 2470 19120
rect 4065 19117 4077 19120
rect 4111 19117 4123 19151
rect 4332 19148 4344 19157
rect 4251 19120 4344 19148
rect 4065 19111 4123 19117
rect 4332 19111 4344 19120
rect 4396 19148 4402 19160
rect 5166 19148 5172 19160
rect 4396 19120 5172 19148
rect 4338 19108 4344 19111
rect 4396 19108 4402 19120
rect 5166 19108 5172 19120
rect 5224 19108 5230 19160
rect 6546 19108 6552 19160
rect 6604 19148 6610 19160
rect 7745 19151 7803 19157
rect 7745 19148 7757 19151
rect 6604 19120 7757 19148
rect 6604 19108 6610 19120
rect 7745 19117 7757 19120
rect 7791 19117 7803 19151
rect 7745 19111 7803 19117
rect 7944 19120 9536 19148
rect 1946 19040 1952 19092
rect 2004 19080 2010 19092
rect 2004 19052 5580 19080
rect 2004 19040 2010 19052
rect 5442 19012 5448 19024
rect 5403 18984 5448 19012
rect 5442 18972 5448 18984
rect 5500 18972 5506 19024
rect 5552 19012 5580 19052
rect 5810 19040 5816 19092
rect 5868 19080 5874 19092
rect 7944 19080 7972 19120
rect 5868 19052 7972 19080
rect 8012 19083 8070 19089
rect 5868 19040 5874 19052
rect 8012 19049 8024 19083
rect 8058 19080 8070 19083
rect 8202 19080 8208 19092
rect 8058 19052 8208 19080
rect 8058 19049 8070 19052
rect 8012 19043 8070 19049
rect 8202 19040 8208 19052
rect 8260 19040 8266 19092
rect 9508 19080 9536 19120
rect 9692 19080 9720 19179
rect 15378 19176 15384 19228
rect 15436 19216 15442 19228
rect 15841 19219 15899 19225
rect 15841 19216 15853 19219
rect 15436 19188 15853 19216
rect 15436 19176 15442 19188
rect 15841 19185 15853 19188
rect 15887 19185 15899 19219
rect 15841 19179 15899 19185
rect 17221 19219 17279 19225
rect 17221 19185 17233 19219
rect 17267 19216 17279 19219
rect 17678 19216 17684 19228
rect 17267 19188 17684 19216
rect 17267 19185 17279 19188
rect 17221 19179 17279 19185
rect 17678 19176 17684 19188
rect 17736 19176 17742 19228
rect 12253 19151 12311 19157
rect 12253 19117 12265 19151
rect 12299 19148 12311 19151
rect 12345 19151 12403 19157
rect 12345 19148 12357 19151
rect 12299 19120 12357 19148
rect 12299 19117 12311 19120
rect 12253 19111 12311 19117
rect 12345 19117 12357 19120
rect 12391 19117 12403 19151
rect 15749 19151 15807 19157
rect 15749 19148 15761 19151
rect 12345 19111 12403 19117
rect 12544 19120 15761 19148
rect 9766 19080 9772 19092
rect 9508 19052 9628 19080
rect 9692 19052 9772 19080
rect 6730 19012 6736 19024
rect 5552 18984 6736 19012
rect 6730 18972 6736 18984
rect 6788 18972 6794 19024
rect 6822 18972 6828 19024
rect 6880 19012 6886 19024
rect 9030 19012 9036 19024
rect 6880 18984 9036 19012
rect 6880 18972 6886 18984
rect 9030 18972 9036 18984
rect 9088 18972 9094 19024
rect 9125 19015 9183 19021
rect 9125 18981 9137 19015
rect 9171 19012 9183 19015
rect 9490 19012 9496 19024
rect 9171 18984 9496 19012
rect 9171 18981 9183 18984
rect 9125 18975 9183 18981
rect 9490 18972 9496 18984
rect 9548 18972 9554 19024
rect 9600 19012 9628 19052
rect 9766 19040 9772 19052
rect 9824 19040 9830 19092
rect 9950 19089 9956 19092
rect 9944 19080 9956 19089
rect 9911 19052 9956 19080
rect 9944 19043 9956 19052
rect 9950 19040 9956 19043
rect 10008 19040 10014 19092
rect 10226 19040 10232 19092
rect 10284 19080 10290 19092
rect 12544 19080 12572 19120
rect 15749 19117 15761 19120
rect 15795 19117 15807 19151
rect 15749 19111 15807 19117
rect 16758 19108 16764 19160
rect 16816 19148 16822 19160
rect 16945 19151 17003 19157
rect 16945 19148 16957 19151
rect 16816 19120 16957 19148
rect 16816 19108 16822 19120
rect 16945 19117 16957 19120
rect 16991 19117 17003 19151
rect 16945 19111 17003 19117
rect 18141 19151 18199 19157
rect 18141 19117 18153 19151
rect 18187 19148 18199 19151
rect 18874 19148 18880 19160
rect 18187 19120 18880 19148
rect 18187 19117 18199 19120
rect 18141 19111 18199 19117
rect 18874 19108 18880 19120
rect 18932 19108 18938 19160
rect 19518 19148 19524 19160
rect 19479 19120 19524 19148
rect 19518 19108 19524 19120
rect 19576 19108 19582 19160
rect 19797 19151 19855 19157
rect 19797 19117 19809 19151
rect 19843 19148 19855 19151
rect 20257 19151 20315 19157
rect 20257 19148 20269 19151
rect 19843 19120 20269 19148
rect 19843 19117 19855 19120
rect 19797 19111 19855 19117
rect 20257 19117 20269 19120
rect 20303 19117 20315 19151
rect 20257 19111 20315 19117
rect 12618 19089 12624 19092
rect 10284 19052 12572 19080
rect 10284 19040 10290 19052
rect 12612 19043 12624 19089
rect 12676 19080 12682 19092
rect 18782 19080 18788 19092
rect 12676 19052 12712 19080
rect 18743 19052 18788 19080
rect 12618 19040 12624 19043
rect 12676 19040 12682 19052
rect 18782 19040 18788 19052
rect 18840 19040 18846 19092
rect 19610 19080 19616 19092
rect 19168 19052 19616 19080
rect 10962 19012 10968 19024
rect 9600 18984 10968 19012
rect 10962 18972 10968 18984
rect 11020 18972 11026 19024
rect 11146 18972 11152 19024
rect 11204 19012 11210 19024
rect 11333 19015 11391 19021
rect 11333 19012 11345 19015
rect 11204 18984 11345 19012
rect 11204 18972 11210 18984
rect 11333 18981 11345 18984
rect 11379 18981 11391 19015
rect 11698 19012 11704 19024
rect 11659 18984 11704 19012
rect 11333 18975 11391 18981
rect 11698 18972 11704 18984
rect 11756 18972 11762 19024
rect 11790 18972 11796 19024
rect 11848 19012 11854 19024
rect 12253 19015 12311 19021
rect 11848 18984 11893 19012
rect 11848 18972 11854 18984
rect 12253 18981 12265 19015
rect 12299 19012 12311 19015
rect 12710 19012 12716 19024
rect 12299 18984 12716 19012
rect 12299 18981 12311 18984
rect 12253 18975 12311 18981
rect 12710 18972 12716 18984
rect 12768 19012 12774 19024
rect 13446 19012 13452 19024
rect 12768 18984 13452 19012
rect 12768 18972 12774 18984
rect 13446 18972 13452 18984
rect 13504 18972 13510 19024
rect 13722 19012 13728 19024
rect 13683 18984 13728 19012
rect 13722 18972 13728 18984
rect 13780 18972 13786 19024
rect 13998 19012 14004 19024
rect 13959 18984 14004 19012
rect 13998 18972 14004 18984
rect 14056 18972 14062 19024
rect 15289 19015 15347 19021
rect 15289 18981 15301 19015
rect 15335 19012 15347 19015
rect 15562 19012 15568 19024
rect 15335 18984 15568 19012
rect 15335 18981 15347 18984
rect 15289 18975 15347 18981
rect 15562 18972 15568 18984
rect 15620 18972 15626 19024
rect 15657 19015 15715 19021
rect 15657 18981 15669 19015
rect 15703 19012 15715 19015
rect 15746 19012 15752 19024
rect 15703 18984 15752 19012
rect 15703 18981 15715 18984
rect 15657 18975 15715 18981
rect 15746 18972 15752 18984
rect 15804 18972 15810 19024
rect 15838 18972 15844 19024
rect 15896 19012 15902 19024
rect 19168 19012 19196 19052
rect 19610 19040 19616 19052
rect 19668 19040 19674 19092
rect 15896 18984 19196 19012
rect 15896 18972 15902 18984
rect 19242 18972 19248 19024
rect 19300 19012 19306 19024
rect 20441 19015 20499 19021
rect 20441 19012 20453 19015
rect 19300 18984 20453 19012
rect 19300 18972 19306 18984
rect 20441 18981 20453 18984
rect 20487 18981 20499 19015
rect 20441 18975 20499 18981
rect 1104 18922 21620 18944
rect 1104 18870 7846 18922
rect 7898 18870 7910 18922
rect 7962 18870 7974 18922
rect 8026 18870 8038 18922
rect 8090 18870 14710 18922
rect 14762 18870 14774 18922
rect 14826 18870 14838 18922
rect 14890 18870 14902 18922
rect 14954 18870 21620 18922
rect 1104 18848 21620 18870
rect 2498 18768 2504 18820
rect 2556 18808 2562 18820
rect 3789 18811 3847 18817
rect 2556 18780 3740 18808
rect 2556 18768 2562 18780
rect 2676 18743 2734 18749
rect 2676 18709 2688 18743
rect 2722 18740 2734 18743
rect 2866 18740 2872 18752
rect 2722 18712 2872 18740
rect 2722 18709 2734 18712
rect 2676 18703 2734 18709
rect 2866 18700 2872 18712
rect 2924 18700 2930 18752
rect 3712 18740 3740 18780
rect 3789 18777 3801 18811
rect 3835 18808 3847 18811
rect 4338 18808 4344 18820
rect 3835 18780 4344 18808
rect 3835 18777 3847 18780
rect 3789 18771 3847 18777
rect 4338 18768 4344 18780
rect 4396 18768 4402 18820
rect 5258 18808 5264 18820
rect 5219 18780 5264 18808
rect 5258 18768 5264 18780
rect 5316 18768 5322 18820
rect 8202 18808 8208 18820
rect 5368 18780 7788 18808
rect 8163 18780 8208 18808
rect 5368 18740 5396 18780
rect 3712 18712 5396 18740
rect 2406 18672 2412 18684
rect 2367 18644 2412 18672
rect 2406 18632 2412 18644
rect 2464 18632 2470 18684
rect 5169 18675 5227 18681
rect 5169 18641 5181 18675
rect 5215 18672 5227 18675
rect 5813 18675 5871 18681
rect 5813 18672 5825 18675
rect 5215 18644 5825 18672
rect 5215 18641 5227 18644
rect 5169 18635 5227 18641
rect 5813 18641 5825 18644
rect 5859 18641 5871 18675
rect 5813 18635 5871 18641
rect 7092 18675 7150 18681
rect 7092 18641 7104 18675
rect 7138 18672 7150 18675
rect 7650 18672 7656 18684
rect 7138 18644 7656 18672
rect 7138 18641 7150 18644
rect 7092 18635 7150 18641
rect 7650 18632 7656 18644
rect 7708 18632 7714 18684
rect 7760 18672 7788 18780
rect 8202 18768 8208 18780
rect 8260 18768 8266 18820
rect 9122 18768 9128 18820
rect 9180 18808 9186 18820
rect 9677 18811 9735 18817
rect 9677 18808 9689 18811
rect 9180 18780 9689 18808
rect 9180 18768 9186 18780
rect 9677 18777 9689 18780
rect 9723 18777 9735 18811
rect 9677 18771 9735 18777
rect 9858 18768 9864 18820
rect 9916 18808 9922 18820
rect 14090 18808 14096 18820
rect 9916 18780 11192 18808
rect 9916 18768 9922 18780
rect 10956 18743 11014 18749
rect 10956 18709 10968 18743
rect 11002 18740 11014 18743
rect 11054 18740 11060 18752
rect 11002 18712 11060 18740
rect 11002 18709 11014 18712
rect 10956 18703 11014 18709
rect 11054 18700 11060 18712
rect 11112 18700 11118 18752
rect 11164 18740 11192 18780
rect 13740 18780 14096 18808
rect 13740 18752 13768 18780
rect 14090 18768 14096 18780
rect 14148 18768 14154 18820
rect 14829 18811 14887 18817
rect 14829 18777 14841 18811
rect 14875 18777 14887 18811
rect 16758 18808 16764 18820
rect 16719 18780 16764 18808
rect 14829 18771 14887 18777
rect 13722 18749 13728 18752
rect 12897 18743 12955 18749
rect 12897 18740 12909 18743
rect 11164 18712 12909 18740
rect 12897 18709 12909 18712
rect 12943 18709 12955 18743
rect 13716 18740 13728 18749
rect 13683 18712 13728 18740
rect 12897 18703 12955 18709
rect 13716 18703 13728 18712
rect 13722 18700 13728 18703
rect 13780 18700 13786 18752
rect 13906 18700 13912 18752
rect 13964 18740 13970 18752
rect 14550 18740 14556 18752
rect 13964 18712 14556 18740
rect 13964 18700 13970 18712
rect 14550 18700 14556 18712
rect 14608 18700 14614 18752
rect 14844 18740 14872 18771
rect 16758 18768 16764 18780
rect 16816 18768 16822 18820
rect 16942 18768 16948 18820
rect 17000 18808 17006 18820
rect 17000 18780 17908 18808
rect 17000 18768 17006 18780
rect 15378 18749 15384 18752
rect 15372 18740 15384 18749
rect 14844 18712 15384 18740
rect 15372 18703 15384 18712
rect 15378 18700 15384 18703
rect 15436 18700 15442 18752
rect 15562 18700 15568 18752
rect 15620 18740 15626 18752
rect 17221 18743 17279 18749
rect 17221 18740 17233 18743
rect 15620 18712 17233 18740
rect 15620 18700 15626 18712
rect 17221 18709 17233 18712
rect 17267 18709 17279 18743
rect 17880 18740 17908 18780
rect 17954 18768 17960 18820
rect 18012 18808 18018 18820
rect 19334 18808 19340 18820
rect 18012 18780 19340 18808
rect 18012 18768 18018 18780
rect 19334 18768 19340 18780
rect 19392 18768 19398 18820
rect 19794 18768 19800 18820
rect 19852 18808 19858 18820
rect 20441 18811 20499 18817
rect 20441 18808 20453 18811
rect 19852 18780 20453 18808
rect 19852 18768 19858 18780
rect 20441 18777 20453 18780
rect 20487 18777 20499 18811
rect 20714 18808 20720 18820
rect 20675 18780 20720 18808
rect 20441 18771 20499 18777
rect 20714 18768 20720 18780
rect 20772 18768 20778 18820
rect 18325 18743 18383 18749
rect 17880 18712 18276 18740
rect 17221 18703 17279 18709
rect 8846 18672 8852 18684
rect 7760 18644 8852 18672
rect 8846 18632 8852 18644
rect 8904 18632 8910 18684
rect 9582 18672 9588 18684
rect 9543 18644 9588 18672
rect 9582 18632 9588 18644
rect 9640 18632 9646 18684
rect 9858 18632 9864 18684
rect 9916 18672 9922 18684
rect 10689 18675 10747 18681
rect 10689 18672 10701 18675
rect 9916 18644 10701 18672
rect 9916 18632 9922 18644
rect 10689 18641 10701 18644
rect 10735 18641 10747 18675
rect 12802 18672 12808 18684
rect 12763 18644 12808 18672
rect 10689 18635 10747 18641
rect 12802 18632 12808 18644
rect 12860 18632 12866 18684
rect 16574 18632 16580 18684
rect 16632 18672 16638 18684
rect 17129 18675 17187 18681
rect 17129 18672 17141 18675
rect 16632 18644 17141 18672
rect 16632 18632 16638 18644
rect 17129 18641 17141 18644
rect 17175 18641 17187 18675
rect 17129 18635 17187 18641
rect 17954 18632 17960 18684
rect 18012 18672 18018 18684
rect 18049 18675 18107 18681
rect 18049 18672 18061 18675
rect 18012 18644 18061 18672
rect 18012 18632 18018 18644
rect 18049 18641 18061 18644
rect 18095 18641 18107 18675
rect 18248 18672 18276 18712
rect 18325 18709 18337 18743
rect 18371 18740 18383 18743
rect 18506 18740 18512 18752
rect 18371 18712 18512 18740
rect 18371 18709 18383 18712
rect 18325 18703 18383 18709
rect 18506 18700 18512 18712
rect 18564 18700 18570 18752
rect 21450 18740 21456 18752
rect 19352 18712 21456 18740
rect 19352 18672 19380 18712
rect 21450 18700 21456 18712
rect 21508 18700 21514 18752
rect 18248 18644 19380 18672
rect 19521 18675 19579 18681
rect 18049 18635 18107 18641
rect 19521 18641 19533 18675
rect 19567 18672 19579 18675
rect 20441 18675 20499 18681
rect 19567 18644 19840 18672
rect 19567 18641 19579 18644
rect 19521 18635 19579 18641
rect 5442 18604 5448 18616
rect 5403 18576 5448 18604
rect 5442 18564 5448 18576
rect 5500 18564 5506 18616
rect 6546 18564 6552 18616
rect 6604 18604 6610 18616
rect 6825 18607 6883 18613
rect 6825 18604 6837 18607
rect 6604 18576 6837 18604
rect 6604 18564 6610 18576
rect 6825 18573 6837 18576
rect 6871 18573 6883 18607
rect 6825 18567 6883 18573
rect 7926 18564 7932 18616
rect 7984 18604 7990 18616
rect 8481 18607 8539 18613
rect 8481 18604 8493 18607
rect 7984 18576 8493 18604
rect 7984 18564 7990 18576
rect 8481 18573 8493 18576
rect 8527 18573 8539 18607
rect 8481 18567 8539 18573
rect 9490 18564 9496 18616
rect 9548 18604 9554 18616
rect 9769 18607 9827 18613
rect 9769 18604 9781 18607
rect 9548 18576 9781 18604
rect 9548 18564 9554 18576
rect 9769 18573 9781 18576
rect 9815 18604 9827 18607
rect 9950 18604 9956 18616
rect 9815 18576 9956 18604
rect 9815 18573 9827 18576
rect 9769 18567 9827 18573
rect 9950 18564 9956 18576
rect 10008 18564 10014 18616
rect 12989 18607 13047 18613
rect 12989 18573 13001 18607
rect 13035 18573 13047 18607
rect 13446 18604 13452 18616
rect 13407 18576 13452 18604
rect 12989 18567 13047 18573
rect 7834 18496 7840 18548
rect 7892 18536 7898 18548
rect 10594 18536 10600 18548
rect 7892 18508 10600 18536
rect 7892 18496 7898 18508
rect 10594 18496 10600 18508
rect 10652 18496 10658 18548
rect 12069 18539 12127 18545
rect 12069 18505 12081 18539
rect 12115 18536 12127 18539
rect 12618 18536 12624 18548
rect 12115 18508 12624 18536
rect 12115 18505 12127 18508
rect 12069 18499 12127 18505
rect 12618 18496 12624 18508
rect 12676 18536 12682 18548
rect 13004 18536 13032 18567
rect 13446 18564 13452 18576
rect 13504 18564 13510 18616
rect 15105 18607 15163 18613
rect 15105 18573 15117 18607
rect 15151 18573 15163 18607
rect 15105 18567 15163 18573
rect 12676 18508 13032 18536
rect 12676 18496 12682 18508
rect 290 18428 296 18480
rect 348 18468 354 18480
rect 3510 18468 3516 18480
rect 348 18440 3516 18468
rect 348 18428 354 18440
rect 3510 18428 3516 18440
rect 3568 18428 3574 18480
rect 3602 18428 3608 18480
rect 3660 18468 3666 18480
rect 4246 18468 4252 18480
rect 3660 18440 4252 18468
rect 3660 18428 3666 18440
rect 4246 18428 4252 18440
rect 4304 18428 4310 18480
rect 4801 18471 4859 18477
rect 4801 18437 4813 18471
rect 4847 18468 4859 18471
rect 5258 18468 5264 18480
rect 4847 18440 5264 18468
rect 4847 18437 4859 18440
rect 4801 18431 4859 18437
rect 5258 18428 5264 18440
rect 5316 18428 5322 18480
rect 7466 18428 7472 18480
rect 7524 18468 7530 18480
rect 8478 18468 8484 18480
rect 7524 18440 8484 18468
rect 7524 18428 7530 18440
rect 8478 18428 8484 18440
rect 8536 18428 8542 18480
rect 9217 18471 9275 18477
rect 9217 18437 9229 18471
rect 9263 18468 9275 18471
rect 11790 18468 11796 18480
rect 9263 18440 11796 18468
rect 9263 18437 9275 18440
rect 9217 18431 9275 18437
rect 11790 18428 11796 18440
rect 11848 18428 11854 18480
rect 12434 18468 12440 18480
rect 12395 18440 12440 18468
rect 12434 18428 12440 18440
rect 12492 18428 12498 18480
rect 13464 18468 13492 18564
rect 15120 18468 15148 18567
rect 16482 18564 16488 18616
rect 16540 18604 16546 18616
rect 17313 18607 17371 18613
rect 17313 18604 17325 18607
rect 16540 18576 17325 18604
rect 16540 18564 16546 18576
rect 17313 18573 17325 18576
rect 17359 18573 17371 18607
rect 19702 18604 19708 18616
rect 19663 18576 19708 18604
rect 17313 18567 17371 18573
rect 19702 18564 19708 18576
rect 19760 18564 19766 18616
rect 19812 18604 19840 18644
rect 20441 18641 20453 18675
rect 20487 18672 20499 18675
rect 20533 18675 20591 18681
rect 20533 18672 20545 18675
rect 20487 18644 20545 18672
rect 20487 18641 20499 18644
rect 20441 18635 20499 18641
rect 20533 18641 20545 18644
rect 20579 18641 20591 18675
rect 20533 18635 20591 18641
rect 19886 18604 19892 18616
rect 19812 18576 19892 18604
rect 19886 18564 19892 18576
rect 19944 18564 19950 18616
rect 16390 18496 16396 18548
rect 16448 18536 16454 18548
rect 20530 18536 20536 18548
rect 16448 18508 20536 18536
rect 16448 18496 16454 18508
rect 20530 18496 20536 18508
rect 20588 18496 20594 18548
rect 16482 18468 16488 18480
rect 13464 18440 15148 18468
rect 16443 18440 16488 18468
rect 16482 18428 16488 18440
rect 16540 18428 16546 18480
rect 17494 18428 17500 18480
rect 17552 18468 17558 18480
rect 21174 18468 21180 18480
rect 17552 18440 21180 18468
rect 17552 18428 17558 18440
rect 21174 18428 21180 18440
rect 21232 18428 21238 18480
rect 1104 18378 21620 18400
rect 1104 18326 4414 18378
rect 4466 18326 4478 18378
rect 4530 18326 4542 18378
rect 4594 18326 4606 18378
rect 4658 18326 11278 18378
rect 11330 18326 11342 18378
rect 11394 18326 11406 18378
rect 11458 18326 11470 18378
rect 11522 18326 18142 18378
rect 18194 18326 18206 18378
rect 18258 18326 18270 18378
rect 18322 18326 18334 18378
rect 18386 18326 21620 18378
rect 1104 18304 21620 18326
rect 6914 18224 6920 18276
rect 6972 18264 6978 18276
rect 6972 18236 11100 18264
rect 6972 18224 6978 18236
rect 7650 18156 7656 18208
rect 7708 18196 7714 18208
rect 11072 18196 11100 18236
rect 11146 18224 11152 18276
rect 11204 18264 11210 18276
rect 19705 18267 19763 18273
rect 11204 18236 19656 18264
rect 11204 18224 11210 18236
rect 13357 18199 13415 18205
rect 7708 18168 8984 18196
rect 11072 18168 11836 18196
rect 7708 18156 7714 18168
rect 3510 18088 3516 18140
rect 3568 18128 3574 18140
rect 7834 18128 7840 18140
rect 3568 18100 7840 18128
rect 3568 18088 3574 18100
rect 7834 18088 7840 18100
rect 7892 18088 7898 18140
rect 8021 18131 8079 18137
rect 8021 18097 8033 18131
rect 8067 18128 8079 18131
rect 8202 18128 8208 18140
rect 8067 18100 8208 18128
rect 8067 18097 8079 18100
rect 8021 18091 8079 18097
rect 8202 18088 8208 18100
rect 8260 18088 8266 18140
rect 8570 18088 8576 18140
rect 8628 18128 8634 18140
rect 8956 18137 8984 18168
rect 8849 18131 8907 18137
rect 8849 18128 8861 18131
rect 8628 18100 8861 18128
rect 8628 18088 8634 18100
rect 8849 18097 8861 18100
rect 8895 18097 8907 18131
rect 8849 18091 8907 18097
rect 8941 18131 8999 18137
rect 8941 18097 8953 18131
rect 8987 18097 8999 18131
rect 8941 18091 8999 18097
rect 10781 18131 10839 18137
rect 10781 18097 10793 18131
rect 10827 18128 10839 18131
rect 11698 18128 11704 18140
rect 10827 18100 11704 18128
rect 10827 18097 10839 18100
rect 10781 18091 10839 18097
rect 11698 18088 11704 18100
rect 11756 18088 11762 18140
rect 11808 18128 11836 18168
rect 13357 18165 13369 18199
rect 13403 18196 13415 18199
rect 19518 18196 19524 18208
rect 13403 18168 19524 18196
rect 13403 18165 13415 18168
rect 13357 18159 13415 18165
rect 19518 18156 19524 18168
rect 19576 18156 19582 18208
rect 19628 18196 19656 18236
rect 19705 18233 19717 18267
rect 19751 18264 19763 18267
rect 19978 18264 19984 18276
rect 19751 18236 19984 18264
rect 19751 18233 19763 18236
rect 19705 18227 19763 18233
rect 19978 18224 19984 18236
rect 20036 18224 20042 18276
rect 19886 18196 19892 18208
rect 19628 18168 19892 18196
rect 19886 18156 19892 18168
rect 19944 18156 19950 18208
rect 14001 18131 14059 18137
rect 11808 18100 13952 18128
rect 5258 18060 5264 18072
rect 5219 18032 5264 18060
rect 5258 18020 5264 18032
rect 5316 18020 5322 18072
rect 7745 18063 7803 18069
rect 7745 18029 7757 18063
rect 7791 18060 7803 18063
rect 7926 18060 7932 18072
rect 7791 18032 7932 18060
rect 7791 18029 7803 18032
rect 7745 18023 7803 18029
rect 7926 18020 7932 18032
rect 7984 18020 7990 18072
rect 8386 18020 8392 18072
rect 8444 18060 8450 18072
rect 8757 18063 8815 18069
rect 8757 18060 8769 18063
rect 8444 18032 8769 18060
rect 8444 18020 8450 18032
rect 8757 18029 8769 18032
rect 8803 18029 8815 18063
rect 8757 18023 8815 18029
rect 9582 18020 9588 18072
rect 9640 18060 9646 18072
rect 11882 18060 11888 18072
rect 9640 18032 11888 18060
rect 9640 18020 9646 18032
rect 11882 18020 11888 18032
rect 11940 18020 11946 18072
rect 12434 18020 12440 18072
rect 12492 18060 12498 18072
rect 13817 18063 13875 18069
rect 13817 18060 13829 18063
rect 12492 18032 13829 18060
rect 12492 18020 12498 18032
rect 13817 18029 13829 18032
rect 13863 18029 13875 18063
rect 13924 18060 13952 18100
rect 14001 18097 14013 18131
rect 14047 18128 14059 18131
rect 14090 18128 14096 18140
rect 14047 18100 14096 18128
rect 14047 18097 14059 18100
rect 14001 18091 14059 18097
rect 14090 18088 14096 18100
rect 14148 18088 14154 18140
rect 16574 18128 16580 18140
rect 16535 18100 16580 18128
rect 16574 18088 16580 18100
rect 16632 18088 16638 18140
rect 19150 18088 19156 18140
rect 19208 18128 19214 18140
rect 20162 18128 20168 18140
rect 19208 18100 20168 18128
rect 19208 18088 19214 18100
rect 20162 18088 20168 18100
rect 20220 18088 20226 18140
rect 16850 18060 16856 18072
rect 13924 18032 16856 18060
rect 13817 18023 13875 18029
rect 16850 18020 16856 18032
rect 16908 18020 16914 18072
rect 19518 18060 19524 18072
rect 19479 18032 19524 18060
rect 19518 18020 19524 18032
rect 19576 18020 19582 18072
rect 19794 18020 19800 18072
rect 19852 18060 19858 18072
rect 21358 18060 21364 18072
rect 19852 18032 21364 18060
rect 19852 18020 19858 18032
rect 21358 18020 21364 18032
rect 21416 18020 21422 18072
rect 5534 17992 5540 18004
rect 5495 17964 5540 17992
rect 5534 17952 5540 17964
rect 5592 17952 5598 18004
rect 13725 17995 13783 18001
rect 7392 17964 13676 17992
rect 3050 17884 3056 17936
rect 3108 17924 3114 17936
rect 5902 17924 5908 17936
rect 3108 17896 5908 17924
rect 3108 17884 3114 17896
rect 5902 17884 5908 17896
rect 5960 17884 5966 17936
rect 7392 17933 7420 17964
rect 7377 17927 7435 17933
rect 7377 17893 7389 17927
rect 7423 17893 7435 17927
rect 7377 17887 7435 17893
rect 7837 17927 7895 17933
rect 7837 17893 7849 17927
rect 7883 17924 7895 17927
rect 8389 17927 8447 17933
rect 8389 17924 8401 17927
rect 7883 17896 8401 17924
rect 7883 17893 7895 17896
rect 7837 17887 7895 17893
rect 8389 17893 8401 17896
rect 8435 17893 8447 17927
rect 8389 17887 8447 17893
rect 8846 17884 8852 17936
rect 8904 17924 8910 17936
rect 11698 17924 11704 17936
rect 8904 17896 11704 17924
rect 8904 17884 8910 17896
rect 11698 17884 11704 17896
rect 11756 17884 11762 17936
rect 12526 17884 12532 17936
rect 12584 17924 12590 17936
rect 12986 17924 12992 17936
rect 12584 17896 12992 17924
rect 12584 17884 12590 17896
rect 12986 17884 12992 17896
rect 13044 17884 13050 17936
rect 13648 17924 13676 17964
rect 13725 17961 13737 17995
rect 13771 17992 13783 17995
rect 13998 17992 14004 18004
rect 13771 17964 14004 17992
rect 13771 17961 13783 17964
rect 13725 17955 13783 17961
rect 13998 17952 14004 17964
rect 14056 17952 14062 18004
rect 19426 17992 19432 18004
rect 14108 17964 19432 17992
rect 14108 17924 14136 17964
rect 19426 17952 19432 17964
rect 19484 17952 19490 18004
rect 21082 17952 21088 18004
rect 21140 17992 21146 18004
rect 22462 17992 22468 18004
rect 21140 17964 22468 17992
rect 21140 17952 21146 17964
rect 22462 17952 22468 17964
rect 22520 17952 22526 18004
rect 13648 17896 14136 17924
rect 14182 17884 14188 17936
rect 14240 17924 14246 17936
rect 15010 17924 15016 17936
rect 14240 17896 15016 17924
rect 14240 17884 14246 17896
rect 15010 17884 15016 17896
rect 15068 17884 15074 17936
rect 15286 17884 15292 17936
rect 15344 17924 15350 17936
rect 16390 17924 16396 17936
rect 15344 17896 16396 17924
rect 15344 17884 15350 17896
rect 16390 17884 16396 17896
rect 16448 17884 16454 17936
rect 19610 17884 19616 17936
rect 19668 17924 19674 17936
rect 20254 17924 20260 17936
rect 19668 17896 20260 17924
rect 19668 17884 19674 17896
rect 20254 17884 20260 17896
rect 20312 17884 20318 17936
rect 20622 17884 20628 17936
rect 20680 17924 20686 17936
rect 21910 17924 21916 17936
rect 20680 17896 21916 17924
rect 20680 17884 20686 17896
rect 21910 17884 21916 17896
rect 21968 17884 21974 17936
rect 1104 17834 21620 17856
rect 1104 17782 7846 17834
rect 7898 17782 7910 17834
rect 7962 17782 7974 17834
rect 8026 17782 8038 17834
rect 8090 17782 14710 17834
rect 14762 17782 14774 17834
rect 14826 17782 14838 17834
rect 14890 17782 14902 17834
rect 14954 17782 21620 17834
rect 1104 17760 21620 17782
rect 2866 17720 2872 17732
rect 2827 17692 2872 17720
rect 2866 17680 2872 17692
rect 2924 17680 2930 17732
rect 4062 17680 4068 17732
rect 4120 17720 4126 17732
rect 12342 17720 12348 17732
rect 4120 17692 12348 17720
rect 4120 17680 4126 17692
rect 12342 17680 12348 17692
rect 12400 17680 12406 17732
rect 20438 17720 20444 17732
rect 20399 17692 20444 17720
rect 20438 17680 20444 17692
rect 20496 17680 20502 17732
rect 20990 17720 20996 17732
rect 20951 17692 20996 17720
rect 20990 17680 20996 17692
rect 21048 17680 21054 17732
rect 1670 17652 1676 17664
rect 1504 17624 1676 17652
rect 1504 17593 1532 17624
rect 1670 17612 1676 17624
rect 1728 17652 1734 17664
rect 2406 17652 2412 17664
rect 1728 17624 2412 17652
rect 1728 17612 1734 17624
rect 2406 17612 2412 17624
rect 2464 17612 2470 17664
rect 5252 17655 5310 17661
rect 5252 17621 5264 17655
rect 5298 17652 5310 17655
rect 5442 17652 5448 17664
rect 5298 17624 5448 17652
rect 5298 17621 5310 17624
rect 5252 17615 5310 17621
rect 5442 17612 5448 17624
rect 5500 17612 5506 17664
rect 1489 17587 1547 17593
rect 1489 17553 1501 17587
rect 1535 17553 1547 17587
rect 1489 17547 1547 17553
rect 1756 17587 1814 17593
rect 1756 17553 1768 17587
rect 1802 17584 1814 17587
rect 3142 17584 3148 17596
rect 1802 17556 3148 17584
rect 1802 17553 1814 17556
rect 1756 17547 1814 17553
rect 3142 17544 3148 17556
rect 3200 17544 3206 17596
rect 5534 17544 5540 17596
rect 5592 17584 5598 17596
rect 19705 17587 19763 17593
rect 19705 17584 19717 17587
rect 5592 17556 19717 17584
rect 5592 17544 5598 17556
rect 19705 17553 19717 17556
rect 19751 17553 19763 17587
rect 20254 17584 20260 17596
rect 20215 17556 20260 17584
rect 19705 17547 19763 17553
rect 20254 17544 20260 17556
rect 20312 17544 20318 17596
rect 20346 17544 20352 17596
rect 20404 17584 20410 17596
rect 20809 17587 20867 17593
rect 20809 17584 20821 17587
rect 20404 17556 20821 17584
rect 20404 17544 20410 17556
rect 20809 17553 20821 17556
rect 20855 17553 20867 17587
rect 20809 17547 20867 17553
rect 3326 17516 3332 17528
rect 3287 17488 3332 17516
rect 3326 17476 3332 17488
rect 3384 17476 3390 17528
rect 4985 17519 5043 17525
rect 4985 17485 4997 17519
rect 5031 17485 5043 17519
rect 4985 17479 5043 17485
rect 5000 17380 5028 17479
rect 10778 17476 10784 17528
rect 10836 17516 10842 17528
rect 17034 17516 17040 17528
rect 10836 17488 17040 17516
rect 10836 17476 10842 17488
rect 17034 17476 17040 17488
rect 17092 17476 17098 17528
rect 6914 17408 6920 17460
rect 6972 17448 6978 17460
rect 18690 17448 18696 17460
rect 6972 17420 18696 17448
rect 6972 17408 6978 17420
rect 18690 17408 18696 17420
rect 18748 17408 18754 17460
rect 5718 17380 5724 17392
rect 5000 17352 5724 17380
rect 5718 17340 5724 17352
rect 5776 17340 5782 17392
rect 6365 17383 6423 17389
rect 6365 17349 6377 17383
rect 6411 17380 6423 17383
rect 9122 17380 9128 17392
rect 6411 17352 9128 17380
rect 6411 17349 6423 17352
rect 6365 17343 6423 17349
rect 9122 17340 9128 17352
rect 9180 17340 9186 17392
rect 12342 17340 12348 17392
rect 12400 17380 12406 17392
rect 17862 17380 17868 17392
rect 12400 17352 17868 17380
rect 12400 17340 12406 17352
rect 17862 17340 17868 17352
rect 17920 17340 17926 17392
rect 19886 17380 19892 17392
rect 19847 17352 19892 17380
rect 19886 17340 19892 17352
rect 19944 17340 19950 17392
rect 21726 17312 21732 17324
rect 1104 17290 21620 17312
rect 1104 17238 4414 17290
rect 4466 17238 4478 17290
rect 4530 17238 4542 17290
rect 4594 17238 4606 17290
rect 4658 17238 11278 17290
rect 11330 17238 11342 17290
rect 11394 17238 11406 17290
rect 11458 17238 11470 17290
rect 11522 17238 18142 17290
rect 18194 17238 18206 17290
rect 18258 17238 18270 17290
rect 18322 17238 18334 17290
rect 18386 17238 21620 17290
rect 21687 17284 21732 17312
rect 21726 17272 21732 17284
rect 21784 17272 21790 17324
rect 1104 17216 21620 17238
rect 7650 17136 7656 17188
rect 7708 17176 7714 17188
rect 7929 17179 7987 17185
rect 7929 17176 7941 17179
rect 7708 17148 7941 17176
rect 7708 17136 7714 17148
rect 7929 17145 7941 17148
rect 7975 17145 7987 17179
rect 7929 17139 7987 17145
rect 12621 17179 12679 17185
rect 12621 17145 12633 17179
rect 12667 17176 12679 17179
rect 15746 17176 15752 17188
rect 12667 17148 15752 17176
rect 12667 17145 12679 17148
rect 12621 17139 12679 17145
rect 15746 17136 15752 17148
rect 15804 17136 15810 17188
rect 17862 17176 17868 17188
rect 17823 17148 17868 17176
rect 17862 17136 17868 17148
rect 17920 17136 17926 17188
rect 17954 17136 17960 17188
rect 18012 17176 18018 17188
rect 18141 17179 18199 17185
rect 18141 17176 18153 17179
rect 18012 17148 18153 17176
rect 18012 17136 18018 17148
rect 18141 17145 18153 17148
rect 18187 17145 18199 17179
rect 18141 17139 18199 17145
rect 3142 17068 3148 17120
rect 3200 17108 3206 17120
rect 9769 17111 9827 17117
rect 3200 17080 4660 17108
rect 3200 17068 3206 17080
rect 2866 17000 2872 17052
rect 2924 17040 2930 17052
rect 3513 17043 3571 17049
rect 3513 17040 3525 17043
rect 2924 17012 3525 17040
rect 2924 17000 2930 17012
rect 3513 17009 3525 17012
rect 3559 17009 3571 17043
rect 3513 17003 3571 17009
rect 4154 17000 4160 17052
rect 4212 17040 4218 17052
rect 4632 17049 4660 17080
rect 9769 17077 9781 17111
rect 9815 17108 9827 17111
rect 9815 17080 15884 17108
rect 9815 17077 9827 17080
rect 9769 17071 9827 17077
rect 4525 17043 4583 17049
rect 4525 17040 4537 17043
rect 4212 17012 4537 17040
rect 4212 17000 4218 17012
rect 4525 17009 4537 17012
rect 4571 17009 4583 17043
rect 4525 17003 4583 17009
rect 4617 17043 4675 17049
rect 4617 17009 4629 17043
rect 4663 17009 4675 17043
rect 4617 17003 4675 17009
rect 5626 17000 5632 17052
rect 5684 17040 5690 17052
rect 9122 17040 9128 17052
rect 5684 17012 6684 17040
rect 9083 17012 9128 17040
rect 5684 17000 5690 17012
rect 3326 16972 3332 16984
rect 3287 16944 3332 16972
rect 3326 16932 3332 16944
rect 3384 16932 3390 16984
rect 5718 16932 5724 16984
rect 5776 16972 5782 16984
rect 6546 16972 6552 16984
rect 5776 16944 6552 16972
rect 5776 16932 5782 16944
rect 6546 16932 6552 16944
rect 6604 16932 6610 16984
rect 6656 16972 6684 17012
rect 9122 17000 9128 17012
rect 9180 17000 9186 17052
rect 10410 17040 10416 17052
rect 10371 17012 10416 17040
rect 10410 17000 10416 17012
rect 10468 17000 10474 17052
rect 12342 17040 12348 17052
rect 12303 17012 12348 17040
rect 12342 17000 12348 17012
rect 12400 17000 12406 17052
rect 12894 17000 12900 17052
rect 12952 17040 12958 17052
rect 13357 17043 13415 17049
rect 13357 17040 13369 17043
rect 12952 17012 13369 17040
rect 12952 17000 12958 17012
rect 13357 17009 13369 17012
rect 13403 17009 13415 17043
rect 15856 17040 15884 17080
rect 17880 17040 17908 17136
rect 18693 17043 18751 17049
rect 18693 17040 18705 17043
rect 15856 17012 16620 17040
rect 17880 17012 18705 17040
rect 13357 17003 13415 17009
rect 9033 16975 9091 16981
rect 9033 16972 9045 16975
rect 6656 16944 9045 16972
rect 9033 16941 9045 16944
rect 9079 16941 9091 16975
rect 9033 16935 9091 16941
rect 10962 16932 10968 16984
rect 11020 16972 11026 16984
rect 12253 16975 12311 16981
rect 12253 16972 12265 16975
rect 11020 16944 12265 16972
rect 11020 16932 11026 16944
rect 12253 16941 12265 16944
rect 12299 16941 12311 16975
rect 12253 16935 12311 16941
rect 12802 16932 12808 16984
rect 12860 16972 12866 16984
rect 14182 16972 14188 16984
rect 12860 16944 14188 16972
rect 12860 16932 12866 16944
rect 14182 16932 14188 16944
rect 14240 16932 14246 16984
rect 15562 16932 15568 16984
rect 15620 16972 15626 16984
rect 16485 16975 16543 16981
rect 16485 16972 16497 16975
rect 15620 16944 16497 16972
rect 15620 16932 15626 16944
rect 16485 16941 16497 16944
rect 16531 16941 16543 16975
rect 16592 16972 16620 17012
rect 18693 17009 18705 17012
rect 18739 17009 18751 17043
rect 20254 17040 20260 17052
rect 20215 17012 20260 17040
rect 18693 17003 18751 17009
rect 20254 17000 20260 17012
rect 20312 17000 20318 17052
rect 19245 16975 19303 16981
rect 19245 16972 19257 16975
rect 16592 16944 19257 16972
rect 16485 16935 16543 16941
rect 19245 16941 19257 16944
rect 19291 16941 19303 16975
rect 19978 16972 19984 16984
rect 19939 16944 19984 16972
rect 19245 16935 19303 16941
rect 19978 16932 19984 16944
rect 20036 16932 20042 16984
rect 6816 16907 6874 16913
rect 6816 16873 6828 16907
rect 6862 16904 6874 16907
rect 7098 16904 7104 16916
rect 6862 16876 7104 16904
rect 6862 16873 6874 16876
rect 6816 16867 6874 16873
rect 7098 16864 7104 16876
rect 7156 16864 7162 16916
rect 10229 16907 10287 16913
rect 10229 16904 10241 16907
rect 8588 16876 10241 16904
rect 2958 16836 2964 16848
rect 2919 16808 2964 16836
rect 2958 16796 2964 16808
rect 3016 16796 3022 16848
rect 3421 16839 3479 16845
rect 3421 16805 3433 16839
rect 3467 16836 3479 16839
rect 4065 16839 4123 16845
rect 4065 16836 4077 16839
rect 3467 16808 4077 16836
rect 3467 16805 3479 16808
rect 3421 16799 3479 16805
rect 4065 16805 4077 16808
rect 4111 16805 4123 16839
rect 4065 16799 4123 16805
rect 4433 16839 4491 16845
rect 4433 16805 4445 16839
rect 4479 16836 4491 16839
rect 8386 16836 8392 16848
rect 4479 16808 8392 16836
rect 4479 16805 4491 16808
rect 4433 16799 4491 16805
rect 8386 16796 8392 16808
rect 8444 16796 8450 16848
rect 8588 16845 8616 16876
rect 10229 16873 10241 16876
rect 10275 16873 10287 16907
rect 13265 16907 13323 16913
rect 13265 16904 13277 16907
rect 10229 16867 10287 16873
rect 11808 16876 13277 16904
rect 8573 16839 8631 16845
rect 8573 16805 8585 16839
rect 8619 16805 8631 16839
rect 8938 16836 8944 16848
rect 8899 16808 8944 16836
rect 8573 16799 8631 16805
rect 8938 16796 8944 16808
rect 8996 16796 9002 16848
rect 10134 16836 10140 16848
rect 10095 16808 10140 16836
rect 10134 16796 10140 16808
rect 10192 16796 10198 16848
rect 11808 16845 11836 16876
rect 13265 16873 13277 16876
rect 13311 16873 13323 16907
rect 13265 16867 13323 16873
rect 16752 16907 16810 16913
rect 16752 16873 16764 16907
rect 16798 16904 16810 16907
rect 16942 16904 16948 16916
rect 16798 16876 16948 16904
rect 16798 16873 16810 16876
rect 16752 16867 16810 16873
rect 16942 16864 16948 16876
rect 17000 16864 17006 16916
rect 17954 16864 17960 16916
rect 18012 16904 18018 16916
rect 18601 16907 18659 16913
rect 18601 16904 18613 16907
rect 18012 16876 18613 16904
rect 18012 16864 18018 16876
rect 18601 16873 18613 16876
rect 18647 16873 18659 16907
rect 18601 16867 18659 16873
rect 19521 16907 19579 16913
rect 19521 16873 19533 16907
rect 19567 16904 19579 16907
rect 20530 16904 20536 16916
rect 19567 16876 20536 16904
rect 19567 16873 19579 16876
rect 19521 16867 19579 16873
rect 20530 16864 20536 16876
rect 20588 16864 20594 16916
rect 11793 16839 11851 16845
rect 11793 16805 11805 16839
rect 11839 16805 11851 16839
rect 11793 16799 11851 16805
rect 12161 16839 12219 16845
rect 12161 16805 12173 16839
rect 12207 16836 12219 16839
rect 12621 16839 12679 16845
rect 12621 16836 12633 16839
rect 12207 16808 12633 16836
rect 12207 16805 12219 16808
rect 12161 16799 12219 16805
rect 12621 16805 12633 16808
rect 12667 16805 12679 16839
rect 12802 16836 12808 16848
rect 12763 16808 12808 16836
rect 12621 16799 12679 16805
rect 12802 16796 12808 16808
rect 12860 16796 12866 16848
rect 13170 16836 13176 16848
rect 13131 16808 13176 16836
rect 13170 16796 13176 16808
rect 13228 16796 13234 16848
rect 18046 16796 18052 16848
rect 18104 16836 18110 16848
rect 18509 16839 18567 16845
rect 18509 16836 18521 16839
rect 18104 16808 18521 16836
rect 18104 16796 18110 16808
rect 18509 16805 18521 16808
rect 18555 16805 18567 16839
rect 18509 16799 18567 16805
rect 1104 16746 21620 16768
rect 1104 16694 7846 16746
rect 7898 16694 7910 16746
rect 7962 16694 7974 16746
rect 8026 16694 8038 16746
rect 8090 16694 14710 16746
rect 14762 16694 14774 16746
rect 14826 16694 14838 16746
rect 14890 16694 14902 16746
rect 14954 16694 21620 16746
rect 1104 16672 21620 16694
rect 6914 16632 6920 16644
rect 6875 16604 6920 16632
rect 6914 16592 6920 16604
rect 6972 16592 6978 16644
rect 10137 16635 10195 16641
rect 10137 16601 10149 16635
rect 10183 16601 10195 16635
rect 11790 16632 11796 16644
rect 11703 16604 11796 16632
rect 10137 16595 10195 16601
rect 6546 16524 6552 16576
rect 6604 16564 6610 16576
rect 9024 16567 9082 16573
rect 6604 16536 8800 16564
rect 6604 16524 6610 16536
rect 2958 16456 2964 16508
rect 3016 16496 3022 16508
rect 8772 16505 8800 16536
rect 9024 16533 9036 16567
rect 9070 16564 9082 16567
rect 9122 16564 9128 16576
rect 9070 16536 9128 16564
rect 9070 16533 9082 16536
rect 9024 16527 9082 16533
rect 9122 16524 9128 16536
rect 9180 16524 9186 16576
rect 10152 16564 10180 16595
rect 11790 16592 11796 16604
rect 11848 16632 11854 16644
rect 12342 16632 12348 16644
rect 11848 16604 12348 16632
rect 11848 16592 11854 16604
rect 12342 16592 12348 16604
rect 12400 16592 12406 16644
rect 12802 16592 12808 16644
rect 12860 16632 12866 16644
rect 16942 16632 16948 16644
rect 12860 16604 16804 16632
rect 16903 16604 16948 16632
rect 12860 16592 12866 16604
rect 10410 16564 10416 16576
rect 10152 16536 10416 16564
rect 10410 16524 10416 16536
rect 10468 16564 10474 16576
rect 10658 16567 10716 16573
rect 10658 16564 10670 16567
rect 10468 16536 10670 16564
rect 10468 16524 10474 16536
rect 10658 16533 10670 16536
rect 10704 16533 10716 16567
rect 15562 16564 15568 16576
rect 10658 16527 10716 16533
rect 12820 16536 15568 16564
rect 3881 16499 3939 16505
rect 3881 16496 3893 16499
rect 3016 16468 3893 16496
rect 3016 16456 3022 16468
rect 3881 16465 3893 16468
rect 3927 16465 3939 16499
rect 3881 16459 3939 16465
rect 7285 16499 7343 16505
rect 7285 16465 7297 16499
rect 7331 16496 7343 16499
rect 7929 16499 7987 16505
rect 7929 16496 7941 16499
rect 7331 16468 7941 16496
rect 7331 16465 7343 16468
rect 7285 16459 7343 16465
rect 7929 16465 7941 16468
rect 7975 16465 7987 16499
rect 7929 16459 7987 16465
rect 8757 16499 8815 16505
rect 8757 16465 8769 16499
rect 8803 16496 8815 16499
rect 9766 16496 9772 16508
rect 8803 16468 9772 16496
rect 8803 16465 8815 16468
rect 8757 16459 8815 16465
rect 9766 16456 9772 16468
rect 9824 16496 9830 16508
rect 9824 16468 10456 16496
rect 9824 16456 9830 16468
rect 4154 16428 4160 16440
rect 4115 16400 4160 16428
rect 4154 16388 4160 16400
rect 4212 16388 4218 16440
rect 7374 16428 7380 16440
rect 7335 16400 7380 16428
rect 7374 16388 7380 16400
rect 7432 16388 7438 16440
rect 10428 16437 10456 16468
rect 7469 16431 7527 16437
rect 7469 16397 7481 16431
rect 7515 16397 7527 16431
rect 7469 16391 7527 16397
rect 10413 16431 10471 16437
rect 10413 16397 10425 16431
rect 10459 16397 10471 16431
rect 10413 16391 10471 16397
rect 7098 16320 7104 16372
rect 7156 16360 7162 16372
rect 7484 16360 7512 16391
rect 12710 16388 12716 16440
rect 12768 16428 12774 16440
rect 12820 16428 12848 16536
rect 15562 16524 15568 16536
rect 15620 16524 15626 16576
rect 15832 16567 15890 16573
rect 15832 16533 15844 16567
rect 15878 16564 15890 16567
rect 16482 16564 16488 16576
rect 15878 16536 16488 16564
rect 15878 16533 15890 16536
rect 15832 16527 15890 16533
rect 16482 16524 16488 16536
rect 16540 16524 16546 16576
rect 16776 16564 16804 16604
rect 16942 16592 16948 16604
rect 17000 16592 17006 16644
rect 18046 16632 18052 16644
rect 18007 16604 18052 16632
rect 18046 16592 18052 16604
rect 18104 16592 18110 16644
rect 20717 16635 20775 16641
rect 20717 16601 20729 16635
rect 20763 16632 20775 16635
rect 21729 16635 21787 16641
rect 21729 16632 21741 16635
rect 20763 16604 21741 16632
rect 20763 16601 20775 16604
rect 20717 16595 20775 16601
rect 21729 16601 21741 16604
rect 21775 16601 21787 16635
rect 21729 16595 21787 16601
rect 18969 16567 19027 16573
rect 16776 16536 18828 16564
rect 12894 16456 12900 16508
rect 12952 16496 12958 16508
rect 13245 16499 13303 16505
rect 13245 16496 13257 16499
rect 12952 16468 13257 16496
rect 12952 16456 12958 16468
rect 13245 16465 13257 16468
rect 13291 16465 13303 16499
rect 13245 16459 13303 16465
rect 15013 16499 15071 16505
rect 15013 16465 15025 16499
rect 15059 16496 15071 16499
rect 15470 16496 15476 16508
rect 15059 16468 15476 16496
rect 15059 16465 15071 16468
rect 15013 16459 15071 16465
rect 15470 16456 15476 16468
rect 15528 16456 15534 16508
rect 15580 16437 15608 16524
rect 18690 16496 18696 16508
rect 18651 16468 18696 16496
rect 18690 16456 18696 16468
rect 18748 16456 18754 16508
rect 18800 16496 18828 16536
rect 18969 16533 18981 16567
rect 19015 16564 19027 16567
rect 19518 16564 19524 16576
rect 19015 16536 19524 16564
rect 19015 16533 19027 16536
rect 18969 16527 19027 16533
rect 19518 16524 19524 16536
rect 19576 16524 19582 16576
rect 19705 16567 19763 16573
rect 19705 16533 19717 16567
rect 19751 16564 19763 16567
rect 20346 16564 20352 16576
rect 19751 16536 20352 16564
rect 19751 16533 19763 16536
rect 19705 16527 19763 16533
rect 20346 16524 20352 16536
rect 20404 16524 20410 16576
rect 19429 16499 19487 16505
rect 19429 16496 19441 16499
rect 18800 16468 19441 16496
rect 19429 16465 19441 16468
rect 19475 16465 19487 16499
rect 20530 16496 20536 16508
rect 20491 16468 20536 16496
rect 19429 16459 19487 16465
rect 20530 16456 20536 16468
rect 20588 16456 20594 16508
rect 12989 16431 13047 16437
rect 12989 16428 13001 16431
rect 12768 16400 13001 16428
rect 12768 16388 12774 16400
rect 12989 16397 13001 16400
rect 13035 16397 13047 16431
rect 12989 16391 13047 16397
rect 15565 16431 15623 16437
rect 15565 16397 15577 16431
rect 15611 16397 15623 16431
rect 15565 16391 15623 16397
rect 7156 16332 7512 16360
rect 7156 16320 7162 16332
rect 14366 16292 14372 16304
rect 14327 16264 14372 16292
rect 14366 16252 14372 16264
rect 14424 16252 14430 16304
rect 1104 16202 21620 16224
rect 1104 16150 4414 16202
rect 4466 16150 4478 16202
rect 4530 16150 4542 16202
rect 4594 16150 4606 16202
rect 4658 16150 11278 16202
rect 11330 16150 11342 16202
rect 11394 16150 11406 16202
rect 11458 16150 11470 16202
rect 11522 16150 18142 16202
rect 18194 16150 18206 16202
rect 18258 16150 18270 16202
rect 18322 16150 18334 16202
rect 18386 16150 21620 16202
rect 1104 16128 21620 16150
rect 3142 16088 3148 16100
rect 3103 16060 3148 16088
rect 3142 16048 3148 16060
rect 3200 16048 3206 16100
rect 4154 16048 4160 16100
rect 4212 16088 4218 16100
rect 7098 16088 7104 16100
rect 4212 16060 6960 16088
rect 7059 16060 7104 16088
rect 4212 16048 4218 16060
rect 6932 16020 6960 16060
rect 7098 16048 7104 16060
rect 7156 16048 7162 16100
rect 7374 16088 7380 16100
rect 7335 16060 7380 16088
rect 7374 16048 7380 16060
rect 7432 16048 7438 16100
rect 12894 16088 12900 16100
rect 8220 16060 12756 16088
rect 12855 16060 12900 16088
rect 8220 16020 8248 16060
rect 6932 15992 8248 16020
rect 12728 16020 12756 16060
rect 12894 16048 12900 16060
rect 12952 16048 12958 16100
rect 16577 16091 16635 16097
rect 16577 16057 16589 16091
rect 16623 16088 16635 16091
rect 17954 16088 17960 16100
rect 16623 16060 17960 16088
rect 16623 16057 16635 16060
rect 16577 16051 16635 16057
rect 17954 16048 17960 16060
rect 18012 16048 18018 16100
rect 20438 16088 20444 16100
rect 20399 16060 20444 16088
rect 20438 16048 20444 16060
rect 20496 16048 20502 16100
rect 12728 15992 20300 16020
rect 1670 15912 1676 15964
rect 1728 15952 1734 15964
rect 1765 15955 1823 15961
rect 1765 15952 1777 15955
rect 1728 15924 1777 15952
rect 1728 15912 1734 15924
rect 1765 15921 1777 15924
rect 1811 15921 1823 15955
rect 1765 15915 1823 15921
rect 1780 15884 1808 15915
rect 7742 15912 7748 15964
rect 7800 15952 7806 15964
rect 7837 15955 7895 15961
rect 7837 15952 7849 15955
rect 7800 15924 7849 15952
rect 7800 15912 7806 15924
rect 7837 15921 7849 15924
rect 7883 15921 7895 15955
rect 7837 15915 7895 15921
rect 7929 15955 7987 15961
rect 7929 15921 7941 15955
rect 7975 15921 7987 15955
rect 10134 15952 10140 15964
rect 10095 15924 10140 15952
rect 7929 15915 7987 15921
rect 3878 15884 3884 15896
rect 1780 15856 3884 15884
rect 3878 15844 3884 15856
rect 3936 15844 3942 15896
rect 5718 15884 5724 15896
rect 5679 15856 5724 15884
rect 5718 15844 5724 15856
rect 5776 15844 5782 15896
rect 5988 15887 6046 15893
rect 5988 15853 6000 15887
rect 6034 15884 6046 15887
rect 7944 15884 7972 15915
rect 10134 15912 10140 15924
rect 10192 15912 10198 15964
rect 13170 15952 13176 15964
rect 13131 15924 13176 15952
rect 13170 15912 13176 15924
rect 13228 15912 13234 15964
rect 14366 15912 14372 15964
rect 14424 15952 14430 15964
rect 14645 15955 14703 15961
rect 14645 15952 14657 15955
rect 14424 15924 14657 15952
rect 14424 15912 14430 15924
rect 14645 15921 14657 15924
rect 14691 15921 14703 15955
rect 15838 15952 15844 15964
rect 15799 15924 15844 15952
rect 14645 15915 14703 15921
rect 15838 15912 15844 15924
rect 15896 15912 15902 15964
rect 16942 15912 16948 15964
rect 17000 15952 17006 15964
rect 17129 15955 17187 15961
rect 17129 15952 17141 15955
rect 17000 15924 17141 15952
rect 17000 15912 17006 15924
rect 17129 15921 17141 15924
rect 17175 15921 17187 15955
rect 17129 15915 17187 15921
rect 6034 15856 7972 15884
rect 6034 15853 6046 15856
rect 5988 15847 6046 15853
rect 6196 15828 6224 15856
rect 11054 15844 11060 15896
rect 11112 15884 11118 15896
rect 11790 15893 11796 15896
rect 11517 15887 11575 15893
rect 11517 15884 11529 15887
rect 11112 15856 11529 15884
rect 11112 15844 11118 15856
rect 11517 15853 11529 15856
rect 11563 15853 11575 15887
rect 11784 15884 11796 15893
rect 11751 15856 11796 15884
rect 11517 15847 11575 15853
rect 11784 15847 11796 15856
rect 11790 15844 11796 15847
rect 11848 15844 11854 15896
rect 14553 15887 14611 15893
rect 14553 15884 14565 15887
rect 11900 15856 14565 15884
rect 2032 15819 2090 15825
rect 2032 15785 2044 15819
rect 2078 15816 2090 15819
rect 2958 15816 2964 15828
rect 2078 15788 2964 15816
rect 2078 15785 2090 15788
rect 2032 15779 2090 15785
rect 2958 15776 2964 15788
rect 3016 15776 3022 15828
rect 6178 15776 6184 15828
rect 6236 15776 6242 15828
rect 9030 15776 9036 15828
rect 9088 15816 9094 15828
rect 11900 15816 11928 15856
rect 14553 15853 14565 15856
rect 14599 15853 14611 15887
rect 14553 15847 14611 15853
rect 15470 15844 15476 15896
rect 15528 15884 15534 15896
rect 15657 15887 15715 15893
rect 15657 15884 15669 15887
rect 15528 15856 15669 15884
rect 15528 15844 15534 15856
rect 15657 15853 15669 15856
rect 15703 15853 15715 15887
rect 17034 15884 17040 15896
rect 16995 15856 17040 15884
rect 15657 15847 15715 15853
rect 17034 15844 17040 15856
rect 17092 15844 17098 15896
rect 18874 15884 18880 15896
rect 18835 15856 18880 15884
rect 18874 15844 18880 15856
rect 18932 15844 18938 15896
rect 19978 15884 19984 15896
rect 18984 15856 19984 15884
rect 15749 15819 15807 15825
rect 15749 15816 15761 15819
rect 9088 15788 11928 15816
rect 14108 15788 15761 15816
rect 9088 15776 9094 15788
rect 7742 15748 7748 15760
rect 7703 15720 7748 15748
rect 7742 15708 7748 15720
rect 7800 15708 7806 15760
rect 14108 15757 14136 15788
rect 15749 15785 15761 15788
rect 15795 15785 15807 15819
rect 18984 15816 19012 15856
rect 19978 15844 19984 15856
rect 20036 15844 20042 15896
rect 20272 15893 20300 15992
rect 20257 15887 20315 15893
rect 20257 15853 20269 15887
rect 20303 15853 20315 15887
rect 20257 15847 20315 15853
rect 15749 15779 15807 15785
rect 16776 15788 19012 15816
rect 19153 15819 19211 15825
rect 14093 15751 14151 15757
rect 14093 15717 14105 15751
rect 14139 15717 14151 15751
rect 14458 15748 14464 15760
rect 14419 15720 14464 15748
rect 14093 15711 14151 15717
rect 14458 15708 14464 15720
rect 14516 15708 14522 15760
rect 15289 15751 15347 15757
rect 15289 15717 15301 15751
rect 15335 15748 15347 15751
rect 16776 15748 16804 15788
rect 19153 15785 19165 15819
rect 19199 15816 19211 15819
rect 20162 15816 20168 15828
rect 19199 15788 20168 15816
rect 19199 15785 19211 15788
rect 19153 15779 19211 15785
rect 20162 15776 20168 15788
rect 20220 15776 20226 15828
rect 16942 15748 16948 15760
rect 15335 15720 16804 15748
rect 16903 15720 16948 15748
rect 15335 15717 15347 15720
rect 15289 15711 15347 15717
rect 16942 15708 16948 15720
rect 17000 15708 17006 15760
rect 1104 15658 21620 15680
rect 1104 15606 7846 15658
rect 7898 15606 7910 15658
rect 7962 15606 7974 15658
rect 8026 15606 8038 15658
rect 8090 15606 14710 15658
rect 14762 15606 14774 15658
rect 14826 15606 14838 15658
rect 14890 15606 14902 15658
rect 14954 15606 21620 15658
rect 1104 15584 21620 15606
rect 2958 15544 2964 15556
rect 2919 15516 2964 15544
rect 2958 15504 2964 15516
rect 3016 15504 3022 15556
rect 3237 15547 3295 15553
rect 3237 15513 3249 15547
rect 3283 15513 3295 15547
rect 6178 15544 6184 15556
rect 6139 15516 6184 15544
rect 3237 15507 3295 15513
rect 1581 15411 1639 15417
rect 1581 15377 1593 15411
rect 1627 15408 1639 15411
rect 1670 15408 1676 15420
rect 1627 15380 1676 15408
rect 1627 15377 1639 15380
rect 1581 15371 1639 15377
rect 1670 15368 1676 15380
rect 1728 15368 1734 15420
rect 1848 15411 1906 15417
rect 1848 15377 1860 15411
rect 1894 15408 1906 15411
rect 1894 15380 2912 15408
rect 1894 15377 1906 15380
rect 1848 15371 1906 15377
rect 2884 15204 2912 15380
rect 2976 15272 3004 15504
rect 3252 15476 3280 15507
rect 6178 15504 6184 15516
rect 6236 15504 6242 15556
rect 14458 15504 14464 15556
rect 14516 15544 14522 15556
rect 16942 15544 16948 15556
rect 14516 15516 16948 15544
rect 14516 15504 14522 15516
rect 16942 15504 16948 15516
rect 17000 15504 17006 15556
rect 19242 15504 19248 15556
rect 19300 15544 19306 15556
rect 20165 15547 20223 15553
rect 20165 15544 20177 15547
rect 19300 15516 20177 15544
rect 19300 15504 19306 15516
rect 20165 15513 20177 15516
rect 20211 15513 20223 15547
rect 20165 15507 20223 15513
rect 20717 15547 20775 15553
rect 20717 15513 20729 15547
rect 20763 15544 20775 15547
rect 21266 15544 21272 15556
rect 20763 15516 21272 15544
rect 20763 15513 20775 15516
rect 20717 15507 20775 15513
rect 21266 15504 21272 15516
rect 21324 15504 21330 15556
rect 18874 15476 18880 15488
rect 3252 15448 18880 15476
rect 18874 15436 18880 15448
rect 18932 15436 18938 15488
rect 3605 15411 3663 15417
rect 3605 15377 3617 15411
rect 3651 15408 3663 15411
rect 4249 15411 4307 15417
rect 4249 15408 4261 15411
rect 3651 15380 4261 15408
rect 3651 15377 3663 15380
rect 3605 15371 3663 15377
rect 4249 15377 4261 15380
rect 4295 15377 4307 15411
rect 4249 15371 4307 15377
rect 5068 15411 5126 15417
rect 5068 15377 5080 15411
rect 5114 15408 5126 15411
rect 6822 15408 6828 15420
rect 5114 15380 6828 15408
rect 5114 15377 5126 15380
rect 5068 15371 5126 15377
rect 6822 15368 6828 15380
rect 6880 15368 6886 15420
rect 7377 15411 7435 15417
rect 7377 15377 7389 15411
rect 7423 15408 7435 15411
rect 8202 15408 8208 15420
rect 7423 15380 8208 15408
rect 7423 15377 7435 15380
rect 7377 15371 7435 15377
rect 8202 15368 8208 15380
rect 8260 15368 8266 15420
rect 15102 15368 15108 15420
rect 15160 15408 15166 15420
rect 18969 15411 19027 15417
rect 18969 15408 18981 15411
rect 15160 15380 18981 15408
rect 15160 15368 15166 15380
rect 18969 15377 18981 15380
rect 19015 15377 19027 15411
rect 19978 15408 19984 15420
rect 19939 15380 19984 15408
rect 18969 15371 19027 15377
rect 19978 15368 19984 15380
rect 20036 15368 20042 15420
rect 20533 15411 20591 15417
rect 20533 15377 20545 15411
rect 20579 15377 20591 15411
rect 20533 15371 20591 15377
rect 3694 15340 3700 15352
rect 3655 15312 3700 15340
rect 3694 15300 3700 15312
rect 3752 15300 3758 15352
rect 3789 15343 3847 15349
rect 3789 15309 3801 15343
rect 3835 15309 3847 15343
rect 3789 15303 3847 15309
rect 3804 15272 3832 15303
rect 3878 15300 3884 15352
rect 3936 15340 3942 15352
rect 4801 15343 4859 15349
rect 4801 15340 4813 15343
rect 3936 15312 4813 15340
rect 3936 15300 3942 15312
rect 4801 15309 4813 15312
rect 4847 15309 4859 15343
rect 4801 15303 4859 15309
rect 19245 15343 19303 15349
rect 19245 15309 19257 15343
rect 19291 15340 19303 15343
rect 20548 15340 20576 15371
rect 19291 15312 20576 15340
rect 19291 15309 19303 15312
rect 19245 15303 19303 15309
rect 2976 15244 3832 15272
rect 3602 15204 3608 15216
rect 2884 15176 3608 15204
rect 3602 15164 3608 15176
rect 3660 15164 3666 15216
rect 4816 15204 4844 15303
rect 5718 15204 5724 15216
rect 4816 15176 5724 15204
rect 5718 15164 5724 15176
rect 5776 15204 5782 15216
rect 7193 15207 7251 15213
rect 7193 15204 7205 15207
rect 5776 15176 7205 15204
rect 5776 15164 5782 15176
rect 7193 15173 7205 15176
rect 7239 15173 7251 15207
rect 7193 15167 7251 15173
rect 10042 15164 10048 15216
rect 10100 15204 10106 15216
rect 18782 15204 18788 15216
rect 10100 15176 18788 15204
rect 10100 15164 10106 15176
rect 18782 15164 18788 15176
rect 18840 15164 18846 15216
rect 19518 15164 19524 15216
rect 19576 15204 19582 15216
rect 19794 15204 19800 15216
rect 19576 15176 19800 15204
rect 19576 15164 19582 15176
rect 19794 15164 19800 15176
rect 19852 15164 19858 15216
rect 1104 15114 21620 15136
rect 1104 15062 4414 15114
rect 4466 15062 4478 15114
rect 4530 15062 4542 15114
rect 4594 15062 4606 15114
rect 4658 15062 11278 15114
rect 11330 15062 11342 15114
rect 11394 15062 11406 15114
rect 11458 15062 11470 15114
rect 11522 15062 18142 15114
rect 18194 15062 18206 15114
rect 18258 15062 18270 15114
rect 18322 15062 18334 15114
rect 18386 15062 21620 15114
rect 1104 15040 21620 15062
rect 3694 14960 3700 15012
rect 3752 15000 3758 15012
rect 4065 15003 4123 15009
rect 4065 15000 4077 15003
rect 3752 14972 4077 15000
rect 3752 14960 3758 14972
rect 4065 14969 4077 14972
rect 4111 14969 4123 15003
rect 4065 14963 4123 14969
rect 9677 15003 9735 15009
rect 9677 14969 9689 15003
rect 9723 15000 9735 15003
rect 15102 15000 15108 15012
rect 9723 14972 15108 15000
rect 9723 14969 9735 14972
rect 9677 14963 9735 14969
rect 15102 14960 15108 14972
rect 15160 14960 15166 15012
rect 19886 15000 19892 15012
rect 19847 14972 19892 15000
rect 19886 14960 19892 14972
rect 19944 14960 19950 15012
rect 20438 15000 20444 15012
rect 20399 14972 20444 15000
rect 20438 14960 20444 14972
rect 20496 14960 20502 15012
rect 8021 14935 8079 14941
rect 8021 14901 8033 14935
rect 8067 14932 8079 14935
rect 8067 14904 10180 14932
rect 8067 14901 8079 14904
rect 8021 14895 8079 14901
rect 3602 14824 3608 14876
rect 3660 14864 3666 14876
rect 4617 14867 4675 14873
rect 4617 14864 4629 14867
rect 3660 14836 4629 14864
rect 3660 14824 3666 14836
rect 4617 14833 4629 14836
rect 4663 14833 4675 14867
rect 8478 14864 8484 14876
rect 8439 14836 8484 14864
rect 4617 14827 4675 14833
rect 8478 14824 8484 14836
rect 8536 14824 8542 14876
rect 8662 14864 8668 14876
rect 8623 14836 8668 14864
rect 8662 14824 8668 14836
rect 8720 14824 8726 14876
rect 10152 14873 10180 14904
rect 10962 14892 10968 14944
rect 11020 14932 11026 14944
rect 12710 14932 12716 14944
rect 11020 14904 12716 14932
rect 11020 14892 11026 14904
rect 12710 14892 12716 14904
rect 12768 14932 12774 14944
rect 13173 14935 13231 14941
rect 13173 14932 13185 14935
rect 12768 14904 13185 14932
rect 12768 14892 12774 14904
rect 13173 14901 13185 14904
rect 13219 14932 13231 14935
rect 14921 14935 14979 14941
rect 13219 14904 13584 14932
rect 13219 14901 13231 14904
rect 13173 14895 13231 14901
rect 10137 14867 10195 14873
rect 10137 14833 10149 14867
rect 10183 14833 10195 14867
rect 10137 14827 10195 14833
rect 10226 14824 10232 14876
rect 10284 14864 10290 14876
rect 10284 14836 10329 14864
rect 10284 14824 10290 14836
rect 11698 14824 11704 14876
rect 11756 14864 11762 14876
rect 13556 14873 13584 14904
rect 14921 14901 14933 14935
rect 14967 14932 14979 14935
rect 15194 14932 15200 14944
rect 14967 14904 15200 14932
rect 14967 14901 14979 14904
rect 14921 14895 14979 14901
rect 15194 14892 15200 14904
rect 15252 14932 15258 14944
rect 15838 14932 15844 14944
rect 15252 14904 15844 14932
rect 15252 14892 15258 14904
rect 15838 14892 15844 14904
rect 15896 14892 15902 14944
rect 12437 14867 12495 14873
rect 12437 14864 12449 14867
rect 11756 14836 12449 14864
rect 11756 14824 11762 14836
rect 12437 14833 12449 14836
rect 12483 14833 12495 14867
rect 12437 14827 12495 14833
rect 12529 14867 12587 14873
rect 12529 14833 12541 14867
rect 12575 14833 12587 14867
rect 12529 14827 12587 14833
rect 13541 14867 13599 14873
rect 13541 14833 13553 14867
rect 13587 14833 13599 14867
rect 17034 14864 17040 14876
rect 16995 14836 17040 14864
rect 13541 14827 13599 14833
rect 4246 14756 4252 14808
rect 4304 14796 4310 14808
rect 4525 14799 4583 14805
rect 4525 14796 4537 14799
rect 4304 14768 4537 14796
rect 4304 14756 4310 14768
rect 4525 14765 4537 14768
rect 4571 14765 4583 14799
rect 4525 14759 4583 14765
rect 7742 14756 7748 14808
rect 7800 14796 7806 14808
rect 12158 14796 12164 14808
rect 7800 14768 12164 14796
rect 7800 14756 7806 14768
rect 12158 14756 12164 14768
rect 12216 14756 12222 14808
rect 12342 14756 12348 14808
rect 12400 14796 12406 14808
rect 12544 14796 12572 14827
rect 13354 14796 13360 14808
rect 12400 14768 12572 14796
rect 13315 14768 13360 14796
rect 12400 14756 12406 14768
rect 13354 14756 13360 14768
rect 13412 14756 13418 14808
rect 4433 14731 4491 14737
rect 4433 14697 4445 14731
rect 4479 14728 4491 14731
rect 7760 14728 7788 14756
rect 4479 14700 7788 14728
rect 10045 14731 10103 14737
rect 4479 14697 4491 14700
rect 4433 14691 4491 14697
rect 10045 14697 10057 14731
rect 10091 14728 10103 14731
rect 10689 14731 10747 14737
rect 10689 14728 10701 14731
rect 10091 14700 10701 14728
rect 10091 14697 10103 14700
rect 10045 14691 10103 14697
rect 10689 14697 10701 14700
rect 10735 14697 10747 14731
rect 13556 14728 13584 14827
rect 17034 14824 17040 14836
rect 17092 14824 17098 14876
rect 19061 14867 19119 14873
rect 19061 14833 19073 14867
rect 19107 14864 19119 14867
rect 19978 14864 19984 14876
rect 19107 14836 19984 14864
rect 19107 14833 19119 14836
rect 19061 14827 19119 14833
rect 19978 14824 19984 14836
rect 20036 14824 20042 14876
rect 13808 14799 13866 14805
rect 13808 14765 13820 14799
rect 13854 14796 13866 14799
rect 14366 14796 14372 14808
rect 13854 14768 14372 14796
rect 13854 14765 13866 14768
rect 13808 14759 13866 14765
rect 14366 14756 14372 14768
rect 14424 14756 14430 14808
rect 18785 14799 18843 14805
rect 18785 14796 18797 14799
rect 16500 14768 18797 14796
rect 13722 14728 13728 14740
rect 13556 14700 13728 14728
rect 10689 14691 10747 14697
rect 13722 14688 13728 14700
rect 13780 14688 13786 14740
rect 8386 14660 8392 14672
rect 8347 14632 8392 14660
rect 8386 14620 8392 14632
rect 8444 14620 8450 14672
rect 11974 14660 11980 14672
rect 11935 14632 11980 14660
rect 11974 14620 11980 14632
rect 12032 14620 12038 14672
rect 12066 14620 12072 14672
rect 12124 14660 12130 14672
rect 16500 14669 16528 14768
rect 18785 14765 18797 14768
rect 18831 14765 18843 14799
rect 19702 14796 19708 14808
rect 19663 14768 19708 14796
rect 18785 14759 18843 14765
rect 19702 14756 19708 14768
rect 19760 14756 19766 14808
rect 20162 14756 20168 14808
rect 20220 14796 20226 14808
rect 20257 14799 20315 14805
rect 20257 14796 20269 14799
rect 20220 14768 20269 14796
rect 20220 14756 20226 14768
rect 20257 14765 20269 14768
rect 20303 14765 20315 14799
rect 20257 14759 20315 14765
rect 16853 14731 16911 14737
rect 16853 14697 16865 14731
rect 16899 14728 16911 14731
rect 17402 14728 17408 14740
rect 16899 14700 17408 14728
rect 16899 14697 16911 14700
rect 16853 14691 16911 14697
rect 17402 14688 17408 14700
rect 17460 14688 17466 14740
rect 12345 14663 12403 14669
rect 12345 14660 12357 14663
rect 12124 14632 12357 14660
rect 12124 14620 12130 14632
rect 12345 14629 12357 14632
rect 12391 14629 12403 14663
rect 12345 14623 12403 14629
rect 16485 14663 16543 14669
rect 16485 14629 16497 14663
rect 16531 14629 16543 14663
rect 16942 14660 16948 14672
rect 16903 14632 16948 14660
rect 16485 14623 16543 14629
rect 16942 14620 16948 14632
rect 17000 14620 17006 14672
rect 1104 14570 21620 14592
rect 1104 14518 7846 14570
rect 7898 14518 7910 14570
rect 7962 14518 7974 14570
rect 8026 14518 8038 14570
rect 8090 14518 14710 14570
rect 14762 14518 14774 14570
rect 14826 14518 14838 14570
rect 14890 14518 14902 14570
rect 14954 14518 21620 14570
rect 1104 14496 21620 14518
rect 6822 14416 6828 14468
rect 6880 14456 6886 14468
rect 9769 14459 9827 14465
rect 9769 14456 9781 14459
rect 6880 14428 9781 14456
rect 6880 14416 6886 14428
rect 9769 14425 9781 14428
rect 9815 14456 9827 14459
rect 10226 14456 10232 14468
rect 9815 14428 10232 14456
rect 9815 14425 9827 14428
rect 9769 14419 9827 14425
rect 10226 14416 10232 14428
rect 10284 14416 10290 14468
rect 11974 14416 11980 14468
rect 12032 14456 12038 14468
rect 12897 14459 12955 14465
rect 12897 14456 12909 14459
rect 12032 14428 12909 14456
rect 12032 14416 12038 14428
rect 12897 14425 12909 14428
rect 12943 14425 12955 14459
rect 16853 14459 16911 14465
rect 16853 14456 16865 14459
rect 12897 14419 12955 14425
rect 13648 14428 16865 14456
rect 4148 14391 4206 14397
rect 4148 14357 4160 14391
rect 4194 14388 4206 14391
rect 12250 14388 12256 14400
rect 4194 14360 12256 14388
rect 4194 14357 4206 14360
rect 4148 14351 4206 14357
rect 12250 14348 12256 14360
rect 12308 14388 12314 14400
rect 12308 14360 13032 14388
rect 12308 14348 12314 14360
rect 3878 14320 3884 14332
rect 3839 14292 3884 14320
rect 3878 14280 3884 14292
rect 3936 14280 3942 14332
rect 6086 14320 6092 14332
rect 6047 14292 6092 14320
rect 6086 14280 6092 14292
rect 6144 14280 6150 14332
rect 8662 14329 8668 14332
rect 8656 14320 8668 14329
rect 8623 14292 8668 14320
rect 8656 14283 8668 14292
rect 8662 14280 8668 14283
rect 8720 14280 8726 14332
rect 12618 14280 12624 14332
rect 12676 14320 12682 14332
rect 12805 14323 12863 14329
rect 12805 14320 12817 14323
rect 12676 14292 12817 14320
rect 12676 14280 12682 14292
rect 12805 14289 12817 14292
rect 12851 14289 12863 14323
rect 12805 14283 12863 14289
rect 6178 14252 6184 14264
rect 6139 14224 6184 14252
rect 6178 14212 6184 14224
rect 6236 14212 6242 14264
rect 6270 14212 6276 14264
rect 6328 14252 6334 14264
rect 6328 14224 6373 14252
rect 6328 14212 6334 14224
rect 7374 14212 7380 14264
rect 7432 14252 7438 14264
rect 13004 14261 13032 14360
rect 8389 14255 8447 14261
rect 8389 14252 8401 14255
rect 7432 14224 8401 14252
rect 7432 14212 7438 14224
rect 8389 14221 8401 14224
rect 8435 14221 8447 14255
rect 8389 14215 8447 14221
rect 12989 14255 13047 14261
rect 12989 14221 13001 14255
rect 13035 14221 13047 14255
rect 12989 14215 13047 14221
rect 9950 14144 9956 14196
rect 10008 14184 10014 14196
rect 13648 14184 13676 14428
rect 16853 14425 16865 14428
rect 16899 14456 16911 14459
rect 17034 14456 17040 14468
rect 16899 14428 17040 14456
rect 16899 14425 16911 14428
rect 16853 14419 16911 14425
rect 17034 14416 17040 14428
rect 17092 14416 17098 14468
rect 20898 14456 20904 14468
rect 20859 14428 20904 14456
rect 20898 14416 20904 14428
rect 20956 14416 20962 14468
rect 14084 14391 14142 14397
rect 14084 14357 14096 14391
rect 14130 14388 14142 14391
rect 15194 14388 15200 14400
rect 14130 14360 15200 14388
rect 14130 14357 14142 14360
rect 14084 14351 14142 14357
rect 15194 14348 15200 14360
rect 15252 14348 15258 14400
rect 19521 14391 19579 14397
rect 19521 14357 19533 14391
rect 19567 14388 19579 14391
rect 19567 14360 20760 14388
rect 19567 14357 19579 14360
rect 19521 14351 19579 14357
rect 13814 14320 13820 14332
rect 13775 14292 13820 14320
rect 13814 14280 13820 14292
rect 13872 14320 13878 14332
rect 15289 14323 15347 14329
rect 13872 14292 14872 14320
rect 13872 14280 13878 14292
rect 14844 14252 14872 14292
rect 15289 14289 15301 14323
rect 15335 14320 15347 14323
rect 15740 14323 15798 14329
rect 15740 14320 15752 14323
rect 15335 14292 15752 14320
rect 15335 14289 15347 14292
rect 15289 14283 15347 14289
rect 15740 14289 15752 14292
rect 15786 14320 15798 14323
rect 17034 14320 17040 14332
rect 15786 14292 17040 14320
rect 15786 14289 15798 14292
rect 15740 14283 15798 14289
rect 17034 14280 17040 14292
rect 17092 14280 17098 14332
rect 17126 14280 17132 14332
rect 17184 14320 17190 14332
rect 20732 14329 20760 14360
rect 19245 14323 19303 14329
rect 19245 14320 19257 14323
rect 17184 14292 19257 14320
rect 17184 14280 17190 14292
rect 19245 14289 19257 14292
rect 19291 14289 19303 14323
rect 19981 14323 20039 14329
rect 19981 14320 19993 14323
rect 19245 14283 19303 14289
rect 19352 14292 19993 14320
rect 15473 14255 15531 14261
rect 15473 14252 15485 14255
rect 14844 14224 15485 14252
rect 15473 14221 15485 14224
rect 15519 14221 15531 14255
rect 15473 14215 15531 14221
rect 17313 14255 17371 14261
rect 17313 14221 17325 14255
rect 17359 14252 17371 14255
rect 17770 14252 17776 14264
rect 17359 14224 17776 14252
rect 17359 14221 17371 14224
rect 17313 14215 17371 14221
rect 17770 14212 17776 14224
rect 17828 14212 17834 14264
rect 10008 14156 13676 14184
rect 15197 14187 15255 14193
rect 10008 14144 10014 14156
rect 15197 14153 15209 14187
rect 15243 14184 15255 14187
rect 15289 14187 15347 14193
rect 15289 14184 15301 14187
rect 15243 14156 15301 14184
rect 15243 14153 15255 14156
rect 15197 14147 15255 14153
rect 15289 14153 15301 14156
rect 15335 14153 15347 14187
rect 19352 14184 19380 14292
rect 19981 14289 19993 14292
rect 20027 14289 20039 14323
rect 19981 14283 20039 14289
rect 20717 14323 20775 14329
rect 20717 14289 20729 14323
rect 20763 14289 20775 14323
rect 20717 14283 20775 14289
rect 19702 14212 19708 14264
rect 19760 14252 19766 14264
rect 20165 14255 20223 14261
rect 20165 14252 20177 14255
rect 19760 14224 20177 14252
rect 19760 14212 19766 14224
rect 20165 14221 20177 14224
rect 20211 14221 20223 14255
rect 20165 14215 20223 14221
rect 15289 14147 15347 14153
rect 16776 14156 19380 14184
rect 5261 14119 5319 14125
rect 5261 14085 5273 14119
rect 5307 14116 5319 14119
rect 5534 14116 5540 14128
rect 5307 14088 5540 14116
rect 5307 14085 5319 14088
rect 5261 14079 5319 14085
rect 5534 14076 5540 14088
rect 5592 14076 5598 14128
rect 5721 14119 5779 14125
rect 5721 14085 5733 14119
rect 5767 14116 5779 14119
rect 11698 14116 11704 14128
rect 5767 14088 11704 14116
rect 5767 14085 5779 14088
rect 5721 14079 5779 14085
rect 11698 14076 11704 14088
rect 11756 14076 11762 14128
rect 12437 14119 12495 14125
rect 12437 14085 12449 14119
rect 12483 14116 12495 14119
rect 16776 14116 16804 14156
rect 12483 14088 16804 14116
rect 12483 14085 12495 14088
rect 12437 14079 12495 14085
rect 1104 14026 21620 14048
rect 1104 13974 4414 14026
rect 4466 13974 4478 14026
rect 4530 13974 4542 14026
rect 4594 13974 4606 14026
rect 4658 13974 11278 14026
rect 11330 13974 11342 14026
rect 11394 13974 11406 14026
rect 11458 13974 11470 14026
rect 11522 13974 18142 14026
rect 18194 13974 18206 14026
rect 18258 13974 18270 14026
rect 18322 13974 18334 14026
rect 18386 13974 21620 14026
rect 1104 13952 21620 13974
rect 2498 13872 2504 13924
rect 2556 13912 2562 13924
rect 6270 13912 6276 13924
rect 2556 13884 6276 13912
rect 2556 13872 2562 13884
rect 6270 13872 6276 13884
rect 6328 13872 6334 13924
rect 8202 13872 8208 13924
rect 8260 13872 8266 13924
rect 8662 13912 8668 13924
rect 8623 13884 8668 13912
rect 8662 13872 8668 13884
rect 8720 13872 8726 13924
rect 8941 13915 8999 13921
rect 8941 13912 8953 13915
rect 8772 13884 8953 13912
rect 3602 13844 3608 13856
rect 3563 13816 3608 13844
rect 3602 13804 3608 13816
rect 3660 13804 3666 13856
rect 8220 13844 8248 13872
rect 8772 13844 8800 13884
rect 8941 13881 8953 13884
rect 8987 13881 8999 13915
rect 8941 13875 8999 13881
rect 12250 13872 12256 13924
rect 12308 13912 12314 13924
rect 12345 13915 12403 13921
rect 12345 13912 12357 13915
rect 12308 13884 12357 13912
rect 12308 13872 12314 13884
rect 12345 13881 12357 13884
rect 12391 13881 12403 13915
rect 12618 13912 12624 13924
rect 12579 13884 12624 13912
rect 12345 13875 12403 13881
rect 12618 13872 12624 13884
rect 12676 13872 12682 13924
rect 13449 13915 13507 13921
rect 13449 13881 13461 13915
rect 13495 13912 13507 13915
rect 17402 13912 17408 13924
rect 13495 13884 17264 13912
rect 17363 13884 17408 13912
rect 13495 13881 13507 13884
rect 13449 13875 13507 13881
rect 9950 13844 9956 13856
rect 8220 13816 8800 13844
rect 8956 13816 9956 13844
rect 6086 13736 6092 13788
rect 6144 13776 6150 13788
rect 6549 13779 6607 13785
rect 6549 13776 6561 13779
rect 6144 13748 6561 13776
rect 6144 13736 6150 13748
rect 6549 13745 6561 13748
rect 6595 13745 6607 13779
rect 6549 13739 6607 13745
rect 2225 13711 2283 13717
rect 2225 13677 2237 13711
rect 2271 13708 2283 13711
rect 4893 13711 4951 13717
rect 4893 13708 4905 13711
rect 2271 13680 4905 13708
rect 2271 13677 2283 13680
rect 2225 13671 2283 13677
rect 4893 13677 4905 13680
rect 4939 13708 4951 13711
rect 5160 13711 5218 13717
rect 4939 13680 5120 13708
rect 4939 13677 4951 13680
rect 4893 13671 4951 13677
rect 2498 13649 2504 13652
rect 2492 13603 2504 13649
rect 2556 13640 2562 13652
rect 5092 13640 5120 13680
rect 5160 13677 5172 13711
rect 5206 13708 5218 13711
rect 5534 13708 5540 13720
rect 5206 13680 5540 13708
rect 5206 13677 5218 13680
rect 5160 13671 5218 13677
rect 5534 13668 5540 13680
rect 5592 13708 5598 13720
rect 6270 13708 6276 13720
rect 5592 13680 6276 13708
rect 5592 13668 5598 13680
rect 6270 13668 6276 13680
rect 6328 13668 6334 13720
rect 7285 13711 7343 13717
rect 7285 13708 7297 13711
rect 6380 13680 7297 13708
rect 6380 13640 6408 13680
rect 7285 13677 7297 13680
rect 7331 13708 7343 13711
rect 7374 13708 7380 13720
rect 7331 13680 7380 13708
rect 7331 13677 7343 13680
rect 7285 13671 7343 13677
rect 7374 13668 7380 13680
rect 7432 13668 7438 13720
rect 7552 13711 7610 13717
rect 7552 13677 7564 13711
rect 7598 13708 7610 13711
rect 8956 13708 8984 13816
rect 9950 13804 9956 13816
rect 10008 13804 10014 13856
rect 16393 13847 16451 13853
rect 16393 13813 16405 13847
rect 16439 13844 16451 13847
rect 16942 13844 16948 13856
rect 16439 13816 16948 13844
rect 16439 13813 16451 13816
rect 16393 13807 16451 13813
rect 16942 13804 16948 13816
rect 17000 13804 17006 13856
rect 17236 13844 17264 13884
rect 17402 13872 17408 13884
rect 17460 13872 17466 13924
rect 18598 13912 18604 13924
rect 18559 13884 18604 13912
rect 18598 13872 18604 13884
rect 18656 13872 18662 13924
rect 20441 13915 20499 13921
rect 20441 13881 20453 13915
rect 20487 13912 20499 13915
rect 20622 13912 20628 13924
rect 20487 13884 20628 13912
rect 20487 13881 20499 13884
rect 20441 13875 20499 13881
rect 20622 13872 20628 13884
rect 20680 13872 20686 13924
rect 17862 13844 17868 13856
rect 17236 13816 17868 13844
rect 17862 13804 17868 13816
rect 17920 13804 17926 13856
rect 11974 13736 11980 13788
rect 12032 13776 12038 13788
rect 12342 13776 12348 13788
rect 12032 13748 12348 13776
rect 12032 13736 12038 13748
rect 12342 13736 12348 13748
rect 12400 13776 12406 13788
rect 13173 13779 13231 13785
rect 13173 13776 13185 13779
rect 12400 13748 13185 13776
rect 12400 13736 12406 13748
rect 13173 13745 13185 13748
rect 13219 13745 13231 13779
rect 16850 13776 16856 13788
rect 16811 13748 16856 13776
rect 13173 13739 13231 13745
rect 16850 13736 16856 13748
rect 16908 13736 16914 13788
rect 17034 13776 17040 13788
rect 16947 13748 17040 13776
rect 17034 13736 17040 13748
rect 17092 13776 17098 13788
rect 17957 13779 18015 13785
rect 17957 13776 17969 13779
rect 17092 13748 17969 13776
rect 17092 13736 17098 13748
rect 17957 13745 17969 13748
rect 18003 13745 18015 13779
rect 17957 13739 18015 13745
rect 20346 13736 20352 13788
rect 20404 13776 20410 13788
rect 20622 13776 20628 13788
rect 20404 13748 20628 13776
rect 20404 13736 20410 13748
rect 20622 13736 20628 13748
rect 20680 13736 20686 13788
rect 7598 13680 8984 13708
rect 9125 13711 9183 13717
rect 7598 13677 7610 13680
rect 7552 13671 7610 13677
rect 9125 13677 9137 13711
rect 9171 13708 9183 13711
rect 10870 13708 10876 13720
rect 9171 13680 10876 13708
rect 9171 13677 9183 13680
rect 9125 13671 9183 13677
rect 10870 13668 10876 13680
rect 10928 13668 10934 13720
rect 10962 13668 10968 13720
rect 11020 13708 11026 13720
rect 11020 13680 11065 13708
rect 11020 13668 11026 13680
rect 11698 13668 11704 13720
rect 11756 13708 11762 13720
rect 17126 13708 17132 13720
rect 11756 13680 17132 13708
rect 11756 13668 11762 13680
rect 17126 13668 17132 13680
rect 17184 13668 17190 13720
rect 17862 13708 17868 13720
rect 17823 13680 17868 13708
rect 17862 13668 17868 13680
rect 17920 13668 17926 13720
rect 18414 13708 18420 13720
rect 18375 13680 18420 13708
rect 18414 13668 18420 13680
rect 18472 13668 18478 13720
rect 20254 13708 20260 13720
rect 20215 13680 20260 13708
rect 20254 13668 20260 13680
rect 20312 13668 20318 13720
rect 2556 13612 2592 13640
rect 5092 13612 6408 13640
rect 2498 13600 2504 13603
rect 2556 13600 2562 13612
rect 11146 13600 11152 13652
rect 11204 13649 11210 13652
rect 11204 13643 11268 13649
rect 11204 13609 11222 13643
rect 11256 13640 11268 13643
rect 11974 13640 11980 13652
rect 11256 13612 11980 13640
rect 11256 13609 11268 13612
rect 11204 13603 11268 13609
rect 11204 13600 11210 13603
rect 11974 13600 11980 13612
rect 12032 13600 12038 13652
rect 12989 13643 13047 13649
rect 12989 13609 13001 13643
rect 13035 13640 13047 13643
rect 13633 13643 13691 13649
rect 13633 13640 13645 13643
rect 13035 13612 13645 13640
rect 13035 13609 13047 13612
rect 12989 13603 13047 13609
rect 13633 13609 13645 13612
rect 13679 13609 13691 13643
rect 17770 13640 17776 13652
rect 17731 13612 17776 13640
rect 13633 13603 13691 13609
rect 17770 13600 17776 13612
rect 17828 13600 17834 13652
rect 13081 13575 13139 13581
rect 13081 13541 13093 13575
rect 13127 13572 13139 13575
rect 13449 13575 13507 13581
rect 13449 13572 13461 13575
rect 13127 13544 13461 13572
rect 13127 13541 13139 13544
rect 13081 13535 13139 13541
rect 13449 13541 13461 13544
rect 13495 13541 13507 13575
rect 16758 13572 16764 13584
rect 16719 13544 16764 13572
rect 13449 13535 13507 13541
rect 16758 13532 16764 13544
rect 16816 13532 16822 13584
rect 1104 13482 21620 13504
rect 1104 13430 7846 13482
rect 7898 13430 7910 13482
rect 7962 13430 7974 13482
rect 8026 13430 8038 13482
rect 8090 13430 14710 13482
rect 14762 13430 14774 13482
rect 14826 13430 14838 13482
rect 14890 13430 14902 13482
rect 14954 13430 21620 13482
rect 1104 13408 21620 13430
rect 5629 13371 5687 13377
rect 5629 13337 5641 13371
rect 5675 13368 5687 13371
rect 6178 13368 6184 13380
rect 5675 13340 6184 13368
rect 5675 13337 5687 13340
rect 5629 13331 5687 13337
rect 6178 13328 6184 13340
rect 6236 13328 6242 13380
rect 10870 13328 10876 13380
rect 10928 13368 10934 13380
rect 11333 13371 11391 13377
rect 11333 13368 11345 13371
rect 10928 13340 11345 13368
rect 10928 13328 10934 13340
rect 11333 13337 11345 13340
rect 11379 13368 11391 13371
rect 12253 13371 12311 13377
rect 12253 13368 12265 13371
rect 11379 13340 12265 13368
rect 11379 13337 11391 13340
rect 11333 13331 11391 13337
rect 12253 13337 12265 13340
rect 12299 13337 12311 13371
rect 12253 13331 12311 13337
rect 19518 13328 19524 13380
rect 19576 13368 19582 13380
rect 19613 13371 19671 13377
rect 19613 13368 19625 13371
rect 19576 13340 19625 13368
rect 19576 13328 19582 13340
rect 19613 13337 19625 13340
rect 19659 13337 19671 13371
rect 20162 13368 20168 13380
rect 20123 13340 20168 13368
rect 19613 13331 19671 13337
rect 20162 13328 20168 13340
rect 20220 13328 20226 13380
rect 20714 13368 20720 13380
rect 20675 13340 20720 13368
rect 20714 13328 20720 13340
rect 20772 13328 20778 13380
rect 5902 13260 5908 13312
rect 5960 13300 5966 13312
rect 6089 13303 6147 13309
rect 6089 13300 6101 13303
rect 5960 13272 6101 13300
rect 5960 13260 5966 13272
rect 6089 13269 6101 13272
rect 6135 13269 6147 13303
rect 6089 13263 6147 13269
rect 10042 13260 10048 13312
rect 10100 13300 10106 13312
rect 10100 13272 10145 13300
rect 10100 13260 10106 13272
rect 18414 13260 18420 13312
rect 18472 13300 18478 13312
rect 18969 13303 19027 13309
rect 18969 13300 18981 13303
rect 18472 13272 18981 13300
rect 18472 13260 18478 13272
rect 18969 13269 18981 13272
rect 19015 13269 19027 13303
rect 18969 13263 19027 13269
rect 5997 13235 6055 13241
rect 5997 13201 6009 13235
rect 6043 13232 6055 13235
rect 8386 13232 8392 13244
rect 6043 13204 8392 13232
rect 6043 13201 6055 13204
rect 5997 13195 6055 13201
rect 8386 13192 8392 13204
rect 8444 13192 8450 13244
rect 8478 13192 8484 13244
rect 8536 13232 8542 13244
rect 14458 13232 14464 13244
rect 8536 13204 14464 13232
rect 8536 13192 8542 13204
rect 14458 13192 14464 13204
rect 14516 13192 14522 13244
rect 18690 13232 18696 13244
rect 18651 13204 18696 13232
rect 18690 13192 18696 13204
rect 18748 13192 18754 13244
rect 19242 13192 19248 13244
rect 19300 13232 19306 13244
rect 19429 13235 19487 13241
rect 19429 13232 19441 13235
rect 19300 13204 19441 13232
rect 19300 13192 19306 13204
rect 19429 13201 19441 13204
rect 19475 13201 19487 13235
rect 19429 13195 19487 13201
rect 19981 13235 20039 13241
rect 19981 13201 19993 13235
rect 20027 13201 20039 13235
rect 20530 13232 20536 13244
rect 20491 13204 20536 13232
rect 19981 13195 20039 13201
rect 6270 13164 6276 13176
rect 6231 13136 6276 13164
rect 6270 13124 6276 13136
rect 6328 13124 6334 13176
rect 11698 13124 11704 13176
rect 11756 13164 11762 13176
rect 19996 13164 20024 13195
rect 20530 13192 20536 13204
rect 20588 13192 20594 13244
rect 11756 13136 20024 13164
rect 11756 13124 11762 13136
rect 12253 13099 12311 13105
rect 12253 13065 12265 13099
rect 12299 13096 12311 13099
rect 12618 13096 12624 13108
rect 12299 13068 12624 13096
rect 12299 13065 12311 13068
rect 12253 13059 12311 13065
rect 12618 13056 12624 13068
rect 12676 13056 12682 13108
rect 842 12988 848 13040
rect 900 13028 906 13040
rect 13446 13028 13452 13040
rect 900 13000 13452 13028
rect 900 12988 906 13000
rect 13446 12988 13452 13000
rect 13504 12988 13510 13040
rect 1104 12938 21620 12960
rect 1104 12886 4414 12938
rect 4466 12886 4478 12938
rect 4530 12886 4542 12938
rect 4594 12886 4606 12938
rect 4658 12886 11278 12938
rect 11330 12886 11342 12938
rect 11394 12886 11406 12938
rect 11458 12886 11470 12938
rect 11522 12886 18142 12938
rect 18194 12886 18206 12938
rect 18258 12886 18270 12938
rect 18322 12886 18334 12938
rect 18386 12886 21620 12938
rect 1104 12864 21620 12886
rect 7374 12784 7380 12836
rect 7432 12824 7438 12836
rect 7558 12824 7564 12836
rect 7432 12796 7564 12824
rect 7432 12784 7438 12796
rect 7558 12784 7564 12796
rect 7616 12784 7622 12836
rect 8386 12784 8392 12836
rect 8444 12824 8450 12836
rect 8444 12796 11100 12824
rect 8444 12784 8450 12796
rect 7558 12648 7564 12700
rect 7616 12688 7622 12700
rect 9953 12691 10011 12697
rect 9953 12688 9965 12691
rect 7616 12660 9965 12688
rect 7616 12648 7622 12660
rect 9953 12657 9965 12660
rect 9999 12657 10011 12691
rect 9953 12651 10011 12657
rect 7745 12623 7803 12629
rect 7745 12589 7757 12623
rect 7791 12620 7803 12623
rect 8202 12620 8208 12632
rect 7791 12592 8208 12620
rect 7791 12589 7803 12592
rect 7745 12583 7803 12589
rect 8202 12580 8208 12592
rect 8260 12580 8266 12632
rect 10226 12561 10232 12564
rect 10220 12515 10232 12561
rect 10284 12552 10290 12564
rect 10284 12524 10320 12552
rect 10226 12512 10232 12515
rect 10284 12512 10290 12524
rect 11072 12484 11100 12796
rect 11146 12784 11152 12836
rect 11204 12824 11210 12836
rect 11333 12827 11391 12833
rect 11333 12824 11345 12827
rect 11204 12796 11345 12824
rect 11204 12784 11210 12796
rect 11333 12793 11345 12796
rect 11379 12793 11391 12827
rect 11333 12787 11391 12793
rect 12437 12827 12495 12833
rect 12437 12793 12449 12827
rect 12483 12824 12495 12827
rect 13354 12824 13360 12836
rect 12483 12796 13360 12824
rect 12483 12793 12495 12796
rect 12437 12787 12495 12793
rect 13354 12784 13360 12796
rect 13412 12784 13418 12836
rect 20162 12824 20168 12836
rect 20123 12796 20168 12824
rect 20162 12784 20168 12796
rect 20220 12784 20226 12836
rect 12989 12759 13047 12765
rect 12989 12725 13001 12759
rect 13035 12756 13047 12759
rect 14550 12756 14556 12768
rect 13035 12728 14556 12756
rect 13035 12725 13047 12728
rect 12989 12719 13047 12725
rect 14550 12716 14556 12728
rect 14608 12716 14614 12768
rect 11698 12688 11704 12700
rect 11659 12660 11704 12688
rect 11698 12648 11704 12660
rect 11756 12648 11762 12700
rect 13446 12688 13452 12700
rect 13407 12660 13452 12688
rect 13446 12648 13452 12660
rect 13504 12648 13510 12700
rect 13538 12648 13544 12700
rect 13596 12688 13602 12700
rect 13633 12691 13691 12697
rect 13633 12688 13645 12691
rect 13596 12660 13645 12688
rect 13596 12648 13602 12660
rect 13633 12657 13645 12660
rect 13679 12688 13691 12691
rect 14645 12691 14703 12697
rect 14645 12688 14657 12691
rect 13679 12660 14657 12688
rect 13679 12657 13691 12660
rect 13633 12651 13691 12657
rect 14645 12657 14657 12660
rect 14691 12688 14703 12691
rect 15102 12688 15108 12700
rect 14691 12660 15108 12688
rect 14691 12657 14703 12660
rect 14645 12651 14703 12657
rect 15102 12648 15108 12660
rect 15160 12648 15166 12700
rect 15194 12648 15200 12700
rect 15252 12688 15258 12700
rect 16577 12691 16635 12697
rect 16577 12688 16589 12691
rect 15252 12660 16589 12688
rect 15252 12648 15258 12660
rect 16577 12657 16589 12660
rect 16623 12657 16635 12691
rect 20530 12688 20536 12700
rect 16577 12651 16635 12657
rect 18064 12660 20536 12688
rect 11422 12620 11428 12632
rect 11383 12592 11428 12620
rect 11422 12580 11428 12592
rect 11480 12580 11486 12632
rect 12618 12580 12624 12632
rect 12676 12629 12682 12632
rect 12676 12620 12687 12629
rect 12676 12592 12721 12620
rect 12676 12583 12687 12592
rect 12676 12580 12682 12583
rect 13814 12580 13820 12632
rect 13872 12620 13878 12632
rect 15289 12623 15347 12629
rect 15289 12620 15301 12623
rect 13872 12592 15301 12620
rect 13872 12580 13878 12592
rect 15289 12589 15301 12592
rect 15335 12589 15347 12623
rect 15289 12583 15347 12589
rect 15565 12623 15623 12629
rect 15565 12589 15577 12623
rect 15611 12620 15623 12623
rect 18064 12620 18092 12660
rect 20530 12648 20536 12660
rect 20588 12648 20594 12700
rect 19150 12620 19156 12632
rect 15611 12592 18092 12620
rect 19111 12592 19156 12620
rect 15611 12589 15623 12592
rect 15565 12583 15623 12589
rect 19150 12580 19156 12592
rect 19208 12580 19214 12632
rect 19429 12623 19487 12629
rect 19429 12589 19441 12623
rect 19475 12620 19487 12623
rect 19981 12623 20039 12629
rect 19981 12620 19993 12623
rect 19475 12592 19993 12620
rect 19475 12589 19487 12592
rect 19429 12583 19487 12589
rect 19981 12589 19993 12592
rect 20027 12589 20039 12623
rect 19981 12583 20039 12589
rect 14458 12552 14464 12564
rect 14419 12524 14464 12552
rect 14458 12512 14464 12524
rect 14516 12512 14522 12564
rect 16844 12555 16902 12561
rect 16844 12521 16856 12555
rect 16890 12552 16902 12555
rect 17494 12552 17500 12564
rect 16890 12524 17500 12552
rect 16890 12521 16902 12524
rect 16844 12515 16902 12521
rect 17494 12512 17500 12524
rect 17552 12512 17558 12564
rect 13357 12487 13415 12493
rect 13357 12484 13369 12487
rect 11072 12456 13369 12484
rect 13357 12453 13369 12456
rect 13403 12484 13415 12487
rect 13446 12484 13452 12496
rect 13403 12456 13452 12484
rect 13403 12453 13415 12456
rect 13357 12447 13415 12453
rect 13446 12444 13452 12456
rect 13504 12444 13510 12496
rect 13998 12484 14004 12496
rect 13959 12456 14004 12484
rect 13998 12444 14004 12456
rect 14056 12444 14062 12496
rect 14182 12444 14188 12496
rect 14240 12484 14246 12496
rect 14369 12487 14427 12493
rect 14369 12484 14381 12487
rect 14240 12456 14381 12484
rect 14240 12444 14246 12456
rect 14369 12453 14381 12456
rect 14415 12453 14427 12487
rect 17954 12484 17960 12496
rect 17915 12456 17960 12484
rect 14369 12447 14427 12453
rect 17954 12444 17960 12456
rect 18012 12444 18018 12496
rect 1104 12394 21620 12416
rect 1104 12342 7846 12394
rect 7898 12342 7910 12394
rect 7962 12342 7974 12394
rect 8026 12342 8038 12394
rect 8090 12342 14710 12394
rect 14762 12342 14774 12394
rect 14826 12342 14838 12394
rect 14890 12342 14902 12394
rect 14954 12342 21620 12394
rect 1104 12320 21620 12342
rect 8938 12240 8944 12292
rect 8996 12240 9002 12292
rect 10413 12283 10471 12289
rect 10413 12249 10425 12283
rect 10459 12280 10471 12283
rect 11422 12280 11428 12292
rect 10459 12252 11428 12280
rect 10459 12249 10471 12252
rect 10413 12243 10471 12249
rect 11422 12240 11428 12252
rect 11480 12240 11486 12292
rect 14182 12280 14188 12292
rect 12636 12252 14188 12280
rect 7190 12212 7196 12224
rect 7024 12184 7196 12212
rect 7024 12153 7052 12184
rect 7190 12172 7196 12184
rect 7248 12212 7254 12224
rect 7558 12212 7564 12224
rect 7248 12184 7564 12212
rect 7248 12172 7254 12184
rect 7558 12172 7564 12184
rect 7616 12212 7622 12224
rect 8956 12212 8984 12240
rect 12636 12212 12664 12252
rect 14182 12240 14188 12252
rect 14240 12240 14246 12292
rect 14550 12280 14556 12292
rect 14511 12252 14556 12280
rect 14550 12240 14556 12252
rect 14608 12240 14614 12292
rect 15102 12240 15108 12292
rect 15160 12280 15166 12292
rect 16577 12283 16635 12289
rect 16577 12280 16589 12283
rect 15160 12252 16589 12280
rect 15160 12240 15166 12252
rect 16577 12249 16589 12252
rect 16623 12249 16635 12283
rect 16577 12243 16635 12249
rect 17954 12240 17960 12292
rect 18012 12240 18018 12292
rect 18049 12283 18107 12289
rect 18049 12249 18061 12283
rect 18095 12280 18107 12283
rect 19150 12280 19156 12292
rect 18095 12252 19156 12280
rect 18095 12249 18107 12252
rect 18049 12243 18107 12249
rect 19150 12240 19156 12252
rect 19208 12240 19214 12292
rect 20165 12283 20223 12289
rect 20165 12249 20177 12283
rect 20211 12280 20223 12283
rect 20990 12280 20996 12292
rect 20211 12252 20996 12280
rect 20211 12249 20223 12252
rect 20165 12243 20223 12249
rect 20990 12240 20996 12252
rect 21048 12240 21054 12292
rect 7616 12184 8800 12212
rect 8956 12184 12664 12212
rect 12704 12215 12762 12221
rect 7616 12172 7622 12184
rect 7282 12153 7288 12156
rect 7009 12147 7067 12153
rect 7009 12113 7021 12147
rect 7055 12113 7067 12147
rect 7009 12107 7067 12113
rect 7276 12107 7288 12153
rect 7340 12144 7346 12156
rect 8772 12153 8800 12184
rect 12704 12181 12716 12215
rect 12750 12212 12762 12215
rect 13538 12212 13544 12224
rect 12750 12184 13544 12212
rect 12750 12181 12762 12184
rect 12704 12175 12762 12181
rect 13538 12172 13544 12184
rect 13596 12172 13602 12224
rect 13998 12172 14004 12224
rect 14056 12212 14062 12224
rect 14461 12215 14519 12221
rect 14461 12212 14473 12215
rect 14056 12184 14473 12212
rect 14056 12172 14062 12184
rect 14461 12181 14473 12184
rect 14507 12181 14519 12215
rect 14461 12175 14519 12181
rect 15464 12215 15522 12221
rect 15464 12181 15476 12215
rect 15510 12212 15522 12215
rect 17972 12212 18000 12240
rect 15510 12184 18552 12212
rect 15510 12181 15522 12184
rect 15464 12175 15522 12181
rect 8757 12147 8815 12153
rect 7340 12116 7376 12144
rect 7282 12104 7288 12107
rect 7340 12104 7346 12116
rect 8757 12113 8769 12147
rect 8803 12113 8815 12147
rect 9013 12147 9071 12153
rect 9013 12144 9025 12147
rect 8757 12107 8815 12113
rect 8864 12116 9025 12144
rect 8864 12076 8892 12116
rect 9013 12113 9025 12116
rect 9059 12113 9071 12147
rect 9013 12107 9071 12113
rect 10410 12104 10416 12156
rect 10468 12144 10474 12156
rect 10781 12147 10839 12153
rect 10781 12144 10793 12147
rect 10468 12116 10793 12144
rect 10468 12104 10474 12116
rect 10781 12113 10793 12116
rect 10827 12113 10839 12147
rect 15194 12144 15200 12156
rect 10781 12107 10839 12113
rect 12452 12116 15200 12144
rect 12452 12088 12480 12116
rect 15194 12104 15200 12116
rect 15252 12104 15258 12156
rect 17954 12104 17960 12156
rect 18012 12144 18018 12156
rect 18417 12147 18475 12153
rect 18417 12144 18429 12147
rect 18012 12116 18429 12144
rect 18012 12104 18018 12116
rect 18417 12113 18429 12116
rect 18463 12113 18475 12147
rect 18524 12144 18552 12184
rect 19978 12144 19984 12156
rect 18524 12116 18644 12144
rect 19939 12116 19984 12144
rect 18417 12107 18475 12113
rect 8680 12048 8892 12076
rect 8680 11952 8708 12048
rect 9766 12036 9772 12088
rect 9824 12076 9830 12088
rect 10873 12079 10931 12085
rect 10873 12076 10885 12079
rect 9824 12048 10885 12076
rect 9824 12036 9830 12048
rect 10873 12045 10885 12048
rect 10919 12045 10931 12079
rect 10873 12039 10931 12045
rect 10965 12079 11023 12085
rect 10965 12045 10977 12079
rect 11011 12045 11023 12079
rect 10965 12039 11023 12045
rect 10137 12011 10195 12017
rect 10137 11977 10149 12011
rect 10183 12008 10195 12011
rect 10226 12008 10232 12020
rect 10183 11980 10232 12008
rect 10183 11977 10195 11980
rect 10137 11971 10195 11977
rect 10226 11968 10232 11980
rect 10284 12008 10290 12020
rect 10980 12008 11008 12039
rect 12434 12036 12440 12088
rect 12492 12076 12498 12088
rect 14645 12079 14703 12085
rect 14645 12076 14657 12079
rect 12492 12048 12537 12076
rect 14292 12048 14657 12076
rect 12492 12036 12498 12048
rect 14292 12020 14320 12048
rect 14645 12045 14657 12048
rect 14691 12045 14703 12079
rect 14645 12039 14703 12045
rect 16942 12036 16948 12088
rect 17000 12076 17006 12088
rect 18616 12085 18644 12116
rect 19978 12104 19984 12116
rect 20036 12104 20042 12156
rect 20530 12144 20536 12156
rect 20491 12116 20536 12144
rect 20530 12104 20536 12116
rect 20588 12104 20594 12156
rect 18509 12079 18567 12085
rect 18509 12076 18521 12079
rect 17000 12048 18521 12076
rect 17000 12036 17006 12048
rect 18509 12045 18521 12048
rect 18555 12045 18567 12079
rect 18509 12039 18567 12045
rect 18601 12079 18659 12085
rect 18601 12045 18613 12079
rect 18647 12045 18659 12079
rect 18601 12039 18659 12045
rect 10284 11980 11008 12008
rect 13817 12011 13875 12017
rect 10284 11968 10290 11980
rect 13817 11977 13829 12011
rect 13863 12008 13875 12011
rect 14274 12008 14280 12020
rect 13863 11980 14280 12008
rect 13863 11977 13875 11980
rect 13817 11971 13875 11977
rect 14274 11968 14280 11980
rect 14332 11968 14338 12020
rect 19610 11968 19616 12020
rect 19668 12008 19674 12020
rect 20717 12011 20775 12017
rect 20717 12008 20729 12011
rect 19668 11980 20729 12008
rect 19668 11968 19674 11980
rect 20717 11977 20729 11980
rect 20763 11977 20775 12011
rect 20717 11971 20775 11977
rect 8389 11943 8447 11949
rect 8389 11909 8401 11943
rect 8435 11940 8447 11943
rect 8662 11940 8668 11952
rect 8435 11912 8668 11940
rect 8435 11909 8447 11912
rect 8389 11903 8447 11909
rect 8662 11900 8668 11912
rect 8720 11900 8726 11952
rect 13998 11900 14004 11952
rect 14056 11940 14062 11952
rect 14093 11943 14151 11949
rect 14093 11940 14105 11943
rect 14056 11912 14105 11940
rect 14056 11900 14062 11912
rect 14093 11909 14105 11912
rect 14139 11909 14151 11943
rect 14093 11903 14151 11909
rect 14182 11900 14188 11952
rect 14240 11940 14246 11952
rect 18598 11940 18604 11952
rect 14240 11912 18604 11940
rect 14240 11900 14246 11912
rect 18598 11900 18604 11912
rect 18656 11900 18662 11952
rect 1104 11850 21620 11872
rect 1104 11798 4414 11850
rect 4466 11798 4478 11850
rect 4530 11798 4542 11850
rect 4594 11798 4606 11850
rect 4658 11798 11278 11850
rect 11330 11798 11342 11850
rect 11394 11798 11406 11850
rect 11458 11798 11470 11850
rect 11522 11798 18142 11850
rect 18194 11798 18206 11850
rect 18258 11798 18270 11850
rect 18322 11798 18334 11850
rect 18386 11798 21620 11850
rect 1104 11776 21620 11798
rect 8021 11739 8079 11745
rect 8021 11705 8033 11739
rect 8067 11736 8079 11739
rect 9766 11736 9772 11748
rect 8067 11708 9772 11736
rect 8067 11705 8079 11708
rect 8021 11699 8079 11705
rect 9766 11696 9772 11708
rect 9824 11696 9830 11748
rect 10410 11736 10416 11748
rect 10371 11708 10416 11736
rect 10410 11696 10416 11708
rect 10468 11696 10474 11748
rect 12434 11696 12440 11748
rect 12492 11736 12498 11748
rect 13265 11739 13323 11745
rect 13265 11736 13277 11739
rect 12492 11708 13277 11736
rect 12492 11696 12498 11708
rect 13265 11705 13277 11708
rect 13311 11705 13323 11739
rect 13265 11699 13323 11705
rect 13541 11739 13599 11745
rect 13541 11705 13553 11739
rect 13587 11736 13599 11739
rect 13814 11736 13820 11748
rect 13587 11708 13820 11736
rect 13587 11705 13599 11708
rect 13541 11699 13599 11705
rect 13814 11696 13820 11708
rect 13872 11696 13878 11748
rect 17954 11696 17960 11748
rect 18012 11736 18018 11748
rect 18049 11739 18107 11745
rect 18049 11736 18061 11739
rect 18012 11708 18061 11736
rect 18012 11696 18018 11708
rect 18049 11705 18061 11708
rect 18095 11705 18107 11739
rect 18049 11699 18107 11705
rect 20070 11696 20076 11748
rect 20128 11736 20134 11748
rect 20441 11739 20499 11745
rect 20441 11736 20453 11739
rect 20128 11708 20453 11736
rect 20128 11696 20134 11708
rect 20441 11705 20453 11708
rect 20487 11705 20499 11739
rect 20441 11699 20499 11705
rect 14366 11668 14372 11680
rect 10888 11640 14372 11668
rect 6822 11560 6828 11612
rect 6880 11600 6886 11612
rect 7193 11603 7251 11609
rect 7193 11600 7205 11603
rect 6880 11572 7205 11600
rect 6880 11560 6886 11572
rect 7193 11569 7205 11572
rect 7239 11569 7251 11603
rect 7193 11563 7251 11569
rect 7282 11560 7288 11612
rect 7340 11600 7346 11612
rect 8662 11600 8668 11612
rect 7340 11572 8524 11600
rect 8575 11572 8668 11600
rect 7340 11560 7346 11572
rect 7101 11535 7159 11541
rect 7101 11501 7113 11535
rect 7147 11532 7159 11535
rect 8386 11532 8392 11544
rect 7147 11504 8392 11532
rect 7147 11501 7159 11504
rect 7101 11495 7159 11501
rect 8386 11492 8392 11504
rect 8444 11492 8450 11544
rect 8496 11532 8524 11572
rect 8662 11560 8668 11572
rect 8720 11560 8726 11612
rect 10888 11609 10916 11640
rect 14366 11628 14372 11640
rect 14424 11628 14430 11680
rect 10873 11603 10931 11609
rect 10873 11569 10885 11603
rect 10919 11569 10931 11603
rect 10873 11563 10931 11569
rect 10965 11603 11023 11609
rect 10965 11569 10977 11603
rect 11011 11569 11023 11603
rect 13998 11600 14004 11612
rect 13959 11572 14004 11600
rect 10965 11563 11023 11569
rect 8570 11532 8576 11544
rect 8496 11504 8576 11532
rect 8570 11492 8576 11504
rect 8628 11492 8634 11544
rect 8680 11532 8708 11560
rect 10980 11532 11008 11563
rect 13998 11560 14004 11572
rect 14056 11560 14062 11612
rect 14090 11560 14096 11612
rect 14148 11600 14154 11612
rect 14148 11572 14193 11600
rect 14148 11560 14154 11572
rect 17494 11560 17500 11612
rect 17552 11600 17558 11612
rect 18601 11603 18659 11609
rect 18601 11600 18613 11603
rect 17552 11572 18613 11600
rect 17552 11560 17558 11572
rect 18601 11569 18613 11572
rect 18647 11569 18659 11603
rect 18601 11563 18659 11569
rect 8680 11504 11008 11532
rect 13354 11492 13360 11544
rect 13412 11532 13418 11544
rect 13449 11535 13507 11541
rect 13449 11532 13461 11535
rect 13412 11504 13461 11532
rect 13412 11492 13418 11504
rect 13449 11501 13461 11504
rect 13495 11501 13507 11535
rect 13449 11495 13507 11501
rect 15746 11492 15752 11544
rect 15804 11532 15810 11544
rect 19150 11532 19156 11544
rect 15804 11504 19156 11532
rect 15804 11492 15810 11504
rect 19150 11492 19156 11504
rect 19208 11492 19214 11544
rect 20254 11532 20260 11544
rect 20215 11504 20260 11532
rect 20254 11492 20260 11504
rect 20312 11492 20318 11544
rect 8481 11467 8539 11473
rect 8481 11464 8493 11467
rect 6748 11436 8493 11464
rect 6748 11405 6776 11436
rect 8481 11433 8493 11436
rect 8527 11433 8539 11467
rect 8481 11427 8539 11433
rect 10781 11467 10839 11473
rect 10781 11433 10793 11467
rect 10827 11464 10839 11467
rect 11425 11467 11483 11473
rect 11425 11464 11437 11467
rect 10827 11436 11437 11464
rect 10827 11433 10839 11436
rect 10781 11427 10839 11433
rect 11425 11433 11437 11436
rect 11471 11433 11483 11467
rect 11425 11427 11483 11433
rect 11606 11424 11612 11476
rect 11664 11464 11670 11476
rect 14550 11464 14556 11476
rect 11664 11436 14556 11464
rect 11664 11424 11670 11436
rect 14550 11424 14556 11436
rect 14608 11424 14614 11476
rect 18417 11467 18475 11473
rect 18417 11433 18429 11467
rect 18463 11464 18475 11467
rect 19061 11467 19119 11473
rect 19061 11464 19073 11467
rect 18463 11436 19073 11464
rect 18463 11433 18475 11436
rect 18417 11427 18475 11433
rect 19061 11433 19073 11436
rect 19107 11433 19119 11467
rect 19061 11427 19119 11433
rect 6733 11399 6791 11405
rect 6733 11365 6745 11399
rect 6779 11365 6791 11399
rect 6733 11359 6791 11365
rect 8294 11356 8300 11408
rect 8352 11396 8358 11408
rect 8389 11399 8447 11405
rect 8389 11396 8401 11399
rect 8352 11368 8401 11396
rect 8352 11356 8358 11368
rect 8389 11365 8401 11368
rect 8435 11365 8447 11399
rect 8389 11359 8447 11365
rect 13722 11356 13728 11408
rect 13780 11396 13786 11408
rect 13909 11399 13967 11405
rect 13909 11396 13921 11399
rect 13780 11368 13921 11396
rect 13780 11356 13786 11368
rect 13909 11365 13921 11368
rect 13955 11365 13967 11399
rect 13909 11359 13967 11365
rect 18509 11399 18567 11405
rect 18509 11365 18521 11399
rect 18555 11396 18567 11399
rect 18782 11396 18788 11408
rect 18555 11368 18788 11396
rect 18555 11365 18567 11368
rect 18509 11359 18567 11365
rect 18782 11356 18788 11368
rect 18840 11356 18846 11408
rect 1104 11306 21620 11328
rect 1104 11254 7846 11306
rect 7898 11254 7910 11306
rect 7962 11254 7974 11306
rect 8026 11254 8038 11306
rect 8090 11254 14710 11306
rect 14762 11254 14774 11306
rect 14826 11254 14838 11306
rect 14890 11254 14902 11306
rect 14954 11254 21620 11306
rect 1104 11232 21620 11254
rect 8294 11192 8300 11204
rect 8255 11164 8300 11192
rect 8294 11152 8300 11164
rect 8352 11152 8358 11204
rect 8478 11152 8484 11204
rect 8536 11192 8542 11204
rect 8757 11195 8815 11201
rect 8757 11192 8769 11195
rect 8536 11164 8769 11192
rect 8536 11152 8542 11164
rect 8757 11161 8769 11164
rect 8803 11161 8815 11195
rect 13722 11192 13728 11204
rect 13683 11164 13728 11192
rect 8757 11155 8815 11161
rect 13722 11152 13728 11164
rect 13780 11152 13786 11204
rect 14182 11152 14188 11204
rect 14240 11192 14246 11204
rect 14366 11192 14372 11204
rect 14240 11164 14372 11192
rect 14240 11152 14246 11164
rect 14366 11152 14372 11164
rect 14424 11152 14430 11204
rect 15933 11195 15991 11201
rect 15933 11161 15945 11195
rect 15979 11192 15991 11195
rect 17405 11195 17463 11201
rect 17405 11192 17417 11195
rect 15979 11164 17417 11192
rect 15979 11161 15991 11164
rect 15933 11155 15991 11161
rect 17405 11161 17417 11164
rect 17451 11161 17463 11195
rect 18782 11192 18788 11204
rect 18743 11164 18788 11192
rect 17405 11155 17463 11161
rect 18782 11152 18788 11164
rect 18840 11152 18846 11204
rect 20165 11195 20223 11201
rect 20165 11161 20177 11195
rect 20211 11192 20223 11195
rect 20622 11192 20628 11204
rect 20211 11164 20628 11192
rect 20211 11161 20223 11164
rect 20165 11155 20223 11161
rect 20622 11152 20628 11164
rect 20680 11152 20686 11204
rect 20717 11195 20775 11201
rect 20717 11161 20729 11195
rect 20763 11192 20775 11195
rect 20806 11192 20812 11204
rect 20763 11164 20812 11192
rect 20763 11161 20775 11164
rect 20717 11155 20775 11161
rect 20806 11152 20812 11164
rect 20864 11152 20870 11204
rect 8665 11127 8723 11133
rect 8665 11093 8677 11127
rect 8711 11124 8723 11127
rect 8938 11124 8944 11136
rect 8711 11096 8944 11124
rect 8711 11093 8723 11096
rect 8665 11087 8723 11093
rect 8938 11084 8944 11096
rect 8996 11084 9002 11136
rect 10965 11127 11023 11133
rect 10965 11093 10977 11127
rect 11011 11124 11023 11127
rect 11011 11096 20576 11124
rect 11011 11093 11023 11096
rect 10965 11087 11023 11093
rect 10042 11016 10048 11068
rect 10100 11056 10106 11068
rect 10689 11059 10747 11065
rect 10689 11056 10701 11059
rect 10100 11028 10701 11056
rect 10100 11016 10106 11028
rect 10689 11025 10701 11028
rect 10735 11025 10747 11059
rect 10689 11019 10747 11025
rect 14093 11059 14151 11065
rect 14093 11025 14105 11059
rect 14139 11056 14151 11059
rect 14737 11059 14795 11065
rect 14737 11056 14749 11059
rect 14139 11028 14749 11056
rect 14139 11025 14151 11028
rect 14093 11019 14151 11025
rect 14737 11025 14749 11028
rect 14783 11025 14795 11059
rect 14737 11019 14795 11025
rect 15749 11059 15807 11065
rect 15749 11025 15761 11059
rect 15795 11056 15807 11059
rect 16301 11059 16359 11065
rect 16301 11056 16313 11059
rect 15795 11028 16313 11056
rect 15795 11025 15807 11028
rect 15749 11019 15807 11025
rect 16301 11025 16313 11028
rect 16347 11056 16359 11059
rect 16758 11056 16764 11068
rect 16347 11028 16764 11056
rect 16347 11025 16359 11028
rect 16301 11019 16359 11025
rect 16758 11016 16764 11028
rect 16816 11056 16822 11068
rect 17126 11056 17132 11068
rect 16816 11028 17132 11056
rect 16816 11016 16822 11028
rect 17126 11016 17132 11028
rect 17184 11016 17190 11068
rect 17310 11056 17316 11068
rect 17271 11028 17316 11056
rect 17310 11016 17316 11028
rect 17368 11016 17374 11068
rect 17862 11016 17868 11068
rect 17920 11056 17926 11068
rect 19153 11059 19211 11065
rect 19153 11056 19165 11059
rect 17920 11028 19165 11056
rect 17920 11016 17926 11028
rect 19153 11025 19165 11028
rect 19199 11025 19211 11059
rect 19978 11056 19984 11068
rect 19939 11028 19984 11056
rect 19153 11019 19211 11025
rect 19978 11016 19984 11028
rect 20036 11016 20042 11068
rect 20548 11065 20576 11096
rect 20533 11059 20591 11065
rect 20533 11025 20545 11059
rect 20579 11025 20591 11059
rect 20533 11019 20591 11025
rect 8570 10948 8576 11000
rect 8628 10988 8634 11000
rect 8849 10991 8907 10997
rect 8849 10988 8861 10991
rect 8628 10960 8861 10988
rect 8628 10948 8634 10960
rect 8849 10957 8861 10960
rect 8895 10957 8907 10991
rect 14182 10988 14188 11000
rect 14143 10960 14188 10988
rect 8849 10951 8907 10957
rect 14182 10948 14188 10960
rect 14240 10948 14246 11000
rect 14274 10948 14280 11000
rect 14332 10988 14338 11000
rect 14332 10960 14377 10988
rect 14332 10948 14338 10960
rect 14550 10948 14556 11000
rect 14608 10988 14614 11000
rect 16393 10991 16451 10997
rect 16393 10988 16405 10991
rect 14608 10960 16405 10988
rect 14608 10948 14614 10960
rect 16393 10957 16405 10960
rect 16439 10957 16451 10991
rect 16393 10951 16451 10957
rect 16577 10991 16635 10997
rect 16577 10957 16589 10991
rect 16623 10957 16635 10991
rect 17494 10988 17500 11000
rect 17455 10960 17500 10988
rect 16577 10951 16635 10957
rect 12066 10880 12072 10932
rect 12124 10920 12130 10932
rect 15749 10923 15807 10929
rect 15749 10920 15761 10923
rect 12124 10892 15761 10920
rect 12124 10880 12130 10892
rect 15749 10889 15761 10892
rect 15795 10889 15807 10923
rect 15749 10883 15807 10889
rect 16482 10880 16488 10932
rect 16540 10920 16546 10932
rect 16592 10920 16620 10951
rect 17494 10948 17500 10960
rect 17552 10948 17558 11000
rect 19245 10991 19303 10997
rect 19245 10957 19257 10991
rect 19291 10957 19303 10991
rect 19245 10951 19303 10957
rect 19337 10991 19395 10997
rect 19337 10957 19349 10991
rect 19383 10957 19395 10991
rect 19337 10951 19395 10957
rect 16942 10920 16948 10932
rect 16540 10892 16620 10920
rect 16903 10892 16948 10920
rect 16540 10880 16546 10892
rect 16942 10880 16948 10892
rect 17000 10880 17006 10932
rect 19150 10880 19156 10932
rect 19208 10920 19214 10932
rect 19260 10920 19288 10951
rect 19208 10892 19288 10920
rect 19208 10880 19214 10892
rect 13446 10812 13452 10864
rect 13504 10852 13510 10864
rect 18506 10852 18512 10864
rect 13504 10824 18512 10852
rect 13504 10812 13510 10824
rect 18506 10812 18512 10824
rect 18564 10812 18570 10864
rect 19242 10812 19248 10864
rect 19300 10852 19306 10864
rect 19352 10852 19380 10951
rect 19300 10824 19380 10852
rect 19300 10812 19306 10824
rect 1104 10762 21620 10784
rect 1104 10710 4414 10762
rect 4466 10710 4478 10762
rect 4530 10710 4542 10762
rect 4594 10710 4606 10762
rect 4658 10710 11278 10762
rect 11330 10710 11342 10762
rect 11394 10710 11406 10762
rect 11458 10710 11470 10762
rect 11522 10710 18142 10762
rect 18194 10710 18206 10762
rect 18258 10710 18270 10762
rect 18322 10710 18334 10762
rect 18386 10710 21620 10762
rect 1104 10688 21620 10710
rect 1670 10608 1676 10660
rect 1728 10648 1734 10660
rect 1728 10620 11560 10648
rect 1728 10608 1734 10620
rect 8570 10580 8576 10592
rect 8531 10552 8576 10580
rect 8570 10540 8576 10552
rect 8628 10540 8634 10592
rect 11532 10521 11560 10620
rect 11698 10608 11704 10660
rect 11756 10648 11762 10660
rect 14090 10648 14096 10660
rect 11756 10620 13952 10648
rect 14051 10620 14096 10648
rect 11756 10608 11762 10620
rect 11517 10515 11575 10521
rect 11517 10481 11529 10515
rect 11563 10481 11575 10515
rect 11517 10475 11575 10481
rect 11701 10515 11759 10521
rect 11701 10481 11713 10515
rect 11747 10512 11759 10515
rect 11790 10512 11796 10524
rect 11747 10484 11796 10512
rect 11747 10481 11759 10484
rect 11701 10475 11759 10481
rect 11790 10472 11796 10484
rect 11848 10472 11854 10524
rect 12434 10472 12440 10524
rect 12492 10512 12498 10524
rect 12710 10512 12716 10524
rect 12492 10484 12716 10512
rect 12492 10472 12498 10484
rect 12710 10472 12716 10484
rect 12768 10472 12774 10524
rect 13924 10512 13952 10620
rect 14090 10608 14096 10620
rect 14148 10608 14154 10660
rect 16577 10651 16635 10657
rect 16577 10617 16589 10651
rect 16623 10648 16635 10651
rect 17310 10648 17316 10660
rect 16623 10620 17316 10648
rect 16623 10617 16635 10620
rect 16577 10611 16635 10617
rect 17310 10608 17316 10620
rect 17368 10608 17374 10660
rect 18417 10651 18475 10657
rect 18417 10617 18429 10651
rect 18463 10648 18475 10651
rect 18690 10648 18696 10660
rect 18463 10620 18696 10648
rect 18463 10617 18475 10620
rect 18417 10611 18475 10617
rect 18690 10608 18696 10620
rect 18748 10608 18754 10660
rect 19334 10608 19340 10660
rect 19392 10648 19398 10660
rect 20441 10651 20499 10657
rect 20441 10648 20453 10651
rect 19392 10620 20453 10648
rect 19392 10608 19398 10620
rect 20441 10617 20453 10620
rect 20487 10617 20499 10651
rect 20441 10611 20499 10617
rect 16482 10540 16488 10592
rect 16540 10580 16546 10592
rect 19242 10580 19248 10592
rect 16540 10552 19248 10580
rect 16540 10540 16546 10552
rect 17236 10521 17264 10552
rect 19242 10540 19248 10552
rect 19300 10540 19306 10592
rect 17221 10515 17279 10521
rect 13924 10484 16988 10512
rect 7190 10444 7196 10456
rect 7151 10416 7196 10444
rect 7190 10404 7196 10416
rect 7248 10404 7254 10456
rect 11425 10447 11483 10453
rect 11425 10413 11437 10447
rect 11471 10444 11483 10447
rect 12066 10444 12072 10456
rect 11471 10416 12072 10444
rect 11471 10413 11483 10416
rect 11425 10407 11483 10413
rect 12066 10404 12072 10416
rect 12124 10404 12130 10456
rect 12980 10447 13038 10453
rect 12980 10413 12992 10447
rect 13026 10444 13038 10447
rect 14274 10444 14280 10456
rect 13026 10416 14280 10444
rect 13026 10413 13038 10416
rect 12980 10407 13038 10413
rect 14274 10404 14280 10416
rect 14332 10404 14338 10456
rect 16960 10453 16988 10484
rect 17221 10481 17233 10515
rect 17267 10481 17279 10515
rect 17221 10475 17279 10481
rect 19061 10515 19119 10521
rect 19061 10481 19073 10515
rect 19107 10512 19119 10515
rect 19334 10512 19340 10524
rect 19107 10484 19340 10512
rect 19107 10481 19119 10484
rect 19061 10475 19119 10481
rect 19334 10472 19340 10484
rect 19392 10472 19398 10524
rect 16945 10447 17003 10453
rect 16945 10413 16957 10447
rect 16991 10444 17003 10447
rect 18966 10444 18972 10456
rect 16991 10416 18972 10444
rect 16991 10413 17003 10416
rect 16945 10407 17003 10413
rect 18966 10404 18972 10416
rect 19024 10404 19030 10456
rect 20254 10444 20260 10456
rect 20215 10416 20260 10444
rect 20254 10404 20260 10416
rect 20312 10404 20318 10456
rect 7460 10379 7518 10385
rect 7460 10345 7472 10379
rect 7506 10376 7518 10379
rect 9306 10376 9312 10388
rect 7506 10348 9312 10376
rect 7506 10345 7518 10348
rect 7460 10339 7518 10345
rect 9306 10336 9312 10348
rect 9364 10336 9370 10388
rect 18785 10379 18843 10385
rect 18785 10345 18797 10379
rect 18831 10376 18843 10379
rect 19702 10376 19708 10388
rect 18831 10348 19708 10376
rect 18831 10345 18843 10348
rect 18785 10339 18843 10345
rect 19702 10336 19708 10348
rect 19760 10336 19766 10388
rect 11054 10308 11060 10320
rect 11015 10280 11060 10308
rect 11054 10268 11060 10280
rect 11112 10268 11118 10320
rect 17034 10268 17040 10320
rect 17092 10308 17098 10320
rect 17092 10280 17137 10308
rect 17092 10268 17098 10280
rect 18874 10268 18880 10320
rect 18932 10308 18938 10320
rect 18932 10280 18977 10308
rect 18932 10268 18938 10280
rect 1104 10218 21620 10240
rect 1104 10166 7846 10218
rect 7898 10166 7910 10218
rect 7962 10166 7974 10218
rect 8026 10166 8038 10218
rect 8090 10166 14710 10218
rect 14762 10166 14774 10218
rect 14826 10166 14838 10218
rect 14890 10166 14902 10218
rect 14954 10166 21620 10218
rect 1104 10144 21620 10166
rect 10042 10104 10048 10116
rect 10003 10076 10048 10104
rect 10042 10064 10048 10076
rect 10100 10064 10106 10116
rect 10413 10107 10471 10113
rect 10413 10073 10425 10107
rect 10459 10104 10471 10107
rect 11057 10107 11115 10113
rect 11057 10104 11069 10107
rect 10459 10076 11069 10104
rect 10459 10073 10471 10076
rect 10413 10067 10471 10073
rect 11057 10073 11069 10076
rect 11103 10073 11115 10107
rect 11057 10067 11115 10073
rect 17313 10107 17371 10113
rect 17313 10073 17325 10107
rect 17359 10104 17371 10107
rect 17494 10104 17500 10116
rect 17359 10076 17500 10104
rect 17359 10073 17371 10076
rect 17313 10067 17371 10073
rect 17494 10064 17500 10076
rect 17552 10064 17558 10116
rect 19242 10064 19248 10116
rect 19300 10104 19306 10116
rect 19889 10107 19947 10113
rect 19889 10104 19901 10107
rect 19300 10076 19901 10104
rect 19300 10064 19306 10076
rect 19889 10073 19901 10076
rect 19935 10073 19947 10107
rect 19889 10067 19947 10073
rect 20717 10107 20775 10113
rect 20717 10073 20729 10107
rect 20763 10104 20775 10107
rect 21174 10104 21180 10116
rect 20763 10076 21180 10104
rect 20763 10073 20775 10076
rect 20717 10067 20775 10073
rect 21174 10064 21180 10076
rect 21232 10064 21238 10116
rect 11425 10039 11483 10045
rect 11425 10005 11437 10039
rect 11471 10036 11483 10039
rect 11606 10036 11612 10048
rect 11471 10008 11612 10036
rect 11471 10005 11483 10008
rect 11425 9999 11483 10005
rect 11606 9996 11612 10008
rect 11664 9996 11670 10048
rect 16200 10039 16258 10045
rect 16200 10005 16212 10039
rect 16246 10036 16258 10039
rect 16482 10036 16488 10048
rect 16246 10008 16488 10036
rect 16246 10005 16258 10008
rect 16200 9999 16258 10005
rect 16482 9996 16488 10008
rect 16540 9996 16546 10048
rect 11517 9971 11575 9977
rect 11517 9937 11529 9971
rect 11563 9968 11575 9971
rect 12342 9968 12348 9980
rect 11563 9940 12348 9968
rect 11563 9937 11575 9940
rect 11517 9931 11575 9937
rect 12342 9928 12348 9940
rect 12400 9928 12406 9980
rect 15194 9928 15200 9980
rect 15252 9968 15258 9980
rect 15930 9968 15936 9980
rect 15252 9940 15936 9968
rect 15252 9928 15258 9940
rect 15930 9928 15936 9940
rect 15988 9928 15994 9980
rect 18776 9971 18834 9977
rect 18776 9937 18788 9971
rect 18822 9968 18834 9971
rect 19334 9968 19340 9980
rect 18822 9940 19340 9968
rect 18822 9937 18834 9940
rect 18776 9931 18834 9937
rect 19334 9928 19340 9940
rect 19392 9928 19398 9980
rect 20530 9968 20536 9980
rect 20491 9940 20536 9968
rect 20530 9928 20536 9940
rect 20588 9928 20594 9980
rect 10502 9900 10508 9912
rect 10463 9872 10508 9900
rect 10502 9860 10508 9872
rect 10560 9860 10566 9912
rect 10597 9903 10655 9909
rect 10597 9869 10609 9903
rect 10643 9869 10655 9903
rect 10597 9863 10655 9869
rect 9306 9792 9312 9844
rect 9364 9832 9370 9844
rect 10612 9832 10640 9863
rect 11146 9860 11152 9912
rect 11204 9900 11210 9912
rect 11609 9903 11667 9909
rect 11609 9900 11621 9903
rect 11204 9872 11621 9900
rect 11204 9860 11210 9872
rect 11609 9869 11621 9872
rect 11655 9869 11667 9903
rect 11609 9863 11667 9869
rect 17954 9860 17960 9912
rect 18012 9900 18018 9912
rect 18509 9903 18567 9909
rect 18509 9900 18521 9903
rect 18012 9872 18521 9900
rect 18012 9860 18018 9872
rect 18509 9869 18521 9872
rect 18555 9869 18567 9903
rect 18509 9863 18567 9869
rect 9364 9804 10640 9832
rect 9364 9792 9370 9804
rect 1104 9674 21620 9696
rect 1104 9622 4414 9674
rect 4466 9622 4478 9674
rect 4530 9622 4542 9674
rect 4594 9622 4606 9674
rect 4658 9622 11278 9674
rect 11330 9622 11342 9674
rect 11394 9622 11406 9674
rect 11458 9622 11470 9674
rect 11522 9622 18142 9674
rect 18194 9622 18206 9674
rect 18258 9622 18270 9674
rect 18322 9622 18334 9674
rect 18386 9622 21620 9674
rect 1104 9600 21620 9622
rect 10502 9560 10508 9572
rect 10463 9532 10508 9560
rect 10502 9520 10508 9532
rect 10560 9520 10566 9572
rect 12342 9560 12348 9572
rect 12303 9532 12348 9560
rect 12342 9520 12348 9532
rect 12400 9520 12406 9572
rect 17034 9560 17040 9572
rect 12452 9532 17040 9560
rect 9306 9492 9312 9504
rect 9267 9464 9312 9492
rect 9306 9452 9312 9464
rect 9364 9452 9370 9504
rect 12158 9452 12164 9504
rect 12216 9492 12222 9504
rect 12452 9492 12480 9532
rect 17034 9520 17040 9532
rect 17092 9520 17098 9572
rect 18693 9563 18751 9569
rect 18693 9529 18705 9563
rect 18739 9560 18751 9563
rect 18874 9560 18880 9572
rect 18739 9532 18880 9560
rect 18739 9529 18751 9532
rect 18693 9523 18751 9529
rect 18874 9520 18880 9532
rect 18932 9520 18938 9572
rect 12216 9464 12480 9492
rect 12216 9452 12222 9464
rect 12710 9452 12716 9504
rect 12768 9492 12774 9504
rect 14921 9495 14979 9501
rect 12768 9464 13584 9492
rect 12768 9452 12774 9464
rect 11146 9424 11152 9436
rect 11107 9396 11152 9424
rect 11146 9384 11152 9396
rect 11204 9384 11210 9436
rect 11517 9427 11575 9433
rect 11517 9393 11529 9427
rect 11563 9424 11575 9427
rect 11606 9424 11612 9436
rect 11563 9396 11612 9424
rect 11563 9393 11575 9396
rect 11517 9387 11575 9393
rect 11606 9384 11612 9396
rect 11664 9384 11670 9436
rect 11790 9384 11796 9436
rect 11848 9424 11854 9436
rect 13556 9433 13584 9464
rect 14921 9461 14933 9495
rect 14967 9461 14979 9495
rect 14921 9455 14979 9461
rect 12989 9427 13047 9433
rect 12989 9424 13001 9427
rect 11848 9396 13001 9424
rect 11848 9384 11854 9396
rect 12989 9393 13001 9396
rect 13035 9393 13047 9427
rect 12989 9387 13047 9393
rect 13541 9427 13599 9433
rect 13541 9393 13553 9427
rect 13587 9393 13599 9427
rect 13541 9387 13599 9393
rect 7190 9316 7196 9368
rect 7248 9356 7254 9368
rect 7929 9359 7987 9365
rect 7929 9356 7941 9359
rect 7248 9328 7941 9356
rect 7248 9316 7254 9328
rect 7929 9325 7941 9328
rect 7975 9325 7987 9359
rect 7929 9319 7987 9325
rect 8196 9359 8254 9365
rect 8196 9325 8208 9359
rect 8242 9356 8254 9359
rect 11164 9356 11192 9384
rect 8242 9328 11192 9356
rect 8242 9325 8254 9328
rect 8196 9319 8254 9325
rect 7944 9220 7972 9319
rect 10965 9291 11023 9297
rect 10965 9257 10977 9291
rect 11011 9288 11023 9291
rect 11054 9288 11060 9300
rect 11011 9260 11060 9288
rect 11011 9257 11023 9260
rect 10965 9251 11023 9257
rect 11054 9248 11060 9260
rect 11112 9248 11118 9300
rect 12713 9291 12771 9297
rect 12713 9257 12725 9291
rect 12759 9288 12771 9291
rect 12894 9288 12900 9300
rect 12759 9260 12900 9288
rect 12759 9257 12771 9260
rect 12713 9251 12771 9257
rect 12894 9248 12900 9260
rect 12952 9248 12958 9300
rect 13004 9288 13032 9387
rect 13808 9359 13866 9365
rect 13808 9325 13820 9359
rect 13854 9356 13866 9359
rect 14090 9356 14096 9368
rect 13854 9328 14096 9356
rect 13854 9325 13866 9328
rect 13808 9319 13866 9325
rect 14090 9316 14096 9328
rect 14148 9316 14154 9368
rect 14936 9288 14964 9455
rect 15010 9452 15016 9504
rect 15068 9492 15074 9504
rect 15473 9495 15531 9501
rect 15473 9492 15485 9495
rect 15068 9464 15485 9492
rect 15068 9452 15074 9464
rect 15473 9461 15485 9464
rect 15519 9461 15531 9495
rect 15473 9455 15531 9461
rect 19245 9427 19303 9433
rect 19245 9393 19257 9427
rect 19291 9424 19303 9427
rect 19426 9424 19432 9436
rect 19291 9396 19432 9424
rect 19291 9393 19303 9396
rect 19245 9387 19303 9393
rect 19426 9384 19432 9396
rect 19484 9384 19490 9436
rect 19702 9424 19708 9436
rect 19663 9396 19708 9424
rect 19702 9384 19708 9396
rect 19760 9384 19766 9436
rect 15286 9356 15292 9368
rect 15247 9328 15292 9356
rect 15286 9316 15292 9328
rect 15344 9316 15350 9368
rect 19058 9356 19064 9368
rect 19019 9328 19064 9356
rect 19058 9316 19064 9328
rect 19116 9316 19122 9368
rect 13004 9260 14964 9288
rect 8202 9220 8208 9232
rect 7944 9192 8208 9220
rect 8202 9180 8208 9192
rect 8260 9180 8266 9232
rect 10870 9220 10876 9232
rect 10831 9192 10876 9220
rect 10870 9180 10876 9192
rect 10928 9180 10934 9232
rect 12805 9223 12863 9229
rect 12805 9189 12817 9223
rect 12851 9220 12863 9223
rect 15746 9220 15752 9232
rect 12851 9192 15752 9220
rect 12851 9189 12863 9192
rect 12805 9183 12863 9189
rect 15746 9180 15752 9192
rect 15804 9180 15810 9232
rect 19150 9220 19156 9232
rect 19111 9192 19156 9220
rect 19150 9180 19156 9192
rect 19208 9180 19214 9232
rect 1104 9130 21620 9152
rect 1104 9078 7846 9130
rect 7898 9078 7910 9130
rect 7962 9078 7974 9130
rect 8026 9078 8038 9130
rect 8090 9078 14710 9130
rect 14762 9078 14774 9130
rect 14826 9078 14838 9130
rect 14890 9078 14902 9130
rect 14954 9078 21620 9130
rect 1104 9056 21620 9078
rect 10870 8976 10876 9028
rect 10928 9016 10934 9028
rect 10965 9019 11023 9025
rect 10965 9016 10977 9019
rect 10928 8988 10977 9016
rect 10928 8976 10934 8988
rect 10965 8985 10977 8988
rect 11011 8985 11023 9019
rect 10965 8979 11023 8985
rect 11425 9019 11483 9025
rect 11425 8985 11437 9019
rect 11471 9016 11483 9019
rect 12158 9016 12164 9028
rect 11471 8988 12164 9016
rect 11471 8985 11483 8988
rect 11425 8979 11483 8985
rect 12158 8976 12164 8988
rect 12216 8976 12222 9028
rect 13262 8976 13268 9028
rect 13320 9016 13326 9028
rect 13449 9019 13507 9025
rect 13449 9016 13461 9019
rect 13320 8988 13461 9016
rect 13320 8976 13326 8988
rect 13449 8985 13461 8988
rect 13495 8985 13507 9019
rect 17862 9016 17868 9028
rect 13449 8979 13507 8985
rect 13556 8988 17868 9016
rect 11333 8951 11391 8957
rect 11333 8917 11345 8951
rect 11379 8948 11391 8951
rect 11698 8948 11704 8960
rect 11379 8920 11704 8948
rect 11379 8917 11391 8920
rect 11333 8911 11391 8917
rect 11698 8908 11704 8920
rect 11756 8908 11762 8960
rect 12894 8908 12900 8960
rect 12952 8948 12958 8960
rect 13556 8948 13584 8988
rect 17862 8976 17868 8988
rect 17920 8976 17926 9028
rect 19334 8976 19340 9028
rect 19392 9016 19398 9028
rect 19705 9019 19763 9025
rect 19705 9016 19717 9019
rect 19392 8988 19717 9016
rect 19392 8976 19398 8988
rect 19705 8985 19717 8988
rect 19751 8985 19763 9019
rect 19705 8979 19763 8985
rect 20165 9019 20223 9025
rect 20165 8985 20177 9019
rect 20211 9016 20223 9019
rect 20346 9016 20352 9028
rect 20211 8988 20352 9016
rect 20211 8985 20223 8988
rect 20165 8979 20223 8985
rect 20346 8976 20352 8988
rect 20404 8976 20410 9028
rect 20717 9019 20775 9025
rect 20717 8985 20729 9019
rect 20763 9016 20775 9019
rect 21450 9016 21456 9028
rect 20763 8988 21456 9016
rect 20763 8985 20775 8988
rect 20717 8979 20775 8985
rect 21450 8976 21456 8988
rect 21508 8976 21514 9028
rect 12952 8920 13584 8948
rect 12952 8908 12958 8920
rect 15286 8908 15292 8960
rect 15344 8948 15350 8960
rect 15749 8951 15807 8957
rect 15749 8948 15761 8951
rect 15344 8920 15761 8948
rect 15344 8908 15350 8920
rect 15749 8917 15761 8920
rect 15795 8917 15807 8951
rect 15749 8911 15807 8917
rect 8472 8883 8530 8889
rect 8472 8849 8484 8883
rect 8518 8880 8530 8883
rect 11790 8880 11796 8892
rect 8518 8852 11796 8880
rect 8518 8849 8530 8852
rect 8472 8843 8530 8849
rect 8202 8812 8208 8824
rect 8163 8784 8208 8812
rect 8202 8772 8208 8784
rect 8260 8772 8266 8824
rect 11532 8821 11560 8852
rect 11790 8840 11796 8852
rect 11848 8840 11854 8892
rect 13265 8883 13323 8889
rect 13265 8849 13277 8883
rect 13311 8880 13323 8883
rect 13538 8880 13544 8892
rect 13311 8852 13544 8880
rect 13311 8849 13323 8852
rect 13265 8843 13323 8849
rect 13538 8840 13544 8852
rect 13596 8840 13602 8892
rect 15473 8883 15531 8889
rect 15473 8849 15485 8883
rect 15519 8880 15531 8883
rect 16298 8880 16304 8892
rect 15519 8852 16304 8880
rect 15519 8849 15531 8852
rect 15473 8843 15531 8849
rect 16298 8840 16304 8852
rect 16356 8840 16362 8892
rect 18592 8883 18650 8889
rect 18592 8849 18604 8883
rect 18638 8880 18650 8883
rect 19426 8880 19432 8892
rect 18638 8852 19432 8880
rect 18638 8849 18650 8852
rect 18592 8843 18650 8849
rect 19426 8840 19432 8852
rect 19484 8840 19490 8892
rect 19978 8880 19984 8892
rect 19939 8852 19984 8880
rect 19978 8840 19984 8852
rect 20036 8840 20042 8892
rect 20530 8880 20536 8892
rect 20491 8852 20536 8880
rect 20530 8840 20536 8852
rect 20588 8840 20594 8892
rect 11517 8815 11575 8821
rect 11517 8781 11529 8815
rect 11563 8781 11575 8815
rect 11517 8775 11575 8781
rect 17954 8772 17960 8824
rect 18012 8812 18018 8824
rect 18325 8815 18383 8821
rect 18325 8812 18337 8815
rect 18012 8784 18337 8812
rect 18012 8772 18018 8784
rect 18325 8781 18337 8784
rect 18371 8781 18383 8815
rect 18325 8775 18383 8781
rect 9585 8747 9643 8753
rect 9585 8713 9597 8747
rect 9631 8744 9643 8747
rect 11146 8744 11152 8756
rect 9631 8716 11152 8744
rect 9631 8713 9643 8716
rect 9585 8707 9643 8713
rect 11146 8704 11152 8716
rect 11204 8704 11210 8756
rect 1104 8586 21620 8608
rect 1104 8534 4414 8586
rect 4466 8534 4478 8586
rect 4530 8534 4542 8586
rect 4594 8534 4606 8586
rect 4658 8534 11278 8586
rect 11330 8534 11342 8586
rect 11394 8534 11406 8586
rect 11458 8534 11470 8586
rect 11522 8534 18142 8586
rect 18194 8534 18206 8586
rect 18258 8534 18270 8586
rect 18322 8534 18334 8586
rect 18386 8534 21620 8586
rect 1104 8512 21620 8534
rect 11517 8475 11575 8481
rect 11517 8441 11529 8475
rect 11563 8472 11575 8475
rect 11882 8472 11888 8484
rect 11563 8444 11888 8472
rect 11563 8441 11575 8444
rect 11517 8435 11575 8441
rect 11882 8432 11888 8444
rect 11940 8432 11946 8484
rect 16298 8472 16304 8484
rect 16259 8444 16304 8472
rect 16298 8432 16304 8444
rect 16356 8432 16362 8484
rect 19794 8432 19800 8484
rect 19852 8472 19858 8484
rect 20441 8475 20499 8481
rect 20441 8472 20453 8475
rect 19852 8444 20453 8472
rect 19852 8432 19858 8444
rect 20441 8441 20453 8444
rect 20487 8441 20499 8475
rect 20441 8435 20499 8441
rect 13538 8336 13544 8348
rect 13499 8308 13544 8336
rect 13538 8296 13544 8308
rect 13596 8296 13602 8348
rect 16945 8339 17003 8345
rect 16945 8305 16957 8339
rect 16991 8336 17003 8339
rect 17678 8336 17684 8348
rect 16991 8308 17684 8336
rect 16991 8305 17003 8308
rect 16945 8299 17003 8305
rect 17678 8296 17684 8308
rect 17736 8296 17742 8348
rect 11330 8268 11336 8280
rect 11291 8240 11336 8268
rect 11330 8228 11336 8240
rect 11388 8228 11394 8280
rect 13354 8268 13360 8280
rect 13315 8240 13360 8268
rect 13354 8228 13360 8240
rect 13412 8228 13418 8280
rect 20254 8268 20260 8280
rect 20215 8240 20260 8268
rect 20254 8228 20260 8240
rect 20312 8228 20318 8280
rect 16669 8203 16727 8209
rect 16669 8169 16681 8203
rect 16715 8200 16727 8203
rect 17313 8203 17371 8209
rect 17313 8200 17325 8203
rect 16715 8172 17325 8200
rect 16715 8169 16727 8172
rect 16669 8163 16727 8169
rect 17313 8169 17325 8172
rect 17359 8169 17371 8203
rect 17313 8163 17371 8169
rect 10686 8132 10692 8144
rect 10647 8104 10692 8132
rect 10686 8092 10692 8104
rect 10744 8092 10750 8144
rect 16758 8132 16764 8144
rect 16719 8104 16764 8132
rect 16758 8092 16764 8104
rect 16816 8092 16822 8144
rect 1104 8042 21620 8064
rect 1104 7990 7846 8042
rect 7898 7990 7910 8042
rect 7962 7990 7974 8042
rect 8026 7990 8038 8042
rect 8090 7990 14710 8042
rect 14762 7990 14774 8042
rect 14826 7990 14838 8042
rect 14890 7990 14902 8042
rect 14954 7990 21620 8042
rect 1104 7968 21620 7990
rect 10686 7888 10692 7940
rect 10744 7928 10750 7940
rect 10781 7931 10839 7937
rect 10781 7928 10793 7931
rect 10744 7900 10793 7928
rect 10744 7888 10750 7900
rect 10781 7897 10793 7900
rect 10827 7897 10839 7931
rect 10781 7891 10839 7897
rect 13354 7888 13360 7940
rect 13412 7928 13418 7940
rect 13725 7931 13783 7937
rect 13725 7928 13737 7931
rect 13412 7900 13737 7928
rect 13412 7888 13418 7900
rect 13725 7897 13737 7900
rect 13771 7897 13783 7931
rect 16666 7928 16672 7940
rect 13725 7891 13783 7897
rect 16592 7900 16672 7928
rect 11330 7820 11336 7872
rect 11388 7860 11394 7872
rect 16592 7869 16620 7900
rect 16666 7888 16672 7900
rect 16724 7888 16730 7940
rect 17678 7928 17684 7940
rect 17639 7900 17684 7928
rect 17678 7888 17684 7900
rect 17736 7888 17742 7940
rect 19426 7928 19432 7940
rect 19387 7900 19432 7928
rect 19426 7888 19432 7900
rect 19484 7888 19490 7940
rect 11701 7863 11759 7869
rect 11701 7860 11713 7863
rect 11388 7832 11713 7860
rect 11388 7820 11394 7832
rect 11701 7829 11713 7832
rect 11747 7829 11759 7863
rect 11701 7823 11759 7829
rect 16568 7863 16626 7869
rect 16568 7829 16580 7863
rect 16614 7829 16626 7863
rect 16568 7823 16626 7829
rect 16850 7820 16856 7872
rect 16908 7860 16914 7872
rect 17696 7860 17724 7888
rect 18294 7863 18352 7869
rect 18294 7860 18306 7863
rect 16908 7832 17632 7860
rect 17696 7832 18306 7860
rect 16908 7820 16914 7832
rect 11425 7795 11483 7801
rect 11425 7792 11437 7795
rect 10428 7764 11437 7792
rect 10428 7665 10456 7764
rect 11425 7761 11437 7764
rect 11471 7761 11483 7795
rect 11425 7755 11483 7761
rect 14093 7795 14151 7801
rect 14093 7761 14105 7795
rect 14139 7792 14151 7795
rect 14642 7792 14648 7804
rect 14139 7764 14648 7792
rect 14139 7761 14151 7764
rect 14093 7755 14151 7761
rect 14642 7752 14648 7764
rect 14700 7752 14706 7804
rect 15930 7752 15936 7804
rect 15988 7792 15994 7804
rect 16301 7795 16359 7801
rect 16301 7792 16313 7795
rect 15988 7764 16313 7792
rect 15988 7752 15994 7764
rect 16301 7761 16313 7764
rect 16347 7792 16359 7795
rect 17604 7792 17632 7832
rect 18294 7829 18306 7832
rect 18340 7829 18352 7863
rect 18294 7823 18352 7829
rect 19978 7792 19984 7804
rect 16347 7764 17356 7792
rect 17604 7764 19104 7792
rect 19939 7764 19984 7792
rect 16347 7761 16359 7764
rect 16301 7755 16359 7761
rect 10870 7724 10876 7736
rect 10831 7696 10876 7724
rect 10870 7684 10876 7696
rect 10928 7684 10934 7736
rect 11054 7724 11060 7736
rect 11015 7696 11060 7724
rect 11054 7684 11060 7696
rect 11112 7684 11118 7736
rect 14182 7724 14188 7736
rect 14143 7696 14188 7724
rect 14182 7684 14188 7696
rect 14240 7684 14246 7736
rect 14366 7724 14372 7736
rect 14327 7696 14372 7724
rect 14366 7684 14372 7696
rect 14424 7684 14430 7736
rect 17328 7724 17356 7764
rect 17954 7724 17960 7736
rect 17328 7696 17960 7724
rect 17954 7684 17960 7696
rect 18012 7724 18018 7736
rect 18049 7727 18107 7733
rect 18049 7724 18061 7727
rect 18012 7696 18061 7724
rect 18012 7684 18018 7696
rect 18049 7693 18061 7696
rect 18095 7693 18107 7727
rect 18049 7687 18107 7693
rect 10413 7659 10471 7665
rect 10413 7625 10425 7659
rect 10459 7625 10471 7659
rect 19076 7656 19104 7764
rect 19978 7752 19984 7764
rect 20036 7752 20042 7804
rect 20530 7792 20536 7804
rect 20491 7764 20536 7792
rect 20530 7752 20536 7764
rect 20588 7752 20594 7804
rect 20717 7659 20775 7665
rect 20717 7656 20729 7659
rect 19076 7628 20729 7656
rect 10413 7619 10471 7625
rect 20717 7625 20729 7628
rect 20763 7625 20775 7659
rect 20717 7619 20775 7625
rect 13906 7548 13912 7600
rect 13964 7588 13970 7600
rect 20165 7591 20223 7597
rect 20165 7588 20177 7591
rect 13964 7560 20177 7588
rect 13964 7548 13970 7560
rect 20165 7557 20177 7560
rect 20211 7557 20223 7591
rect 20165 7551 20223 7557
rect 1104 7498 21620 7520
rect 1104 7446 4414 7498
rect 4466 7446 4478 7498
rect 4530 7446 4542 7498
rect 4594 7446 4606 7498
rect 4658 7446 11278 7498
rect 11330 7446 11342 7498
rect 11394 7446 11406 7498
rect 11458 7446 11470 7498
rect 11522 7446 18142 7498
rect 18194 7446 18206 7498
rect 18258 7446 18270 7498
rect 18322 7446 18334 7498
rect 18386 7446 21620 7498
rect 1104 7424 21620 7446
rect 11054 7384 11060 7396
rect 11015 7356 11060 7384
rect 11054 7344 11060 7356
rect 11112 7344 11118 7396
rect 16666 7384 16672 7396
rect 16627 7356 16672 7384
rect 16666 7344 16672 7356
rect 16724 7344 16730 7396
rect 16758 7344 16764 7396
rect 16816 7384 16822 7396
rect 16945 7387 17003 7393
rect 16945 7384 16957 7387
rect 16816 7356 16957 7384
rect 16816 7344 16822 7356
rect 16945 7353 16957 7356
rect 16991 7353 17003 7387
rect 16945 7347 17003 7353
rect 7374 7140 7380 7192
rect 7432 7180 7438 7192
rect 8202 7180 8208 7192
rect 7432 7152 8208 7180
rect 7432 7140 7438 7152
rect 8202 7140 8208 7152
rect 8260 7180 8266 7192
rect 9677 7183 9735 7189
rect 9677 7180 9689 7183
rect 8260 7152 9689 7180
rect 8260 7140 8266 7152
rect 9677 7149 9689 7152
rect 9723 7149 9735 7183
rect 9677 7143 9735 7149
rect 9858 7072 9864 7124
rect 9916 7121 9922 7124
rect 9916 7115 9980 7121
rect 9916 7081 9934 7115
rect 9968 7081 9980 7115
rect 11072 7112 11100 7344
rect 14366 7316 14372 7328
rect 14279 7288 14372 7316
rect 14366 7276 14372 7288
rect 14424 7316 14430 7328
rect 14424 7288 14780 7316
rect 14424 7276 14430 7288
rect 11241 7251 11299 7257
rect 11241 7217 11253 7251
rect 11287 7248 11299 7251
rect 11333 7251 11391 7257
rect 11333 7248 11345 7251
rect 11287 7220 11345 7248
rect 11287 7217 11299 7220
rect 11241 7211 11299 7217
rect 11333 7217 11345 7220
rect 11379 7217 11391 7251
rect 14642 7248 14648 7260
rect 14603 7220 14648 7248
rect 11333 7211 11391 7217
rect 14642 7208 14648 7220
rect 14700 7208 14706 7260
rect 12710 7140 12716 7192
rect 12768 7180 12774 7192
rect 12989 7183 13047 7189
rect 12989 7180 13001 7183
rect 12768 7152 13001 7180
rect 12768 7140 12774 7152
rect 12989 7149 13001 7152
rect 13035 7149 13047 7183
rect 13256 7183 13314 7189
rect 13256 7180 13268 7183
rect 12989 7143 13047 7149
rect 13188 7152 13268 7180
rect 11578 7115 11636 7121
rect 11578 7112 11590 7115
rect 11072 7084 11590 7112
rect 9916 7075 9980 7081
rect 11578 7081 11590 7084
rect 11624 7081 11636 7115
rect 12728 7112 12756 7140
rect 11578 7075 11636 7081
rect 12360 7084 12756 7112
rect 9916 7072 9922 7075
rect 11241 7047 11299 7053
rect 11241 7013 11253 7047
rect 11287 7044 11299 7047
rect 12360 7044 12388 7084
rect 11287 7016 12388 7044
rect 12713 7047 12771 7053
rect 11287 7013 11299 7016
rect 11241 7007 11299 7013
rect 12713 7013 12725 7047
rect 12759 7044 12771 7047
rect 13188 7044 13216 7152
rect 13256 7149 13268 7152
rect 13302 7180 13314 7183
rect 14550 7180 14556 7192
rect 13302 7152 14556 7180
rect 13302 7149 13314 7152
rect 13256 7143 13314 7149
rect 14550 7140 14556 7152
rect 14608 7140 14614 7192
rect 14752 7112 14780 7288
rect 16684 7248 16712 7344
rect 17497 7251 17555 7257
rect 17497 7248 17509 7251
rect 16684 7220 17509 7248
rect 17497 7217 17509 7220
rect 17543 7217 17555 7251
rect 17497 7211 17555 7217
rect 15289 7183 15347 7189
rect 15289 7149 15301 7183
rect 15335 7180 15347 7183
rect 15930 7180 15936 7192
rect 15335 7152 15936 7180
rect 15335 7149 15347 7152
rect 15289 7143 15347 7149
rect 15930 7140 15936 7152
rect 15988 7140 15994 7192
rect 17402 7180 17408 7192
rect 17315 7152 17408 7180
rect 17402 7140 17408 7152
rect 17460 7180 17466 7192
rect 19150 7180 19156 7192
rect 17460 7152 19156 7180
rect 17460 7140 17466 7152
rect 19150 7140 19156 7152
rect 19208 7140 19214 7192
rect 15534 7115 15592 7121
rect 15534 7112 15546 7115
rect 14752 7084 15546 7112
rect 15534 7081 15546 7084
rect 15580 7081 15592 7115
rect 15534 7075 15592 7081
rect 17313 7115 17371 7121
rect 17313 7081 17325 7115
rect 17359 7112 17371 7115
rect 18506 7112 18512 7124
rect 17359 7084 18512 7112
rect 17359 7081 17371 7084
rect 17313 7075 17371 7081
rect 18506 7072 18512 7084
rect 18564 7072 18570 7124
rect 12759 7016 13216 7044
rect 12759 7013 12771 7016
rect 12713 7007 12771 7013
rect 1104 6954 21620 6976
rect 1104 6902 7846 6954
rect 7898 6902 7910 6954
rect 7962 6902 7974 6954
rect 8026 6902 8038 6954
rect 8090 6902 14710 6954
rect 14762 6902 14774 6954
rect 14826 6902 14838 6954
rect 14890 6902 14902 6954
rect 14954 6902 21620 6954
rect 1104 6880 21620 6902
rect 10597 6843 10655 6849
rect 10597 6809 10609 6843
rect 10643 6840 10655 6843
rect 10870 6840 10876 6852
rect 10643 6812 10876 6840
rect 10643 6809 10655 6812
rect 10597 6803 10655 6809
rect 10870 6800 10876 6812
rect 10928 6800 10934 6852
rect 14093 6843 14151 6849
rect 14093 6809 14105 6843
rect 14139 6840 14151 6843
rect 14182 6840 14188 6852
rect 14139 6812 14188 6840
rect 14139 6809 14151 6812
rect 14093 6803 14151 6809
rect 14182 6800 14188 6812
rect 14240 6800 14246 6852
rect 16482 6840 16488 6852
rect 14384 6812 16488 6840
rect 10965 6775 11023 6781
rect 10965 6741 10977 6775
rect 11011 6772 11023 6775
rect 14384 6772 14412 6812
rect 16482 6800 16488 6812
rect 16540 6800 16546 6852
rect 11011 6744 14412 6772
rect 14461 6775 14519 6781
rect 11011 6741 11023 6744
rect 10965 6735 11023 6741
rect 14461 6741 14473 6775
rect 14507 6772 14519 6775
rect 14507 6744 16528 6772
rect 14507 6741 14519 6744
rect 14461 6735 14519 6741
rect 4062 6664 4068 6716
rect 4120 6704 4126 6716
rect 7633 6707 7691 6713
rect 7633 6704 7645 6707
rect 4120 6676 7645 6704
rect 4120 6664 4126 6676
rect 7633 6673 7645 6676
rect 7679 6673 7691 6707
rect 7633 6667 7691 6673
rect 10594 6664 10600 6716
rect 10652 6704 10658 6716
rect 11057 6707 11115 6713
rect 11057 6704 11069 6707
rect 10652 6676 11069 6704
rect 10652 6664 10658 6676
rect 11057 6673 11069 6676
rect 11103 6704 11115 6707
rect 14553 6707 14611 6713
rect 14553 6704 14565 6707
rect 11103 6676 14565 6704
rect 11103 6673 11115 6676
rect 11057 6667 11115 6673
rect 14553 6673 14565 6676
rect 14599 6704 14611 6707
rect 16500 6704 16528 6744
rect 18598 6704 18604 6716
rect 14599 6676 15884 6704
rect 16500 6676 18604 6704
rect 14599 6673 14611 6676
rect 14553 6667 14611 6673
rect 7374 6636 7380 6648
rect 7335 6608 7380 6636
rect 7374 6596 7380 6608
rect 7432 6596 7438 6648
rect 11149 6639 11207 6645
rect 11149 6605 11161 6639
rect 11195 6605 11207 6639
rect 11149 6599 11207 6605
rect 8757 6571 8815 6577
rect 8757 6537 8769 6571
rect 8803 6568 8815 6571
rect 9858 6568 9864 6580
rect 8803 6540 9864 6568
rect 8803 6537 8815 6540
rect 8757 6531 8815 6537
rect 9858 6528 9864 6540
rect 9916 6568 9922 6580
rect 11164 6568 11192 6599
rect 14642 6596 14648 6648
rect 14700 6636 14706 6648
rect 15856 6636 15884 6676
rect 18598 6664 18604 6676
rect 18656 6664 18662 6716
rect 20530 6704 20536 6716
rect 20491 6676 20536 6704
rect 20530 6664 20536 6676
rect 20588 6664 20594 6716
rect 17402 6636 17408 6648
rect 14700 6608 14745 6636
rect 15856 6608 17408 6636
rect 14700 6596 14706 6608
rect 17402 6596 17408 6608
rect 17460 6596 17466 6648
rect 9916 6540 11192 6568
rect 9916 6528 9922 6540
rect 13630 6528 13636 6580
rect 13688 6568 13694 6580
rect 20717 6571 20775 6577
rect 20717 6568 20729 6571
rect 13688 6540 20729 6568
rect 13688 6528 13694 6540
rect 20717 6537 20729 6540
rect 20763 6537 20775 6571
rect 20717 6531 20775 6537
rect 1104 6410 21620 6432
rect 1104 6358 4414 6410
rect 4466 6358 4478 6410
rect 4530 6358 4542 6410
rect 4594 6358 4606 6410
rect 4658 6358 11278 6410
rect 11330 6358 11342 6410
rect 11394 6358 11406 6410
rect 11458 6358 11470 6410
rect 11522 6358 18142 6410
rect 18194 6358 18206 6410
rect 18258 6358 18270 6410
rect 18322 6358 18334 6410
rect 18386 6358 21620 6410
rect 1104 6336 21620 6358
rect 1104 5866 21620 5888
rect 1104 5814 7846 5866
rect 7898 5814 7910 5866
rect 7962 5814 7974 5866
rect 8026 5814 8038 5866
rect 8090 5814 14710 5866
rect 14762 5814 14774 5866
rect 14826 5814 14838 5866
rect 14890 5814 14902 5866
rect 14954 5814 21620 5866
rect 1104 5792 21620 5814
rect 12986 5712 12992 5764
rect 13044 5752 13050 5764
rect 20717 5755 20775 5761
rect 20717 5752 20729 5755
rect 13044 5724 20729 5752
rect 13044 5712 13050 5724
rect 20717 5721 20729 5724
rect 20763 5721 20775 5755
rect 20717 5715 20775 5721
rect 20530 5616 20536 5628
rect 20491 5588 20536 5616
rect 20530 5576 20536 5588
rect 20588 5576 20594 5628
rect 1104 5322 21620 5344
rect 1104 5270 4414 5322
rect 4466 5270 4478 5322
rect 4530 5270 4542 5322
rect 4594 5270 4606 5322
rect 4658 5270 11278 5322
rect 11330 5270 11342 5322
rect 11394 5270 11406 5322
rect 11458 5270 11470 5322
rect 11522 5270 18142 5322
rect 18194 5270 18206 5322
rect 18258 5270 18270 5322
rect 18322 5270 18334 5322
rect 18386 5270 21620 5322
rect 1104 5248 21620 5270
rect 16482 5168 16488 5220
rect 16540 5208 16546 5220
rect 17954 5208 17960 5220
rect 16540 5180 17960 5208
rect 16540 5168 16546 5180
rect 17954 5168 17960 5180
rect 18012 5168 18018 5220
rect 1104 4778 21620 4800
rect 1104 4726 7846 4778
rect 7898 4726 7910 4778
rect 7962 4726 7974 4778
rect 8026 4726 8038 4778
rect 8090 4726 14710 4778
rect 14762 4726 14774 4778
rect 14826 4726 14838 4778
rect 14890 4726 14902 4778
rect 14954 4726 21620 4778
rect 1104 4704 21620 4726
rect 20717 4667 20775 4673
rect 20717 4633 20729 4667
rect 20763 4664 20775 4667
rect 21082 4664 21088 4676
rect 20763 4636 21088 4664
rect 20763 4633 20775 4636
rect 20717 4627 20775 4633
rect 21082 4624 21088 4636
rect 21140 4624 21146 4676
rect 20530 4528 20536 4540
rect 20491 4500 20536 4528
rect 20530 4488 20536 4500
rect 20588 4488 20594 4540
rect 1104 4234 21620 4256
rect 1104 4182 4414 4234
rect 4466 4182 4478 4234
rect 4530 4182 4542 4234
rect 4594 4182 4606 4234
rect 4658 4182 11278 4234
rect 11330 4182 11342 4234
rect 11394 4182 11406 4234
rect 11458 4182 11470 4234
rect 11522 4182 18142 4234
rect 18194 4182 18206 4234
rect 18258 4182 18270 4234
rect 18322 4182 18334 4234
rect 18386 4182 21620 4234
rect 1104 4160 21620 4182
rect 14274 3944 14280 3996
rect 14332 3984 14338 3996
rect 18506 3984 18512 3996
rect 14332 3956 18512 3984
rect 14332 3944 14338 3956
rect 18506 3944 18512 3956
rect 18564 3944 18570 3996
rect 1104 3690 21620 3712
rect 1104 3638 7846 3690
rect 7898 3638 7910 3690
rect 7962 3638 7974 3690
rect 8026 3638 8038 3690
rect 8090 3638 14710 3690
rect 14762 3638 14774 3690
rect 14826 3638 14838 3690
rect 14890 3638 14902 3690
rect 14954 3638 21620 3690
rect 1104 3616 21620 3638
rect 1104 3146 21620 3168
rect 1104 3094 4414 3146
rect 4466 3094 4478 3146
rect 4530 3094 4542 3146
rect 4594 3094 4606 3146
rect 4658 3094 11278 3146
rect 11330 3094 11342 3146
rect 11394 3094 11406 3146
rect 11458 3094 11470 3146
rect 11522 3094 18142 3146
rect 18194 3094 18206 3146
rect 18258 3094 18270 3146
rect 18322 3094 18334 3146
rect 18386 3094 21620 3146
rect 1104 3072 21620 3094
rect 1104 2602 21620 2624
rect 1104 2550 7846 2602
rect 7898 2550 7910 2602
rect 7962 2550 7974 2602
rect 8026 2550 8038 2602
rect 8090 2550 14710 2602
rect 14762 2550 14774 2602
rect 14826 2550 14838 2602
rect 14890 2550 14902 2602
rect 14954 2550 21620 2602
rect 1104 2528 21620 2550
rect 14458 2448 14464 2500
rect 14516 2488 14522 2500
rect 18598 2488 18604 2500
rect 14516 2460 18604 2488
rect 14516 2448 14522 2460
rect 18598 2448 18604 2460
rect 18656 2448 18662 2500
rect 1104 2058 21620 2080
rect 1104 2006 4414 2058
rect 4466 2006 4478 2058
rect 4530 2006 4542 2058
rect 4594 2006 4606 2058
rect 4658 2006 11278 2058
rect 11330 2006 11342 2058
rect 11394 2006 11406 2058
rect 11458 2006 11470 2058
rect 11522 2006 18142 2058
rect 18194 2006 18206 2058
rect 18258 2006 18270 2058
rect 18322 2006 18334 2058
rect 18386 2006 21620 2058
rect 1104 1984 21620 2006
rect 17034 1156 17040 1208
rect 17092 1196 17098 1208
rect 19058 1196 19064 1208
rect 17092 1168 19064 1196
rect 17092 1156 17098 1168
rect 19058 1156 19064 1168
rect 19116 1156 19122 1208
<< via1 >>
rect 7846 19958 7898 20010
rect 7910 19958 7962 20010
rect 7974 19958 8026 20010
rect 8038 19958 8090 20010
rect 14710 19958 14762 20010
rect 14774 19958 14826 20010
rect 14838 19958 14890 20010
rect 14902 19958 14954 20010
rect 4712 19856 4764 19908
rect 17960 19856 18012 19908
rect 18696 19856 18748 19908
rect 20628 19856 20680 19908
rect 9588 19720 9640 19772
rect 17684 19763 17736 19772
rect 17684 19729 17693 19763
rect 17693 19729 17727 19763
rect 17727 19729 17736 19763
rect 17684 19720 17736 19729
rect 18512 19720 18564 19772
rect 19432 19720 19484 19772
rect 19708 19720 19760 19772
rect 5172 19695 5224 19704
rect 5172 19661 5181 19695
rect 5181 19661 5215 19695
rect 5215 19661 5224 19695
rect 5172 19652 5224 19661
rect 19800 19695 19852 19704
rect 19800 19661 19809 19695
rect 19809 19661 19843 19695
rect 19843 19661 19852 19695
rect 19800 19652 19852 19661
rect 5264 19516 5316 19568
rect 4414 19414 4466 19466
rect 4478 19414 4530 19466
rect 4542 19414 4594 19466
rect 4606 19414 4658 19466
rect 11278 19414 11330 19466
rect 11342 19414 11394 19466
rect 11406 19414 11458 19466
rect 11470 19414 11522 19466
rect 18142 19414 18194 19466
rect 18206 19414 18258 19466
rect 18270 19414 18322 19466
rect 18334 19414 18386 19466
rect 11060 19355 11112 19364
rect 11060 19321 11069 19355
rect 11069 19321 11103 19355
rect 11103 19321 11112 19355
rect 11060 19312 11112 19321
rect 2412 19108 2464 19160
rect 4344 19151 4396 19160
rect 4344 19117 4378 19151
rect 4378 19117 4396 19151
rect 4344 19108 4396 19117
rect 5172 19108 5224 19160
rect 6552 19108 6604 19160
rect 1952 19040 2004 19092
rect 5448 19015 5500 19024
rect 5448 18981 5457 19015
rect 5457 18981 5491 19015
rect 5491 18981 5500 19015
rect 5448 18972 5500 18981
rect 5816 19040 5868 19092
rect 8208 19040 8260 19092
rect 15384 19176 15436 19228
rect 17684 19176 17736 19228
rect 6736 18972 6788 19024
rect 6828 18972 6880 19024
rect 9036 18972 9088 19024
rect 9496 18972 9548 19024
rect 9772 19040 9824 19092
rect 9956 19083 10008 19092
rect 9956 19049 9990 19083
rect 9990 19049 10008 19083
rect 9956 19040 10008 19049
rect 10232 19040 10284 19092
rect 16764 19108 16816 19160
rect 18880 19108 18932 19160
rect 19524 19151 19576 19160
rect 19524 19117 19533 19151
rect 19533 19117 19567 19151
rect 19567 19117 19576 19151
rect 19524 19108 19576 19117
rect 12624 19083 12676 19092
rect 12624 19049 12658 19083
rect 12658 19049 12676 19083
rect 18788 19083 18840 19092
rect 12624 19040 12676 19049
rect 18788 19049 18797 19083
rect 18797 19049 18831 19083
rect 18831 19049 18840 19083
rect 18788 19040 18840 19049
rect 10968 18972 11020 19024
rect 11152 18972 11204 19024
rect 11704 19015 11756 19024
rect 11704 18981 11713 19015
rect 11713 18981 11747 19015
rect 11747 18981 11756 19015
rect 11704 18972 11756 18981
rect 11796 19015 11848 19024
rect 11796 18981 11805 19015
rect 11805 18981 11839 19015
rect 11839 18981 11848 19015
rect 11796 18972 11848 18981
rect 12716 18972 12768 19024
rect 13452 18972 13504 19024
rect 13728 19015 13780 19024
rect 13728 18981 13737 19015
rect 13737 18981 13771 19015
rect 13771 18981 13780 19015
rect 13728 18972 13780 18981
rect 14004 19015 14056 19024
rect 14004 18981 14013 19015
rect 14013 18981 14047 19015
rect 14047 18981 14056 19015
rect 14004 18972 14056 18981
rect 15568 18972 15620 19024
rect 15752 18972 15804 19024
rect 15844 18972 15896 19024
rect 19616 19040 19668 19092
rect 19248 18972 19300 19024
rect 7846 18870 7898 18922
rect 7910 18870 7962 18922
rect 7974 18870 8026 18922
rect 8038 18870 8090 18922
rect 14710 18870 14762 18922
rect 14774 18870 14826 18922
rect 14838 18870 14890 18922
rect 14902 18870 14954 18922
rect 2504 18768 2556 18820
rect 2872 18700 2924 18752
rect 4344 18768 4396 18820
rect 5264 18811 5316 18820
rect 5264 18777 5273 18811
rect 5273 18777 5307 18811
rect 5307 18777 5316 18811
rect 5264 18768 5316 18777
rect 8208 18811 8260 18820
rect 2412 18675 2464 18684
rect 2412 18641 2421 18675
rect 2421 18641 2455 18675
rect 2455 18641 2464 18675
rect 2412 18632 2464 18641
rect 7656 18632 7708 18684
rect 8208 18777 8217 18811
rect 8217 18777 8251 18811
rect 8251 18777 8260 18811
rect 8208 18768 8260 18777
rect 9128 18768 9180 18820
rect 9864 18768 9916 18820
rect 11060 18700 11112 18752
rect 14096 18768 14148 18820
rect 16764 18811 16816 18820
rect 13728 18743 13780 18752
rect 13728 18709 13762 18743
rect 13762 18709 13780 18743
rect 13728 18700 13780 18709
rect 13912 18700 13964 18752
rect 14556 18700 14608 18752
rect 16764 18777 16773 18811
rect 16773 18777 16807 18811
rect 16807 18777 16816 18811
rect 16764 18768 16816 18777
rect 16948 18768 17000 18820
rect 15384 18743 15436 18752
rect 15384 18709 15418 18743
rect 15418 18709 15436 18743
rect 15384 18700 15436 18709
rect 15568 18700 15620 18752
rect 17960 18768 18012 18820
rect 19340 18768 19392 18820
rect 19800 18768 19852 18820
rect 20720 18811 20772 18820
rect 20720 18777 20729 18811
rect 20729 18777 20763 18811
rect 20763 18777 20772 18811
rect 20720 18768 20772 18777
rect 8852 18632 8904 18684
rect 9588 18675 9640 18684
rect 9588 18641 9597 18675
rect 9597 18641 9631 18675
rect 9631 18641 9640 18675
rect 9588 18632 9640 18641
rect 9864 18632 9916 18684
rect 12808 18675 12860 18684
rect 12808 18641 12817 18675
rect 12817 18641 12851 18675
rect 12851 18641 12860 18675
rect 12808 18632 12860 18641
rect 16580 18632 16632 18684
rect 17960 18632 18012 18684
rect 18512 18700 18564 18752
rect 21456 18700 21508 18752
rect 5448 18607 5500 18616
rect 5448 18573 5457 18607
rect 5457 18573 5491 18607
rect 5491 18573 5500 18607
rect 5448 18564 5500 18573
rect 6552 18564 6604 18616
rect 7932 18564 7984 18616
rect 9496 18564 9548 18616
rect 9956 18564 10008 18616
rect 13452 18607 13504 18616
rect 7840 18496 7892 18548
rect 10600 18496 10652 18548
rect 12624 18496 12676 18548
rect 13452 18573 13461 18607
rect 13461 18573 13495 18607
rect 13495 18573 13504 18607
rect 13452 18564 13504 18573
rect 296 18428 348 18480
rect 3516 18428 3568 18480
rect 3608 18428 3660 18480
rect 4252 18428 4304 18480
rect 5264 18428 5316 18480
rect 7472 18428 7524 18480
rect 8484 18428 8536 18480
rect 11796 18428 11848 18480
rect 12440 18471 12492 18480
rect 12440 18437 12449 18471
rect 12449 18437 12483 18471
rect 12483 18437 12492 18471
rect 12440 18428 12492 18437
rect 16488 18564 16540 18616
rect 19708 18607 19760 18616
rect 19708 18573 19717 18607
rect 19717 18573 19751 18607
rect 19751 18573 19760 18607
rect 19708 18564 19760 18573
rect 19892 18564 19944 18616
rect 16396 18496 16448 18548
rect 20536 18496 20588 18548
rect 16488 18471 16540 18480
rect 16488 18437 16497 18471
rect 16497 18437 16531 18471
rect 16531 18437 16540 18471
rect 16488 18428 16540 18437
rect 17500 18428 17552 18480
rect 21180 18428 21232 18480
rect 4414 18326 4466 18378
rect 4478 18326 4530 18378
rect 4542 18326 4594 18378
rect 4606 18326 4658 18378
rect 11278 18326 11330 18378
rect 11342 18326 11394 18378
rect 11406 18326 11458 18378
rect 11470 18326 11522 18378
rect 18142 18326 18194 18378
rect 18206 18326 18258 18378
rect 18270 18326 18322 18378
rect 18334 18326 18386 18378
rect 6920 18224 6972 18276
rect 7656 18156 7708 18208
rect 11152 18224 11204 18276
rect 3516 18088 3568 18140
rect 7840 18088 7892 18140
rect 8208 18088 8260 18140
rect 8576 18088 8628 18140
rect 11704 18088 11756 18140
rect 19524 18156 19576 18208
rect 19984 18224 20036 18276
rect 19892 18156 19944 18208
rect 5264 18063 5316 18072
rect 5264 18029 5273 18063
rect 5273 18029 5307 18063
rect 5307 18029 5316 18063
rect 5264 18020 5316 18029
rect 7932 18020 7984 18072
rect 8392 18020 8444 18072
rect 9588 18020 9640 18072
rect 11888 18020 11940 18072
rect 12440 18020 12492 18072
rect 14096 18088 14148 18140
rect 16580 18131 16632 18140
rect 16580 18097 16589 18131
rect 16589 18097 16623 18131
rect 16623 18097 16632 18131
rect 16580 18088 16632 18097
rect 19156 18088 19208 18140
rect 20168 18088 20220 18140
rect 16856 18020 16908 18072
rect 19524 18063 19576 18072
rect 19524 18029 19533 18063
rect 19533 18029 19567 18063
rect 19567 18029 19576 18063
rect 19524 18020 19576 18029
rect 19800 18020 19852 18072
rect 21364 18020 21416 18072
rect 5540 17995 5592 18004
rect 5540 17961 5549 17995
rect 5549 17961 5583 17995
rect 5583 17961 5592 17995
rect 5540 17952 5592 17961
rect 3056 17884 3108 17936
rect 5908 17884 5960 17936
rect 8852 17884 8904 17936
rect 11704 17884 11756 17936
rect 12532 17884 12584 17936
rect 12992 17884 13044 17936
rect 14004 17952 14056 18004
rect 19432 17952 19484 18004
rect 21088 17952 21140 18004
rect 22468 17952 22520 18004
rect 14188 17884 14240 17936
rect 15016 17884 15068 17936
rect 15292 17884 15344 17936
rect 16396 17884 16448 17936
rect 19616 17884 19668 17936
rect 20260 17884 20312 17936
rect 20628 17884 20680 17936
rect 21916 17884 21968 17936
rect 7846 17782 7898 17834
rect 7910 17782 7962 17834
rect 7974 17782 8026 17834
rect 8038 17782 8090 17834
rect 14710 17782 14762 17834
rect 14774 17782 14826 17834
rect 14838 17782 14890 17834
rect 14902 17782 14954 17834
rect 2872 17723 2924 17732
rect 2872 17689 2881 17723
rect 2881 17689 2915 17723
rect 2915 17689 2924 17723
rect 2872 17680 2924 17689
rect 4068 17680 4120 17732
rect 12348 17680 12400 17732
rect 20444 17723 20496 17732
rect 20444 17689 20453 17723
rect 20453 17689 20487 17723
rect 20487 17689 20496 17723
rect 20444 17680 20496 17689
rect 20996 17723 21048 17732
rect 20996 17689 21005 17723
rect 21005 17689 21039 17723
rect 21039 17689 21048 17723
rect 20996 17680 21048 17689
rect 1676 17612 1728 17664
rect 2412 17612 2464 17664
rect 5448 17612 5500 17664
rect 3148 17544 3200 17596
rect 5540 17544 5592 17596
rect 20260 17587 20312 17596
rect 20260 17553 20269 17587
rect 20269 17553 20303 17587
rect 20303 17553 20312 17587
rect 20260 17544 20312 17553
rect 20352 17544 20404 17596
rect 3332 17519 3384 17528
rect 3332 17485 3341 17519
rect 3341 17485 3375 17519
rect 3375 17485 3384 17519
rect 3332 17476 3384 17485
rect 10784 17476 10836 17528
rect 17040 17476 17092 17528
rect 6920 17408 6972 17460
rect 18696 17408 18748 17460
rect 5724 17340 5776 17392
rect 9128 17340 9180 17392
rect 12348 17340 12400 17392
rect 17868 17340 17920 17392
rect 19892 17383 19944 17392
rect 19892 17349 19901 17383
rect 19901 17349 19935 17383
rect 19935 17349 19944 17383
rect 19892 17340 19944 17349
rect 21732 17315 21784 17324
rect 4414 17238 4466 17290
rect 4478 17238 4530 17290
rect 4542 17238 4594 17290
rect 4606 17238 4658 17290
rect 11278 17238 11330 17290
rect 11342 17238 11394 17290
rect 11406 17238 11458 17290
rect 11470 17238 11522 17290
rect 18142 17238 18194 17290
rect 18206 17238 18258 17290
rect 18270 17238 18322 17290
rect 18334 17238 18386 17290
rect 21732 17281 21741 17315
rect 21741 17281 21775 17315
rect 21775 17281 21784 17315
rect 21732 17272 21784 17281
rect 7656 17136 7708 17188
rect 15752 17136 15804 17188
rect 17868 17179 17920 17188
rect 17868 17145 17877 17179
rect 17877 17145 17911 17179
rect 17911 17145 17920 17179
rect 17868 17136 17920 17145
rect 17960 17136 18012 17188
rect 3148 17068 3200 17120
rect 2872 17000 2924 17052
rect 4160 17000 4212 17052
rect 5632 17000 5684 17052
rect 9128 17043 9180 17052
rect 3332 16975 3384 16984
rect 3332 16941 3341 16975
rect 3341 16941 3375 16975
rect 3375 16941 3384 16975
rect 3332 16932 3384 16941
rect 5724 16932 5776 16984
rect 6552 16975 6604 16984
rect 6552 16941 6561 16975
rect 6561 16941 6595 16975
rect 6595 16941 6604 16975
rect 6552 16932 6604 16941
rect 9128 17009 9137 17043
rect 9137 17009 9171 17043
rect 9171 17009 9180 17043
rect 9128 17000 9180 17009
rect 10416 17043 10468 17052
rect 10416 17009 10425 17043
rect 10425 17009 10459 17043
rect 10459 17009 10468 17043
rect 10416 17000 10468 17009
rect 12348 17043 12400 17052
rect 12348 17009 12357 17043
rect 12357 17009 12391 17043
rect 12391 17009 12400 17043
rect 12348 17000 12400 17009
rect 12900 17000 12952 17052
rect 10968 16932 11020 16984
rect 12808 16932 12860 16984
rect 14188 16932 14240 16984
rect 15568 16932 15620 16984
rect 20260 17043 20312 17052
rect 20260 17009 20269 17043
rect 20269 17009 20303 17043
rect 20303 17009 20312 17043
rect 20260 17000 20312 17009
rect 19984 16975 20036 16984
rect 19984 16941 19993 16975
rect 19993 16941 20027 16975
rect 20027 16941 20036 16975
rect 19984 16932 20036 16941
rect 7104 16864 7156 16916
rect 2964 16839 3016 16848
rect 2964 16805 2973 16839
rect 2973 16805 3007 16839
rect 3007 16805 3016 16839
rect 2964 16796 3016 16805
rect 8392 16796 8444 16848
rect 8944 16839 8996 16848
rect 8944 16805 8953 16839
rect 8953 16805 8987 16839
rect 8987 16805 8996 16839
rect 8944 16796 8996 16805
rect 10140 16839 10192 16848
rect 10140 16805 10149 16839
rect 10149 16805 10183 16839
rect 10183 16805 10192 16839
rect 10140 16796 10192 16805
rect 16948 16864 17000 16916
rect 17960 16864 18012 16916
rect 20536 16864 20588 16916
rect 12808 16839 12860 16848
rect 12808 16805 12817 16839
rect 12817 16805 12851 16839
rect 12851 16805 12860 16839
rect 12808 16796 12860 16805
rect 13176 16839 13228 16848
rect 13176 16805 13185 16839
rect 13185 16805 13219 16839
rect 13219 16805 13228 16839
rect 13176 16796 13228 16805
rect 18052 16796 18104 16848
rect 7846 16694 7898 16746
rect 7910 16694 7962 16746
rect 7974 16694 8026 16746
rect 8038 16694 8090 16746
rect 14710 16694 14762 16746
rect 14774 16694 14826 16746
rect 14838 16694 14890 16746
rect 14902 16694 14954 16746
rect 6920 16635 6972 16644
rect 6920 16601 6929 16635
rect 6929 16601 6963 16635
rect 6963 16601 6972 16635
rect 6920 16592 6972 16601
rect 11796 16635 11848 16644
rect 6552 16524 6604 16576
rect 2964 16456 3016 16508
rect 9128 16524 9180 16576
rect 11796 16601 11805 16635
rect 11805 16601 11839 16635
rect 11839 16601 11848 16635
rect 11796 16592 11848 16601
rect 12348 16592 12400 16644
rect 12808 16592 12860 16644
rect 16948 16635 17000 16644
rect 10416 16524 10468 16576
rect 9772 16456 9824 16508
rect 4160 16431 4212 16440
rect 4160 16397 4169 16431
rect 4169 16397 4203 16431
rect 4203 16397 4212 16431
rect 4160 16388 4212 16397
rect 7380 16431 7432 16440
rect 7380 16397 7389 16431
rect 7389 16397 7423 16431
rect 7423 16397 7432 16431
rect 7380 16388 7432 16397
rect 7104 16320 7156 16372
rect 12716 16388 12768 16440
rect 15568 16524 15620 16576
rect 16488 16524 16540 16576
rect 16948 16601 16957 16635
rect 16957 16601 16991 16635
rect 16991 16601 17000 16635
rect 16948 16592 17000 16601
rect 18052 16635 18104 16644
rect 18052 16601 18061 16635
rect 18061 16601 18095 16635
rect 18095 16601 18104 16635
rect 18052 16592 18104 16601
rect 12900 16456 12952 16508
rect 15476 16456 15528 16508
rect 18696 16499 18748 16508
rect 18696 16465 18705 16499
rect 18705 16465 18739 16499
rect 18739 16465 18748 16499
rect 18696 16456 18748 16465
rect 19524 16524 19576 16576
rect 20352 16524 20404 16576
rect 20536 16499 20588 16508
rect 20536 16465 20545 16499
rect 20545 16465 20579 16499
rect 20579 16465 20588 16499
rect 20536 16456 20588 16465
rect 14372 16295 14424 16304
rect 14372 16261 14381 16295
rect 14381 16261 14415 16295
rect 14415 16261 14424 16295
rect 14372 16252 14424 16261
rect 4414 16150 4466 16202
rect 4478 16150 4530 16202
rect 4542 16150 4594 16202
rect 4606 16150 4658 16202
rect 11278 16150 11330 16202
rect 11342 16150 11394 16202
rect 11406 16150 11458 16202
rect 11470 16150 11522 16202
rect 18142 16150 18194 16202
rect 18206 16150 18258 16202
rect 18270 16150 18322 16202
rect 18334 16150 18386 16202
rect 3148 16091 3200 16100
rect 3148 16057 3157 16091
rect 3157 16057 3191 16091
rect 3191 16057 3200 16091
rect 3148 16048 3200 16057
rect 4160 16048 4212 16100
rect 7104 16091 7156 16100
rect 7104 16057 7113 16091
rect 7113 16057 7147 16091
rect 7147 16057 7156 16091
rect 7104 16048 7156 16057
rect 7380 16091 7432 16100
rect 7380 16057 7389 16091
rect 7389 16057 7423 16091
rect 7423 16057 7432 16091
rect 7380 16048 7432 16057
rect 12900 16091 12952 16100
rect 12900 16057 12909 16091
rect 12909 16057 12943 16091
rect 12943 16057 12952 16091
rect 12900 16048 12952 16057
rect 17960 16048 18012 16100
rect 20444 16091 20496 16100
rect 20444 16057 20453 16091
rect 20453 16057 20487 16091
rect 20487 16057 20496 16091
rect 20444 16048 20496 16057
rect 1676 15912 1728 15964
rect 7748 15912 7800 15964
rect 10140 15955 10192 15964
rect 3884 15844 3936 15896
rect 5724 15887 5776 15896
rect 5724 15853 5733 15887
rect 5733 15853 5767 15887
rect 5767 15853 5776 15887
rect 5724 15844 5776 15853
rect 10140 15921 10149 15955
rect 10149 15921 10183 15955
rect 10183 15921 10192 15955
rect 10140 15912 10192 15921
rect 13176 15955 13228 15964
rect 13176 15921 13185 15955
rect 13185 15921 13219 15955
rect 13219 15921 13228 15955
rect 13176 15912 13228 15921
rect 14372 15912 14424 15964
rect 15844 15955 15896 15964
rect 15844 15921 15853 15955
rect 15853 15921 15887 15955
rect 15887 15921 15896 15955
rect 15844 15912 15896 15921
rect 16948 15912 17000 15964
rect 11060 15844 11112 15896
rect 11796 15887 11848 15896
rect 11796 15853 11830 15887
rect 11830 15853 11848 15887
rect 11796 15844 11848 15853
rect 2964 15776 3016 15828
rect 6184 15776 6236 15828
rect 9036 15776 9088 15828
rect 15476 15844 15528 15896
rect 17040 15887 17092 15896
rect 17040 15853 17049 15887
rect 17049 15853 17083 15887
rect 17083 15853 17092 15887
rect 17040 15844 17092 15853
rect 18880 15887 18932 15896
rect 18880 15853 18889 15887
rect 18889 15853 18923 15887
rect 18923 15853 18932 15887
rect 18880 15844 18932 15853
rect 7748 15751 7800 15760
rect 7748 15717 7757 15751
rect 7757 15717 7791 15751
rect 7791 15717 7800 15751
rect 7748 15708 7800 15717
rect 19984 15844 20036 15896
rect 14464 15751 14516 15760
rect 14464 15717 14473 15751
rect 14473 15717 14507 15751
rect 14507 15717 14516 15751
rect 14464 15708 14516 15717
rect 20168 15776 20220 15828
rect 16948 15751 17000 15760
rect 16948 15717 16957 15751
rect 16957 15717 16991 15751
rect 16991 15717 17000 15751
rect 16948 15708 17000 15717
rect 7846 15606 7898 15658
rect 7910 15606 7962 15658
rect 7974 15606 8026 15658
rect 8038 15606 8090 15658
rect 14710 15606 14762 15658
rect 14774 15606 14826 15658
rect 14838 15606 14890 15658
rect 14902 15606 14954 15658
rect 2964 15547 3016 15556
rect 2964 15513 2973 15547
rect 2973 15513 3007 15547
rect 3007 15513 3016 15547
rect 2964 15504 3016 15513
rect 6184 15547 6236 15556
rect 1676 15368 1728 15420
rect 6184 15513 6193 15547
rect 6193 15513 6227 15547
rect 6227 15513 6236 15547
rect 6184 15504 6236 15513
rect 14464 15504 14516 15556
rect 16948 15504 17000 15556
rect 19248 15504 19300 15556
rect 21272 15504 21324 15556
rect 18880 15436 18932 15488
rect 6828 15368 6880 15420
rect 8208 15368 8260 15420
rect 15108 15368 15160 15420
rect 19984 15411 20036 15420
rect 19984 15377 19993 15411
rect 19993 15377 20027 15411
rect 20027 15377 20036 15411
rect 19984 15368 20036 15377
rect 3700 15343 3752 15352
rect 3700 15309 3709 15343
rect 3709 15309 3743 15343
rect 3743 15309 3752 15343
rect 3700 15300 3752 15309
rect 3884 15300 3936 15352
rect 3608 15164 3660 15216
rect 5724 15164 5776 15216
rect 10048 15164 10100 15216
rect 18788 15164 18840 15216
rect 19524 15164 19576 15216
rect 19800 15164 19852 15216
rect 4414 15062 4466 15114
rect 4478 15062 4530 15114
rect 4542 15062 4594 15114
rect 4606 15062 4658 15114
rect 11278 15062 11330 15114
rect 11342 15062 11394 15114
rect 11406 15062 11458 15114
rect 11470 15062 11522 15114
rect 18142 15062 18194 15114
rect 18206 15062 18258 15114
rect 18270 15062 18322 15114
rect 18334 15062 18386 15114
rect 3700 14960 3752 15012
rect 15108 14960 15160 15012
rect 19892 15003 19944 15012
rect 19892 14969 19901 15003
rect 19901 14969 19935 15003
rect 19935 14969 19944 15003
rect 19892 14960 19944 14969
rect 20444 15003 20496 15012
rect 20444 14969 20453 15003
rect 20453 14969 20487 15003
rect 20487 14969 20496 15003
rect 20444 14960 20496 14969
rect 3608 14824 3660 14876
rect 8484 14867 8536 14876
rect 8484 14833 8493 14867
rect 8493 14833 8527 14867
rect 8527 14833 8536 14867
rect 8484 14824 8536 14833
rect 8668 14867 8720 14876
rect 8668 14833 8677 14867
rect 8677 14833 8711 14867
rect 8711 14833 8720 14867
rect 8668 14824 8720 14833
rect 10968 14892 11020 14944
rect 12716 14892 12768 14944
rect 10232 14867 10284 14876
rect 10232 14833 10241 14867
rect 10241 14833 10275 14867
rect 10275 14833 10284 14867
rect 10232 14824 10284 14833
rect 11704 14824 11756 14876
rect 15200 14892 15252 14944
rect 15844 14892 15896 14944
rect 17040 14867 17092 14876
rect 4252 14756 4304 14808
rect 7748 14756 7800 14808
rect 12164 14756 12216 14808
rect 12348 14756 12400 14808
rect 13360 14799 13412 14808
rect 13360 14765 13369 14799
rect 13369 14765 13403 14799
rect 13403 14765 13412 14799
rect 13360 14756 13412 14765
rect 17040 14833 17049 14867
rect 17049 14833 17083 14867
rect 17083 14833 17092 14867
rect 17040 14824 17092 14833
rect 19984 14824 20036 14876
rect 14372 14756 14424 14808
rect 13728 14688 13780 14740
rect 8392 14663 8444 14672
rect 8392 14629 8401 14663
rect 8401 14629 8435 14663
rect 8435 14629 8444 14663
rect 8392 14620 8444 14629
rect 11980 14663 12032 14672
rect 11980 14629 11989 14663
rect 11989 14629 12023 14663
rect 12023 14629 12032 14663
rect 11980 14620 12032 14629
rect 12072 14620 12124 14672
rect 19708 14799 19760 14808
rect 19708 14765 19717 14799
rect 19717 14765 19751 14799
rect 19751 14765 19760 14799
rect 19708 14756 19760 14765
rect 20168 14756 20220 14808
rect 17408 14688 17460 14740
rect 16948 14663 17000 14672
rect 16948 14629 16957 14663
rect 16957 14629 16991 14663
rect 16991 14629 17000 14663
rect 16948 14620 17000 14629
rect 7846 14518 7898 14570
rect 7910 14518 7962 14570
rect 7974 14518 8026 14570
rect 8038 14518 8090 14570
rect 14710 14518 14762 14570
rect 14774 14518 14826 14570
rect 14838 14518 14890 14570
rect 14902 14518 14954 14570
rect 6828 14416 6880 14468
rect 10232 14416 10284 14468
rect 11980 14416 12032 14468
rect 12256 14348 12308 14400
rect 3884 14323 3936 14332
rect 3884 14289 3893 14323
rect 3893 14289 3927 14323
rect 3927 14289 3936 14323
rect 3884 14280 3936 14289
rect 6092 14323 6144 14332
rect 6092 14289 6101 14323
rect 6101 14289 6135 14323
rect 6135 14289 6144 14323
rect 6092 14280 6144 14289
rect 8668 14323 8720 14332
rect 8668 14289 8702 14323
rect 8702 14289 8720 14323
rect 8668 14280 8720 14289
rect 12624 14280 12676 14332
rect 6184 14255 6236 14264
rect 6184 14221 6193 14255
rect 6193 14221 6227 14255
rect 6227 14221 6236 14255
rect 6184 14212 6236 14221
rect 6276 14255 6328 14264
rect 6276 14221 6285 14255
rect 6285 14221 6319 14255
rect 6319 14221 6328 14255
rect 6276 14212 6328 14221
rect 7380 14212 7432 14264
rect 9956 14144 10008 14196
rect 17040 14416 17092 14468
rect 20904 14459 20956 14468
rect 20904 14425 20913 14459
rect 20913 14425 20947 14459
rect 20947 14425 20956 14459
rect 20904 14416 20956 14425
rect 15200 14348 15252 14400
rect 13820 14323 13872 14332
rect 13820 14289 13829 14323
rect 13829 14289 13863 14323
rect 13863 14289 13872 14323
rect 13820 14280 13872 14289
rect 17040 14280 17092 14332
rect 17132 14280 17184 14332
rect 17776 14212 17828 14264
rect 19708 14212 19760 14264
rect 5540 14076 5592 14128
rect 11704 14076 11756 14128
rect 4414 13974 4466 14026
rect 4478 13974 4530 14026
rect 4542 13974 4594 14026
rect 4606 13974 4658 14026
rect 11278 13974 11330 14026
rect 11342 13974 11394 14026
rect 11406 13974 11458 14026
rect 11470 13974 11522 14026
rect 18142 13974 18194 14026
rect 18206 13974 18258 14026
rect 18270 13974 18322 14026
rect 18334 13974 18386 14026
rect 2504 13872 2556 13924
rect 6276 13915 6328 13924
rect 6276 13881 6285 13915
rect 6285 13881 6319 13915
rect 6319 13881 6328 13915
rect 6276 13872 6328 13881
rect 8208 13872 8260 13924
rect 8668 13915 8720 13924
rect 8668 13881 8677 13915
rect 8677 13881 8711 13915
rect 8711 13881 8720 13915
rect 8668 13872 8720 13881
rect 3608 13847 3660 13856
rect 3608 13813 3617 13847
rect 3617 13813 3651 13847
rect 3651 13813 3660 13847
rect 3608 13804 3660 13813
rect 12256 13872 12308 13924
rect 12624 13915 12676 13924
rect 12624 13881 12633 13915
rect 12633 13881 12667 13915
rect 12667 13881 12676 13915
rect 12624 13872 12676 13881
rect 17408 13915 17460 13924
rect 6092 13736 6144 13788
rect 2504 13643 2556 13652
rect 2504 13609 2538 13643
rect 2538 13609 2556 13643
rect 5540 13668 5592 13720
rect 6276 13668 6328 13720
rect 7380 13668 7432 13720
rect 9956 13804 10008 13856
rect 16948 13804 17000 13856
rect 17408 13881 17417 13915
rect 17417 13881 17451 13915
rect 17451 13881 17460 13915
rect 17408 13872 17460 13881
rect 18604 13915 18656 13924
rect 18604 13881 18613 13915
rect 18613 13881 18647 13915
rect 18647 13881 18656 13915
rect 18604 13872 18656 13881
rect 20628 13872 20680 13924
rect 17868 13804 17920 13856
rect 11980 13736 12032 13788
rect 12348 13736 12400 13788
rect 16856 13779 16908 13788
rect 16856 13745 16865 13779
rect 16865 13745 16899 13779
rect 16899 13745 16908 13779
rect 16856 13736 16908 13745
rect 17040 13779 17092 13788
rect 17040 13745 17049 13779
rect 17049 13745 17083 13779
rect 17083 13745 17092 13779
rect 17040 13736 17092 13745
rect 20352 13736 20404 13788
rect 20628 13736 20680 13788
rect 10876 13668 10928 13720
rect 10968 13711 11020 13720
rect 10968 13677 10977 13711
rect 10977 13677 11011 13711
rect 11011 13677 11020 13711
rect 10968 13668 11020 13677
rect 11704 13668 11756 13720
rect 17132 13668 17184 13720
rect 17868 13711 17920 13720
rect 17868 13677 17877 13711
rect 17877 13677 17911 13711
rect 17911 13677 17920 13711
rect 17868 13668 17920 13677
rect 18420 13711 18472 13720
rect 18420 13677 18429 13711
rect 18429 13677 18463 13711
rect 18463 13677 18472 13711
rect 18420 13668 18472 13677
rect 20260 13711 20312 13720
rect 20260 13677 20269 13711
rect 20269 13677 20303 13711
rect 20303 13677 20312 13711
rect 20260 13668 20312 13677
rect 2504 13600 2556 13609
rect 11152 13600 11204 13652
rect 11980 13600 12032 13652
rect 17776 13643 17828 13652
rect 17776 13609 17785 13643
rect 17785 13609 17819 13643
rect 17819 13609 17828 13643
rect 17776 13600 17828 13609
rect 16764 13575 16816 13584
rect 16764 13541 16773 13575
rect 16773 13541 16807 13575
rect 16807 13541 16816 13575
rect 16764 13532 16816 13541
rect 7846 13430 7898 13482
rect 7910 13430 7962 13482
rect 7974 13430 8026 13482
rect 8038 13430 8090 13482
rect 14710 13430 14762 13482
rect 14774 13430 14826 13482
rect 14838 13430 14890 13482
rect 14902 13430 14954 13482
rect 6184 13328 6236 13380
rect 10876 13328 10928 13380
rect 19524 13328 19576 13380
rect 20168 13371 20220 13380
rect 20168 13337 20177 13371
rect 20177 13337 20211 13371
rect 20211 13337 20220 13371
rect 20168 13328 20220 13337
rect 20720 13371 20772 13380
rect 20720 13337 20729 13371
rect 20729 13337 20763 13371
rect 20763 13337 20772 13371
rect 20720 13328 20772 13337
rect 5908 13260 5960 13312
rect 10048 13303 10100 13312
rect 10048 13269 10059 13303
rect 10059 13269 10093 13303
rect 10093 13269 10100 13303
rect 10048 13260 10100 13269
rect 18420 13260 18472 13312
rect 8392 13192 8444 13244
rect 8484 13192 8536 13244
rect 14464 13192 14516 13244
rect 18696 13235 18748 13244
rect 18696 13201 18705 13235
rect 18705 13201 18739 13235
rect 18739 13201 18748 13235
rect 18696 13192 18748 13201
rect 19248 13192 19300 13244
rect 20536 13235 20588 13244
rect 6276 13167 6328 13176
rect 6276 13133 6285 13167
rect 6285 13133 6319 13167
rect 6319 13133 6328 13167
rect 6276 13124 6328 13133
rect 11704 13124 11756 13176
rect 20536 13201 20545 13235
rect 20545 13201 20579 13235
rect 20579 13201 20588 13235
rect 20536 13192 20588 13201
rect 12624 13056 12676 13108
rect 848 12988 900 13040
rect 13452 12988 13504 13040
rect 4414 12886 4466 12938
rect 4478 12886 4530 12938
rect 4542 12886 4594 12938
rect 4606 12886 4658 12938
rect 11278 12886 11330 12938
rect 11342 12886 11394 12938
rect 11406 12886 11458 12938
rect 11470 12886 11522 12938
rect 18142 12886 18194 12938
rect 18206 12886 18258 12938
rect 18270 12886 18322 12938
rect 18334 12886 18386 12938
rect 7380 12784 7432 12836
rect 7564 12827 7616 12836
rect 7564 12793 7573 12827
rect 7573 12793 7607 12827
rect 7607 12793 7616 12827
rect 7564 12784 7616 12793
rect 8392 12784 8444 12836
rect 7564 12648 7616 12700
rect 8208 12580 8260 12632
rect 10232 12555 10284 12564
rect 10232 12521 10266 12555
rect 10266 12521 10284 12555
rect 10232 12512 10284 12521
rect 11152 12784 11204 12836
rect 13360 12784 13412 12836
rect 20168 12827 20220 12836
rect 20168 12793 20177 12827
rect 20177 12793 20211 12827
rect 20211 12793 20220 12827
rect 20168 12784 20220 12793
rect 14556 12716 14608 12768
rect 11704 12691 11756 12700
rect 11704 12657 11713 12691
rect 11713 12657 11747 12691
rect 11747 12657 11756 12691
rect 11704 12648 11756 12657
rect 13452 12691 13504 12700
rect 13452 12657 13461 12691
rect 13461 12657 13495 12691
rect 13495 12657 13504 12691
rect 13452 12648 13504 12657
rect 13544 12648 13596 12700
rect 15108 12648 15160 12700
rect 15200 12648 15252 12700
rect 11428 12623 11480 12632
rect 11428 12589 11437 12623
rect 11437 12589 11471 12623
rect 11471 12589 11480 12623
rect 11428 12580 11480 12589
rect 12624 12623 12676 12632
rect 12624 12589 12641 12623
rect 12641 12589 12675 12623
rect 12675 12589 12676 12623
rect 12624 12580 12676 12589
rect 13820 12580 13872 12632
rect 20536 12648 20588 12700
rect 19156 12623 19208 12632
rect 19156 12589 19165 12623
rect 19165 12589 19199 12623
rect 19199 12589 19208 12623
rect 19156 12580 19208 12589
rect 14464 12555 14516 12564
rect 14464 12521 14473 12555
rect 14473 12521 14507 12555
rect 14507 12521 14516 12555
rect 14464 12512 14516 12521
rect 17500 12512 17552 12564
rect 13452 12444 13504 12496
rect 14004 12487 14056 12496
rect 14004 12453 14013 12487
rect 14013 12453 14047 12487
rect 14047 12453 14056 12487
rect 14004 12444 14056 12453
rect 14188 12444 14240 12496
rect 17960 12487 18012 12496
rect 17960 12453 17969 12487
rect 17969 12453 18003 12487
rect 18003 12453 18012 12487
rect 17960 12444 18012 12453
rect 7846 12342 7898 12394
rect 7910 12342 7962 12394
rect 7974 12342 8026 12394
rect 8038 12342 8090 12394
rect 14710 12342 14762 12394
rect 14774 12342 14826 12394
rect 14838 12342 14890 12394
rect 14902 12342 14954 12394
rect 8944 12240 8996 12292
rect 11428 12240 11480 12292
rect 7196 12172 7248 12224
rect 7564 12172 7616 12224
rect 14188 12240 14240 12292
rect 14556 12283 14608 12292
rect 14556 12249 14565 12283
rect 14565 12249 14599 12283
rect 14599 12249 14608 12283
rect 14556 12240 14608 12249
rect 15108 12240 15160 12292
rect 17960 12240 18012 12292
rect 19156 12240 19208 12292
rect 20996 12240 21048 12292
rect 7288 12147 7340 12156
rect 7288 12113 7322 12147
rect 7322 12113 7340 12147
rect 13544 12172 13596 12224
rect 14004 12172 14056 12224
rect 7288 12104 7340 12113
rect 10416 12104 10468 12156
rect 15200 12147 15252 12156
rect 15200 12113 15209 12147
rect 15209 12113 15243 12147
rect 15243 12113 15252 12147
rect 15200 12104 15252 12113
rect 17960 12104 18012 12156
rect 19984 12147 20036 12156
rect 9772 12036 9824 12088
rect 10232 11968 10284 12020
rect 12440 12079 12492 12088
rect 12440 12045 12449 12079
rect 12449 12045 12483 12079
rect 12483 12045 12492 12079
rect 12440 12036 12492 12045
rect 16948 12036 17000 12088
rect 19984 12113 19993 12147
rect 19993 12113 20027 12147
rect 20027 12113 20036 12147
rect 19984 12104 20036 12113
rect 20536 12147 20588 12156
rect 20536 12113 20545 12147
rect 20545 12113 20579 12147
rect 20579 12113 20588 12147
rect 20536 12104 20588 12113
rect 14280 11968 14332 12020
rect 19616 11968 19668 12020
rect 8668 11900 8720 11952
rect 14004 11900 14056 11952
rect 14188 11900 14240 11952
rect 18604 11900 18656 11952
rect 4414 11798 4466 11850
rect 4478 11798 4530 11850
rect 4542 11798 4594 11850
rect 4606 11798 4658 11850
rect 11278 11798 11330 11850
rect 11342 11798 11394 11850
rect 11406 11798 11458 11850
rect 11470 11798 11522 11850
rect 18142 11798 18194 11850
rect 18206 11798 18258 11850
rect 18270 11798 18322 11850
rect 18334 11798 18386 11850
rect 9772 11696 9824 11748
rect 10416 11739 10468 11748
rect 10416 11705 10425 11739
rect 10425 11705 10459 11739
rect 10459 11705 10468 11739
rect 10416 11696 10468 11705
rect 12440 11696 12492 11748
rect 13820 11696 13872 11748
rect 17960 11696 18012 11748
rect 20076 11696 20128 11748
rect 6828 11560 6880 11612
rect 7288 11603 7340 11612
rect 7288 11569 7297 11603
rect 7297 11569 7331 11603
rect 7331 11569 7340 11603
rect 8668 11603 8720 11612
rect 7288 11560 7340 11569
rect 8392 11492 8444 11544
rect 8668 11569 8677 11603
rect 8677 11569 8711 11603
rect 8711 11569 8720 11603
rect 8668 11560 8720 11569
rect 14372 11628 14424 11680
rect 14004 11603 14056 11612
rect 8576 11492 8628 11544
rect 14004 11569 14013 11603
rect 14013 11569 14047 11603
rect 14047 11569 14056 11603
rect 14004 11560 14056 11569
rect 14096 11603 14148 11612
rect 14096 11569 14105 11603
rect 14105 11569 14139 11603
rect 14139 11569 14148 11603
rect 14096 11560 14148 11569
rect 17500 11560 17552 11612
rect 13360 11492 13412 11544
rect 15752 11492 15804 11544
rect 19156 11492 19208 11544
rect 20260 11535 20312 11544
rect 20260 11501 20269 11535
rect 20269 11501 20303 11535
rect 20303 11501 20312 11535
rect 20260 11492 20312 11501
rect 11612 11424 11664 11476
rect 14556 11424 14608 11476
rect 8300 11356 8352 11408
rect 13728 11356 13780 11408
rect 18788 11356 18840 11408
rect 7846 11254 7898 11306
rect 7910 11254 7962 11306
rect 7974 11254 8026 11306
rect 8038 11254 8090 11306
rect 14710 11254 14762 11306
rect 14774 11254 14826 11306
rect 14838 11254 14890 11306
rect 14902 11254 14954 11306
rect 8300 11195 8352 11204
rect 8300 11161 8309 11195
rect 8309 11161 8343 11195
rect 8343 11161 8352 11195
rect 8300 11152 8352 11161
rect 8484 11152 8536 11204
rect 13728 11195 13780 11204
rect 13728 11161 13737 11195
rect 13737 11161 13771 11195
rect 13771 11161 13780 11195
rect 13728 11152 13780 11161
rect 14188 11152 14240 11204
rect 14372 11152 14424 11204
rect 18788 11195 18840 11204
rect 18788 11161 18797 11195
rect 18797 11161 18831 11195
rect 18831 11161 18840 11195
rect 18788 11152 18840 11161
rect 20628 11152 20680 11204
rect 20812 11152 20864 11204
rect 8944 11084 8996 11136
rect 10048 11016 10100 11068
rect 16764 11016 16816 11068
rect 17132 11016 17184 11068
rect 17316 11059 17368 11068
rect 17316 11025 17325 11059
rect 17325 11025 17359 11059
rect 17359 11025 17368 11059
rect 17316 11016 17368 11025
rect 17868 11016 17920 11068
rect 19984 11059 20036 11068
rect 19984 11025 19993 11059
rect 19993 11025 20027 11059
rect 20027 11025 20036 11059
rect 19984 11016 20036 11025
rect 8576 10948 8628 11000
rect 14188 10991 14240 11000
rect 14188 10957 14197 10991
rect 14197 10957 14231 10991
rect 14231 10957 14240 10991
rect 14188 10948 14240 10957
rect 14280 10991 14332 11000
rect 14280 10957 14289 10991
rect 14289 10957 14323 10991
rect 14323 10957 14332 10991
rect 14280 10948 14332 10957
rect 14556 10948 14608 11000
rect 17500 10991 17552 11000
rect 12072 10880 12124 10932
rect 16488 10880 16540 10932
rect 17500 10957 17509 10991
rect 17509 10957 17543 10991
rect 17543 10957 17552 10991
rect 17500 10948 17552 10957
rect 16948 10923 17000 10932
rect 16948 10889 16957 10923
rect 16957 10889 16991 10923
rect 16991 10889 17000 10923
rect 16948 10880 17000 10889
rect 19156 10880 19208 10932
rect 13452 10812 13504 10864
rect 18512 10812 18564 10864
rect 19248 10812 19300 10864
rect 4414 10710 4466 10762
rect 4478 10710 4530 10762
rect 4542 10710 4594 10762
rect 4606 10710 4658 10762
rect 11278 10710 11330 10762
rect 11342 10710 11394 10762
rect 11406 10710 11458 10762
rect 11470 10710 11522 10762
rect 18142 10710 18194 10762
rect 18206 10710 18258 10762
rect 18270 10710 18322 10762
rect 18334 10710 18386 10762
rect 1676 10608 1728 10660
rect 8576 10583 8628 10592
rect 8576 10549 8585 10583
rect 8585 10549 8619 10583
rect 8619 10549 8628 10583
rect 8576 10540 8628 10549
rect 11704 10608 11756 10660
rect 14096 10651 14148 10660
rect 11796 10472 11848 10524
rect 12440 10472 12492 10524
rect 12716 10515 12768 10524
rect 12716 10481 12725 10515
rect 12725 10481 12759 10515
rect 12759 10481 12768 10515
rect 12716 10472 12768 10481
rect 14096 10617 14105 10651
rect 14105 10617 14139 10651
rect 14139 10617 14148 10651
rect 14096 10608 14148 10617
rect 17316 10608 17368 10660
rect 18696 10608 18748 10660
rect 19340 10608 19392 10660
rect 16488 10540 16540 10592
rect 19248 10540 19300 10592
rect 7196 10447 7248 10456
rect 7196 10413 7205 10447
rect 7205 10413 7239 10447
rect 7239 10413 7248 10447
rect 7196 10404 7248 10413
rect 12072 10404 12124 10456
rect 14280 10404 14332 10456
rect 19340 10472 19392 10524
rect 18972 10404 19024 10456
rect 20260 10447 20312 10456
rect 20260 10413 20269 10447
rect 20269 10413 20303 10447
rect 20303 10413 20312 10447
rect 20260 10404 20312 10413
rect 9312 10336 9364 10388
rect 19708 10336 19760 10388
rect 11060 10311 11112 10320
rect 11060 10277 11069 10311
rect 11069 10277 11103 10311
rect 11103 10277 11112 10311
rect 11060 10268 11112 10277
rect 17040 10311 17092 10320
rect 17040 10277 17049 10311
rect 17049 10277 17083 10311
rect 17083 10277 17092 10311
rect 17040 10268 17092 10277
rect 18880 10311 18932 10320
rect 18880 10277 18889 10311
rect 18889 10277 18923 10311
rect 18923 10277 18932 10311
rect 18880 10268 18932 10277
rect 7846 10166 7898 10218
rect 7910 10166 7962 10218
rect 7974 10166 8026 10218
rect 8038 10166 8090 10218
rect 14710 10166 14762 10218
rect 14774 10166 14826 10218
rect 14838 10166 14890 10218
rect 14902 10166 14954 10218
rect 10048 10107 10100 10116
rect 10048 10073 10057 10107
rect 10057 10073 10091 10107
rect 10091 10073 10100 10107
rect 10048 10064 10100 10073
rect 17500 10064 17552 10116
rect 19248 10064 19300 10116
rect 21180 10064 21232 10116
rect 11612 9996 11664 10048
rect 16488 9996 16540 10048
rect 12348 9928 12400 9980
rect 15200 9928 15252 9980
rect 15936 9971 15988 9980
rect 15936 9937 15945 9971
rect 15945 9937 15979 9971
rect 15979 9937 15988 9971
rect 15936 9928 15988 9937
rect 19340 9928 19392 9980
rect 20536 9971 20588 9980
rect 20536 9937 20545 9971
rect 20545 9937 20579 9971
rect 20579 9937 20588 9971
rect 20536 9928 20588 9937
rect 10508 9903 10560 9912
rect 10508 9869 10517 9903
rect 10517 9869 10551 9903
rect 10551 9869 10560 9903
rect 10508 9860 10560 9869
rect 9312 9792 9364 9844
rect 11152 9860 11204 9912
rect 17960 9860 18012 9912
rect 4414 9622 4466 9674
rect 4478 9622 4530 9674
rect 4542 9622 4594 9674
rect 4606 9622 4658 9674
rect 11278 9622 11330 9674
rect 11342 9622 11394 9674
rect 11406 9622 11458 9674
rect 11470 9622 11522 9674
rect 18142 9622 18194 9674
rect 18206 9622 18258 9674
rect 18270 9622 18322 9674
rect 18334 9622 18386 9674
rect 10508 9563 10560 9572
rect 10508 9529 10517 9563
rect 10517 9529 10551 9563
rect 10551 9529 10560 9563
rect 10508 9520 10560 9529
rect 12348 9563 12400 9572
rect 12348 9529 12357 9563
rect 12357 9529 12391 9563
rect 12391 9529 12400 9563
rect 12348 9520 12400 9529
rect 9312 9495 9364 9504
rect 9312 9461 9321 9495
rect 9321 9461 9355 9495
rect 9355 9461 9364 9495
rect 9312 9452 9364 9461
rect 12164 9452 12216 9504
rect 17040 9520 17092 9572
rect 18880 9520 18932 9572
rect 12716 9452 12768 9504
rect 11152 9427 11204 9436
rect 11152 9393 11161 9427
rect 11161 9393 11195 9427
rect 11195 9393 11204 9427
rect 11152 9384 11204 9393
rect 11612 9384 11664 9436
rect 11796 9384 11848 9436
rect 7196 9316 7248 9368
rect 11060 9248 11112 9300
rect 12900 9248 12952 9300
rect 14096 9316 14148 9368
rect 15016 9452 15068 9504
rect 19432 9384 19484 9436
rect 19708 9427 19760 9436
rect 19708 9393 19717 9427
rect 19717 9393 19751 9427
rect 19751 9393 19760 9427
rect 19708 9384 19760 9393
rect 15292 9359 15344 9368
rect 15292 9325 15301 9359
rect 15301 9325 15335 9359
rect 15335 9325 15344 9359
rect 15292 9316 15344 9325
rect 19064 9359 19116 9368
rect 19064 9325 19073 9359
rect 19073 9325 19107 9359
rect 19107 9325 19116 9359
rect 19064 9316 19116 9325
rect 8208 9180 8260 9232
rect 10876 9223 10928 9232
rect 10876 9189 10885 9223
rect 10885 9189 10919 9223
rect 10919 9189 10928 9223
rect 10876 9180 10928 9189
rect 15752 9180 15804 9232
rect 19156 9223 19208 9232
rect 19156 9189 19165 9223
rect 19165 9189 19199 9223
rect 19199 9189 19208 9223
rect 19156 9180 19208 9189
rect 7846 9078 7898 9130
rect 7910 9078 7962 9130
rect 7974 9078 8026 9130
rect 8038 9078 8090 9130
rect 14710 9078 14762 9130
rect 14774 9078 14826 9130
rect 14838 9078 14890 9130
rect 14902 9078 14954 9130
rect 10876 8976 10928 9028
rect 12164 8976 12216 9028
rect 13268 8976 13320 9028
rect 11704 8908 11756 8960
rect 12900 8908 12952 8960
rect 17868 8976 17920 9028
rect 19340 8976 19392 9028
rect 20352 8976 20404 9028
rect 21456 8976 21508 9028
rect 15292 8908 15344 8960
rect 8208 8815 8260 8824
rect 8208 8781 8217 8815
rect 8217 8781 8251 8815
rect 8251 8781 8260 8815
rect 8208 8772 8260 8781
rect 11796 8840 11848 8892
rect 13544 8840 13596 8892
rect 16304 8840 16356 8892
rect 19432 8840 19484 8892
rect 19984 8883 20036 8892
rect 19984 8849 19993 8883
rect 19993 8849 20027 8883
rect 20027 8849 20036 8883
rect 19984 8840 20036 8849
rect 20536 8883 20588 8892
rect 20536 8849 20545 8883
rect 20545 8849 20579 8883
rect 20579 8849 20588 8883
rect 20536 8840 20588 8849
rect 17960 8772 18012 8824
rect 11152 8704 11204 8756
rect 4414 8534 4466 8586
rect 4478 8534 4530 8586
rect 4542 8534 4594 8586
rect 4606 8534 4658 8586
rect 11278 8534 11330 8586
rect 11342 8534 11394 8586
rect 11406 8534 11458 8586
rect 11470 8534 11522 8586
rect 18142 8534 18194 8586
rect 18206 8534 18258 8586
rect 18270 8534 18322 8586
rect 18334 8534 18386 8586
rect 11888 8432 11940 8484
rect 16304 8475 16356 8484
rect 16304 8441 16313 8475
rect 16313 8441 16347 8475
rect 16347 8441 16356 8475
rect 16304 8432 16356 8441
rect 19800 8432 19852 8484
rect 13544 8339 13596 8348
rect 13544 8305 13553 8339
rect 13553 8305 13587 8339
rect 13587 8305 13596 8339
rect 13544 8296 13596 8305
rect 17684 8296 17736 8348
rect 11336 8271 11388 8280
rect 11336 8237 11345 8271
rect 11345 8237 11379 8271
rect 11379 8237 11388 8271
rect 11336 8228 11388 8237
rect 13360 8271 13412 8280
rect 13360 8237 13369 8271
rect 13369 8237 13403 8271
rect 13403 8237 13412 8271
rect 13360 8228 13412 8237
rect 20260 8271 20312 8280
rect 20260 8237 20269 8271
rect 20269 8237 20303 8271
rect 20303 8237 20312 8271
rect 20260 8228 20312 8237
rect 10692 8135 10744 8144
rect 10692 8101 10701 8135
rect 10701 8101 10735 8135
rect 10735 8101 10744 8135
rect 10692 8092 10744 8101
rect 16764 8135 16816 8144
rect 16764 8101 16773 8135
rect 16773 8101 16807 8135
rect 16807 8101 16816 8135
rect 16764 8092 16816 8101
rect 7846 7990 7898 8042
rect 7910 7990 7962 8042
rect 7974 7990 8026 8042
rect 8038 7990 8090 8042
rect 14710 7990 14762 8042
rect 14774 7990 14826 8042
rect 14838 7990 14890 8042
rect 14902 7990 14954 8042
rect 10692 7888 10744 7940
rect 13360 7888 13412 7940
rect 11336 7820 11388 7872
rect 16672 7888 16724 7940
rect 17684 7931 17736 7940
rect 17684 7897 17693 7931
rect 17693 7897 17727 7931
rect 17727 7897 17736 7931
rect 17684 7888 17736 7897
rect 19432 7931 19484 7940
rect 19432 7897 19441 7931
rect 19441 7897 19475 7931
rect 19475 7897 19484 7931
rect 19432 7888 19484 7897
rect 16856 7820 16908 7872
rect 14648 7752 14700 7804
rect 15936 7752 15988 7804
rect 19984 7795 20036 7804
rect 10876 7727 10928 7736
rect 10876 7693 10885 7727
rect 10885 7693 10919 7727
rect 10919 7693 10928 7727
rect 10876 7684 10928 7693
rect 11060 7727 11112 7736
rect 11060 7693 11069 7727
rect 11069 7693 11103 7727
rect 11103 7693 11112 7727
rect 11060 7684 11112 7693
rect 14188 7727 14240 7736
rect 14188 7693 14197 7727
rect 14197 7693 14231 7727
rect 14231 7693 14240 7727
rect 14188 7684 14240 7693
rect 14372 7727 14424 7736
rect 14372 7693 14381 7727
rect 14381 7693 14415 7727
rect 14415 7693 14424 7727
rect 14372 7684 14424 7693
rect 17960 7684 18012 7736
rect 19984 7761 19993 7795
rect 19993 7761 20027 7795
rect 20027 7761 20036 7795
rect 19984 7752 20036 7761
rect 20536 7795 20588 7804
rect 20536 7761 20545 7795
rect 20545 7761 20579 7795
rect 20579 7761 20588 7795
rect 20536 7752 20588 7761
rect 13912 7548 13964 7600
rect 4414 7446 4466 7498
rect 4478 7446 4530 7498
rect 4542 7446 4594 7498
rect 4606 7446 4658 7498
rect 11278 7446 11330 7498
rect 11342 7446 11394 7498
rect 11406 7446 11458 7498
rect 11470 7446 11522 7498
rect 18142 7446 18194 7498
rect 18206 7446 18258 7498
rect 18270 7446 18322 7498
rect 18334 7446 18386 7498
rect 11060 7387 11112 7396
rect 11060 7353 11069 7387
rect 11069 7353 11103 7387
rect 11103 7353 11112 7387
rect 11060 7344 11112 7353
rect 16672 7387 16724 7396
rect 16672 7353 16681 7387
rect 16681 7353 16715 7387
rect 16715 7353 16724 7387
rect 16672 7344 16724 7353
rect 16764 7344 16816 7396
rect 7380 7140 7432 7192
rect 8208 7140 8260 7192
rect 9864 7072 9916 7124
rect 14372 7319 14424 7328
rect 14372 7285 14381 7319
rect 14381 7285 14415 7319
rect 14415 7285 14424 7319
rect 14372 7276 14424 7285
rect 14648 7251 14700 7260
rect 14648 7217 14657 7251
rect 14657 7217 14691 7251
rect 14691 7217 14700 7251
rect 14648 7208 14700 7217
rect 12716 7140 12768 7192
rect 14556 7140 14608 7192
rect 15936 7140 15988 7192
rect 17408 7183 17460 7192
rect 17408 7149 17417 7183
rect 17417 7149 17451 7183
rect 17451 7149 17460 7183
rect 17408 7140 17460 7149
rect 19156 7140 19208 7192
rect 18512 7072 18564 7124
rect 7846 6902 7898 6954
rect 7910 6902 7962 6954
rect 7974 6902 8026 6954
rect 8038 6902 8090 6954
rect 14710 6902 14762 6954
rect 14774 6902 14826 6954
rect 14838 6902 14890 6954
rect 14902 6902 14954 6954
rect 10876 6800 10928 6852
rect 14188 6800 14240 6852
rect 16488 6800 16540 6852
rect 4068 6664 4120 6716
rect 10600 6664 10652 6716
rect 7380 6639 7432 6648
rect 7380 6605 7389 6639
rect 7389 6605 7423 6639
rect 7423 6605 7432 6639
rect 7380 6596 7432 6605
rect 9864 6528 9916 6580
rect 14648 6639 14700 6648
rect 14648 6605 14657 6639
rect 14657 6605 14691 6639
rect 14691 6605 14700 6639
rect 18604 6664 18656 6716
rect 20536 6707 20588 6716
rect 20536 6673 20545 6707
rect 20545 6673 20579 6707
rect 20579 6673 20588 6707
rect 20536 6664 20588 6673
rect 14648 6596 14700 6605
rect 17408 6596 17460 6648
rect 13636 6528 13688 6580
rect 4414 6358 4466 6410
rect 4478 6358 4530 6410
rect 4542 6358 4594 6410
rect 4606 6358 4658 6410
rect 11278 6358 11330 6410
rect 11342 6358 11394 6410
rect 11406 6358 11458 6410
rect 11470 6358 11522 6410
rect 18142 6358 18194 6410
rect 18206 6358 18258 6410
rect 18270 6358 18322 6410
rect 18334 6358 18386 6410
rect 7846 5814 7898 5866
rect 7910 5814 7962 5866
rect 7974 5814 8026 5866
rect 8038 5814 8090 5866
rect 14710 5814 14762 5866
rect 14774 5814 14826 5866
rect 14838 5814 14890 5866
rect 14902 5814 14954 5866
rect 12992 5712 13044 5764
rect 20536 5619 20588 5628
rect 20536 5585 20545 5619
rect 20545 5585 20579 5619
rect 20579 5585 20588 5619
rect 20536 5576 20588 5585
rect 4414 5270 4466 5322
rect 4478 5270 4530 5322
rect 4542 5270 4594 5322
rect 4606 5270 4658 5322
rect 11278 5270 11330 5322
rect 11342 5270 11394 5322
rect 11406 5270 11458 5322
rect 11470 5270 11522 5322
rect 18142 5270 18194 5322
rect 18206 5270 18258 5322
rect 18270 5270 18322 5322
rect 18334 5270 18386 5322
rect 16488 5168 16540 5220
rect 17960 5168 18012 5220
rect 7846 4726 7898 4778
rect 7910 4726 7962 4778
rect 7974 4726 8026 4778
rect 8038 4726 8090 4778
rect 14710 4726 14762 4778
rect 14774 4726 14826 4778
rect 14838 4726 14890 4778
rect 14902 4726 14954 4778
rect 21088 4624 21140 4676
rect 20536 4531 20588 4540
rect 20536 4497 20545 4531
rect 20545 4497 20579 4531
rect 20579 4497 20588 4531
rect 20536 4488 20588 4497
rect 4414 4182 4466 4234
rect 4478 4182 4530 4234
rect 4542 4182 4594 4234
rect 4606 4182 4658 4234
rect 11278 4182 11330 4234
rect 11342 4182 11394 4234
rect 11406 4182 11458 4234
rect 11470 4182 11522 4234
rect 18142 4182 18194 4234
rect 18206 4182 18258 4234
rect 18270 4182 18322 4234
rect 18334 4182 18386 4234
rect 14280 3944 14332 3996
rect 18512 3944 18564 3996
rect 7846 3638 7898 3690
rect 7910 3638 7962 3690
rect 7974 3638 8026 3690
rect 8038 3638 8090 3690
rect 14710 3638 14762 3690
rect 14774 3638 14826 3690
rect 14838 3638 14890 3690
rect 14902 3638 14954 3690
rect 4414 3094 4466 3146
rect 4478 3094 4530 3146
rect 4542 3094 4594 3146
rect 4606 3094 4658 3146
rect 11278 3094 11330 3146
rect 11342 3094 11394 3146
rect 11406 3094 11458 3146
rect 11470 3094 11522 3146
rect 18142 3094 18194 3146
rect 18206 3094 18258 3146
rect 18270 3094 18322 3146
rect 18334 3094 18386 3146
rect 7846 2550 7898 2602
rect 7910 2550 7962 2602
rect 7974 2550 8026 2602
rect 8038 2550 8090 2602
rect 14710 2550 14762 2602
rect 14774 2550 14826 2602
rect 14838 2550 14890 2602
rect 14902 2550 14954 2602
rect 14464 2448 14516 2500
rect 18604 2448 18656 2500
rect 4414 2006 4466 2058
rect 4478 2006 4530 2058
rect 4542 2006 4594 2058
rect 4606 2006 4658 2058
rect 11278 2006 11330 2058
rect 11342 2006 11394 2058
rect 11406 2006 11458 2058
rect 11470 2006 11522 2058
rect 18142 2006 18194 2058
rect 18206 2006 18258 2058
rect 18270 2006 18322 2058
rect 18334 2006 18386 2058
rect 17040 1156 17092 1208
rect 19064 1156 19116 1208
<< metal2 >>
rect 294 22176 350 22656
rect 846 22176 902 22656
rect 1398 22176 1454 22656
rect 1950 22176 2006 22656
rect 2502 22176 2558 22656
rect 3054 22176 3110 22656
rect 3606 22176 3662 22656
rect 4158 22176 4214 22656
rect 4710 22176 4766 22656
rect 5262 22176 5318 22656
rect 5814 22176 5870 22656
rect 6366 22176 6422 22656
rect 6918 22176 6974 22656
rect 7470 22176 7526 22656
rect 8022 22176 8078 22656
rect 8574 22176 8630 22656
rect 9126 22176 9182 22656
rect 9678 22176 9734 22656
rect 10230 22176 10286 22656
rect 10782 22176 10838 22656
rect 11334 22176 11390 22656
rect 11978 22176 12034 22656
rect 12530 22176 12586 22656
rect 13082 22176 13138 22656
rect 13634 22176 13690 22656
rect 14186 22176 14242 22656
rect 14738 22176 14794 22656
rect 15290 22176 15346 22656
rect 15842 22176 15898 22656
rect 16394 22176 16450 22656
rect 16946 22176 17002 22656
rect 17498 22176 17554 22656
rect 18050 22176 18106 22656
rect 18602 22176 18658 22656
rect 18878 22392 18934 22401
rect 18878 22327 18934 22336
rect 308 18486 336 22176
rect 296 18480 348 18486
rect 296 18422 348 18428
rect 860 13046 888 22176
rect 1412 22106 1440 22176
rect 1412 22078 1624 22106
rect 1596 13810 1624 22078
rect 1964 19098 1992 22176
rect 2412 19160 2464 19166
rect 2412 19102 2464 19108
rect 1952 19092 2004 19098
rect 1952 19034 2004 19040
rect 2424 18690 2452 19102
rect 2516 18826 2544 22176
rect 2504 18820 2556 18826
rect 2504 18762 2556 18768
rect 2872 18752 2924 18758
rect 2872 18694 2924 18700
rect 2412 18684 2464 18690
rect 2412 18626 2464 18632
rect 2424 17670 2452 18626
rect 2884 17738 2912 18694
rect 3068 17942 3096 22176
rect 3620 18486 3648 22176
rect 3516 18480 3568 18486
rect 3516 18422 3568 18428
rect 3608 18480 3660 18486
rect 3608 18422 3660 18428
rect 3528 18146 3556 18422
rect 3516 18140 3568 18146
rect 3516 18082 3568 18088
rect 3056 17936 3108 17942
rect 3056 17878 3108 17884
rect 2872 17732 2924 17738
rect 2872 17674 2924 17680
rect 4068 17732 4120 17738
rect 4068 17674 4120 17680
rect 1676 17664 1728 17670
rect 1676 17606 1728 17612
rect 2412 17664 2464 17670
rect 2412 17606 2464 17612
rect 1688 15970 1716 17606
rect 2884 17058 2912 17674
rect 3148 17596 3200 17602
rect 3148 17538 3200 17544
rect 3160 17126 3188 17538
rect 3332 17528 3384 17534
rect 3332 17470 3384 17476
rect 3148 17120 3200 17126
rect 3148 17062 3200 17068
rect 2872 17052 2924 17058
rect 2872 16994 2924 17000
rect 2964 16848 3016 16854
rect 2964 16790 3016 16796
rect 2976 16514 3004 16790
rect 2964 16508 3016 16514
rect 2964 16450 3016 16456
rect 3160 16106 3188 17062
rect 3344 16990 3372 17470
rect 4080 17097 4108 17674
rect 4066 17088 4122 17097
rect 4172 17058 4200 22176
rect 4724 19914 4752 22176
rect 4712 19908 4764 19914
rect 4712 19850 4764 19856
rect 5172 19704 5224 19710
rect 5172 19646 5224 19652
rect 5276 19658 5304 22176
rect 4388 19468 4684 19488
rect 4444 19466 4468 19468
rect 4524 19466 4548 19468
rect 4604 19466 4628 19468
rect 4466 19414 4468 19466
rect 4530 19414 4542 19466
rect 4604 19414 4606 19466
rect 4444 19412 4468 19414
rect 4524 19412 4548 19414
rect 4604 19412 4628 19414
rect 4388 19392 4684 19412
rect 5184 19166 5212 19646
rect 5276 19630 5396 19658
rect 5264 19568 5316 19574
rect 5264 19510 5316 19516
rect 4344 19160 4396 19166
rect 4344 19102 4396 19108
rect 5172 19160 5224 19166
rect 5172 19102 5224 19108
rect 4356 18826 4384 19102
rect 5276 18826 5304 19510
rect 5368 19114 5396 19630
rect 5368 19086 5672 19114
rect 5828 19098 5856 22176
rect 6380 19250 6408 22176
rect 6380 19222 6868 19250
rect 6552 19160 6604 19166
rect 6552 19102 6604 19108
rect 5448 19024 5500 19030
rect 5448 18966 5500 18972
rect 4344 18820 4396 18826
rect 4344 18762 4396 18768
rect 5264 18820 5316 18826
rect 5264 18762 5316 18768
rect 5460 18622 5488 18966
rect 5448 18616 5500 18622
rect 5448 18558 5500 18564
rect 4252 18480 4304 18486
rect 4252 18422 4304 18428
rect 5264 18480 5316 18486
rect 5264 18422 5316 18428
rect 4066 17023 4122 17032
rect 4160 17052 4212 17058
rect 4160 16994 4212 17000
rect 3332 16984 3384 16990
rect 3332 16926 3384 16932
rect 4160 16440 4212 16446
rect 4160 16382 4212 16388
rect 4172 16106 4200 16382
rect 3148 16100 3200 16106
rect 3148 16042 3200 16048
rect 4160 16100 4212 16106
rect 4160 16042 4212 16048
rect 1676 15964 1728 15970
rect 1676 15906 1728 15912
rect 1688 15426 1716 15906
rect 3884 15896 3936 15902
rect 3884 15838 3936 15844
rect 2964 15828 3016 15834
rect 2964 15770 3016 15776
rect 2976 15562 3004 15770
rect 2964 15556 3016 15562
rect 2964 15498 3016 15504
rect 1676 15420 1728 15426
rect 1676 15362 1728 15368
rect 3896 15358 3924 15838
rect 3700 15352 3752 15358
rect 3700 15294 3752 15300
rect 3884 15352 3936 15358
rect 3884 15294 3936 15300
rect 3608 15216 3660 15222
rect 3608 15158 3660 15164
rect 3620 14882 3648 15158
rect 3712 15018 3740 15294
rect 3700 15012 3752 15018
rect 3700 14954 3752 14960
rect 3608 14876 3660 14882
rect 3608 14818 3660 14824
rect 2504 13924 2556 13930
rect 2504 13866 2556 13872
rect 1596 13782 1716 13810
rect 848 13040 900 13046
rect 848 12982 900 12988
rect 1688 10666 1716 13782
rect 2516 13658 2544 13866
rect 3620 13862 3648 14818
rect 3896 14338 3924 15294
rect 4264 14814 4292 18422
rect 4388 18380 4684 18400
rect 4444 18378 4468 18380
rect 4524 18378 4548 18380
rect 4604 18378 4628 18380
rect 4466 18326 4468 18378
rect 4530 18326 4542 18378
rect 4604 18326 4606 18378
rect 4444 18324 4468 18326
rect 4524 18324 4548 18326
rect 4604 18324 4628 18326
rect 4388 18304 4684 18324
rect 5276 18078 5304 18422
rect 5264 18072 5316 18078
rect 5264 18014 5316 18020
rect 5460 17670 5488 18558
rect 5540 18004 5592 18010
rect 5540 17946 5592 17952
rect 5448 17664 5500 17670
rect 5448 17606 5500 17612
rect 5552 17602 5580 17946
rect 5540 17596 5592 17602
rect 5540 17538 5592 17544
rect 4388 17292 4684 17312
rect 4444 17290 4468 17292
rect 4524 17290 4548 17292
rect 4604 17290 4628 17292
rect 4466 17238 4468 17290
rect 4530 17238 4542 17290
rect 4604 17238 4606 17290
rect 4444 17236 4468 17238
rect 4524 17236 4548 17238
rect 4604 17236 4628 17238
rect 4388 17216 4684 17236
rect 5644 17058 5672 19086
rect 5816 19092 5868 19098
rect 5816 19034 5868 19040
rect 6564 18622 6592 19102
rect 6840 19030 6868 19222
rect 6736 19024 6788 19030
rect 6736 18966 6788 18972
rect 6828 19024 6880 19030
rect 6828 18966 6880 18972
rect 6552 18616 6604 18622
rect 6552 18558 6604 18564
rect 5908 17936 5960 17942
rect 5908 17878 5960 17884
rect 5724 17392 5776 17398
rect 5724 17334 5776 17340
rect 5632 17052 5684 17058
rect 5632 16994 5684 17000
rect 5736 16990 5764 17334
rect 5724 16984 5776 16990
rect 5724 16926 5776 16932
rect 4388 16204 4684 16224
rect 4444 16202 4468 16204
rect 4524 16202 4548 16204
rect 4604 16202 4628 16204
rect 4466 16150 4468 16202
rect 4530 16150 4542 16202
rect 4604 16150 4606 16202
rect 4444 16148 4468 16150
rect 4524 16148 4548 16150
rect 4604 16148 4628 16150
rect 4388 16128 4684 16148
rect 5736 15902 5764 16926
rect 5724 15896 5776 15902
rect 5724 15838 5776 15844
rect 5736 15222 5764 15838
rect 5724 15216 5776 15222
rect 5724 15158 5776 15164
rect 4388 15116 4684 15136
rect 4444 15114 4468 15116
rect 4524 15114 4548 15116
rect 4604 15114 4628 15116
rect 4466 15062 4468 15114
rect 4530 15062 4542 15114
rect 4604 15062 4606 15114
rect 4444 15060 4468 15062
rect 4524 15060 4548 15062
rect 4604 15060 4628 15062
rect 4388 15040 4684 15060
rect 4252 14808 4304 14814
rect 4252 14750 4304 14756
rect 3884 14332 3936 14338
rect 3884 14274 3936 14280
rect 5540 14128 5592 14134
rect 5540 14070 5592 14076
rect 4388 14028 4684 14048
rect 4444 14026 4468 14028
rect 4524 14026 4548 14028
rect 4604 14026 4628 14028
rect 4466 13974 4468 14026
rect 4530 13974 4542 14026
rect 4604 13974 4606 14026
rect 4444 13972 4468 13974
rect 4524 13972 4548 13974
rect 4604 13972 4628 13974
rect 4388 13952 4684 13972
rect 3608 13856 3660 13862
rect 3608 13798 3660 13804
rect 5552 13726 5580 14070
rect 5540 13720 5592 13726
rect 5540 13662 5592 13668
rect 2504 13652 2556 13658
rect 2504 13594 2556 13600
rect 5920 13318 5948 17878
rect 6564 16990 6592 18558
rect 6552 16984 6604 16990
rect 6552 16926 6604 16932
rect 6564 16582 6592 16926
rect 6552 16576 6604 16582
rect 6552 16518 6604 16524
rect 6184 15828 6236 15834
rect 6184 15770 6236 15776
rect 6196 15562 6224 15770
rect 6184 15556 6236 15562
rect 6184 15498 6236 15504
rect 6748 14354 6776 18966
rect 6932 18282 6960 22176
rect 7484 18486 7512 22176
rect 8036 20202 8064 22176
rect 7760 20174 8064 20202
rect 7656 18684 7708 18690
rect 7656 18626 7708 18632
rect 7472 18480 7524 18486
rect 7472 18422 7524 18428
rect 6920 18276 6972 18282
rect 6920 18218 6972 18224
rect 7668 18214 7696 18626
rect 7656 18208 7708 18214
rect 7656 18150 7708 18156
rect 6920 17460 6972 17466
rect 6920 17402 6972 17408
rect 6932 16650 6960 17402
rect 7668 17194 7696 18150
rect 7656 17188 7708 17194
rect 7656 17130 7708 17136
rect 7104 16916 7156 16922
rect 7104 16858 7156 16864
rect 6920 16644 6972 16650
rect 6920 16586 6972 16592
rect 7116 16378 7144 16858
rect 7380 16440 7432 16446
rect 7380 16382 7432 16388
rect 7104 16372 7156 16378
rect 7104 16314 7156 16320
rect 7116 16106 7144 16314
rect 7392 16106 7420 16382
rect 7104 16100 7156 16106
rect 7104 16042 7156 16048
rect 7380 16100 7432 16106
rect 7380 16042 7432 16048
rect 7760 15970 7788 20174
rect 7820 20012 8116 20032
rect 7876 20010 7900 20012
rect 7956 20010 7980 20012
rect 8036 20010 8060 20012
rect 7898 19958 7900 20010
rect 7962 19958 7974 20010
rect 8036 19958 8038 20010
rect 7876 19956 7900 19958
rect 7956 19956 7980 19958
rect 8036 19956 8060 19958
rect 7820 19936 8116 19956
rect 8208 19092 8260 19098
rect 8208 19034 8260 19040
rect 7820 18924 8116 18944
rect 7876 18922 7900 18924
rect 7956 18922 7980 18924
rect 8036 18922 8060 18924
rect 7898 18870 7900 18922
rect 7962 18870 7974 18922
rect 8036 18870 8038 18922
rect 7876 18868 7900 18870
rect 7956 18868 7980 18870
rect 8036 18868 8060 18870
rect 7820 18848 8116 18868
rect 8220 18826 8248 19034
rect 8208 18820 8260 18826
rect 8208 18762 8260 18768
rect 7932 18616 7984 18622
rect 7932 18558 7984 18564
rect 7840 18548 7892 18554
rect 7840 18490 7892 18496
rect 7852 18146 7880 18490
rect 7840 18140 7892 18146
rect 7840 18082 7892 18088
rect 7944 18078 7972 18558
rect 8220 18146 8248 18762
rect 8484 18480 8536 18486
rect 8484 18422 8536 18428
rect 8208 18140 8260 18146
rect 8208 18082 8260 18088
rect 7932 18072 7984 18078
rect 7932 18014 7984 18020
rect 8392 18072 8444 18078
rect 8392 18014 8444 18020
rect 7820 17836 8116 17856
rect 7876 17834 7900 17836
rect 7956 17834 7980 17836
rect 8036 17834 8060 17836
rect 7898 17782 7900 17834
rect 7962 17782 7974 17834
rect 8036 17782 8038 17834
rect 7876 17780 7900 17782
rect 7956 17780 7980 17782
rect 8036 17780 8060 17782
rect 7820 17760 8116 17780
rect 8404 16854 8432 18014
rect 8392 16848 8444 16854
rect 8392 16790 8444 16796
rect 7820 16748 8116 16768
rect 7876 16746 7900 16748
rect 7956 16746 7980 16748
rect 8036 16746 8060 16748
rect 7898 16694 7900 16746
rect 7962 16694 7974 16746
rect 8036 16694 8038 16746
rect 7876 16692 7900 16694
rect 7956 16692 7980 16694
rect 8036 16692 8060 16694
rect 7820 16672 8116 16692
rect 7748 15964 7800 15970
rect 7748 15906 7800 15912
rect 7748 15760 7800 15766
rect 7748 15702 7800 15708
rect 6828 15420 6880 15426
rect 6828 15362 6880 15368
rect 6840 14474 6868 15362
rect 7760 14814 7788 15702
rect 7820 15660 8116 15680
rect 7876 15658 7900 15660
rect 7956 15658 7980 15660
rect 8036 15658 8060 15660
rect 7898 15606 7900 15658
rect 7962 15606 7974 15658
rect 8036 15606 8038 15658
rect 7876 15604 7900 15606
rect 7956 15604 7980 15606
rect 8036 15604 8060 15606
rect 7820 15584 8116 15604
rect 8208 15420 8260 15426
rect 8208 15362 8260 15368
rect 7748 14808 7800 14814
rect 7748 14750 7800 14756
rect 7820 14572 8116 14592
rect 7876 14570 7900 14572
rect 7956 14570 7980 14572
rect 8036 14570 8060 14572
rect 7898 14518 7900 14570
rect 7962 14518 7974 14570
rect 8036 14518 8038 14570
rect 7876 14516 7900 14518
rect 7956 14516 7980 14518
rect 8036 14516 8060 14518
rect 7820 14496 8116 14516
rect 6828 14468 6880 14474
rect 6828 14410 6880 14416
rect 6092 14332 6144 14338
rect 6748 14326 6868 14354
rect 6092 14274 6144 14280
rect 6104 13794 6132 14274
rect 6184 14264 6236 14270
rect 6184 14206 6236 14212
rect 6276 14264 6328 14270
rect 6276 14206 6328 14212
rect 6092 13788 6144 13794
rect 6092 13730 6144 13736
rect 6196 13386 6224 14206
rect 6288 13930 6316 14206
rect 6276 13924 6328 13930
rect 6276 13866 6328 13872
rect 6276 13720 6328 13726
rect 6276 13662 6328 13668
rect 6184 13380 6236 13386
rect 6184 13322 6236 13328
rect 5908 13312 5960 13318
rect 5908 13254 5960 13260
rect 6288 13182 6316 13662
rect 6276 13176 6328 13182
rect 6276 13118 6328 13124
rect 4388 12940 4684 12960
rect 4444 12938 4468 12940
rect 4524 12938 4548 12940
rect 4604 12938 4628 12940
rect 4466 12886 4468 12938
rect 4530 12886 4542 12938
rect 4604 12886 4606 12938
rect 4444 12884 4468 12886
rect 4524 12884 4548 12886
rect 4604 12884 4628 12886
rect 4388 12864 4684 12884
rect 4388 11852 4684 11872
rect 4444 11850 4468 11852
rect 4524 11850 4548 11852
rect 4604 11850 4628 11852
rect 4466 11798 4468 11850
rect 4530 11798 4542 11850
rect 4604 11798 4606 11850
rect 4444 11796 4468 11798
rect 4524 11796 4548 11798
rect 4604 11796 4628 11798
rect 4388 11776 4684 11796
rect 6840 11618 6868 14326
rect 7380 14264 7432 14270
rect 7380 14206 7432 14212
rect 7392 13726 7420 14206
rect 8220 13930 8248 15362
rect 8404 14762 8432 16790
rect 8496 14882 8524 18422
rect 8588 18146 8616 22176
rect 9036 19024 9088 19030
rect 9036 18966 9088 18972
rect 8852 18684 8904 18690
rect 8852 18626 8904 18632
rect 8576 18140 8628 18146
rect 8576 18082 8628 18088
rect 8864 17942 8892 18626
rect 8852 17936 8904 17942
rect 8852 17878 8904 17884
rect 8944 16848 8996 16854
rect 8944 16790 8996 16796
rect 8484 14876 8536 14882
rect 8484 14818 8536 14824
rect 8668 14876 8720 14882
rect 8668 14818 8720 14824
rect 8404 14734 8524 14762
rect 8392 14672 8444 14678
rect 8392 14614 8444 14620
rect 8208 13924 8260 13930
rect 8208 13866 8260 13872
rect 7380 13720 7432 13726
rect 7380 13662 7432 13668
rect 7392 12842 7420 13662
rect 7820 13484 8116 13504
rect 7876 13482 7900 13484
rect 7956 13482 7980 13484
rect 8036 13482 8060 13484
rect 7898 13430 7900 13482
rect 7962 13430 7974 13482
rect 8036 13430 8038 13482
rect 7876 13428 7900 13430
rect 7956 13428 7980 13430
rect 8036 13428 8060 13430
rect 7820 13408 8116 13428
rect 7380 12836 7432 12842
rect 7380 12778 7432 12784
rect 7564 12836 7616 12842
rect 7564 12778 7616 12784
rect 7576 12706 7604 12778
rect 7564 12700 7616 12706
rect 7564 12642 7616 12648
rect 7576 12230 7604 12642
rect 8220 12638 8248 13866
rect 8404 13250 8432 14614
rect 8496 13250 8524 14734
rect 8680 14338 8708 14818
rect 8668 14332 8720 14338
rect 8668 14274 8720 14280
rect 8680 13930 8708 14274
rect 8668 13924 8720 13930
rect 8668 13866 8720 13872
rect 8392 13244 8444 13250
rect 8392 13186 8444 13192
rect 8484 13244 8536 13250
rect 8484 13186 8536 13192
rect 8404 12842 8432 13186
rect 8392 12836 8444 12842
rect 8392 12778 8444 12784
rect 8208 12632 8260 12638
rect 8208 12574 8260 12580
rect 7820 12396 8116 12416
rect 7876 12394 7900 12396
rect 7956 12394 7980 12396
rect 8036 12394 8060 12396
rect 7898 12342 7900 12394
rect 7962 12342 7974 12394
rect 8036 12342 8038 12394
rect 7876 12340 7900 12342
rect 7956 12340 7980 12342
rect 8036 12340 8060 12342
rect 7820 12320 8116 12340
rect 7196 12224 7248 12230
rect 7196 12166 7248 12172
rect 7564 12224 7616 12230
rect 7564 12166 7616 12172
rect 6828 11612 6880 11618
rect 6828 11554 6880 11560
rect 4388 10764 4684 10784
rect 4444 10762 4468 10764
rect 4524 10762 4548 10764
rect 4604 10762 4628 10764
rect 4466 10710 4468 10762
rect 4530 10710 4542 10762
rect 4604 10710 4606 10762
rect 4444 10708 4468 10710
rect 4524 10708 4548 10710
rect 4604 10708 4628 10710
rect 4388 10688 4684 10708
rect 1676 10660 1728 10666
rect 1676 10602 1728 10608
rect 7208 10462 7236 12166
rect 7288 12156 7340 12162
rect 7288 12098 7340 12104
rect 7300 11618 7328 12098
rect 7288 11612 7340 11618
rect 7288 11554 7340 11560
rect 8404 11550 8432 12778
rect 8392 11544 8444 11550
rect 8392 11486 8444 11492
rect 8300 11408 8352 11414
rect 8300 11350 8352 11356
rect 7820 11308 8116 11328
rect 7876 11306 7900 11308
rect 7956 11306 7980 11308
rect 8036 11306 8060 11308
rect 7898 11254 7900 11306
rect 7962 11254 7974 11306
rect 8036 11254 8038 11306
rect 7876 11252 7900 11254
rect 7956 11252 7980 11254
rect 8036 11252 8060 11254
rect 7820 11232 8116 11252
rect 8312 11210 8340 11350
rect 8496 11210 8524 13186
rect 8956 12298 8984 16790
rect 9048 15834 9076 18966
rect 9140 18826 9168 22176
rect 9588 19772 9640 19778
rect 9588 19714 9640 19720
rect 9496 19024 9548 19030
rect 9496 18966 9548 18972
rect 9128 18820 9180 18826
rect 9128 18762 9180 18768
rect 9508 18622 9536 18966
rect 9600 18690 9628 19714
rect 9692 19250 9720 22176
rect 9692 19222 9904 19250
rect 9772 19092 9824 19098
rect 9772 19034 9824 19040
rect 9588 18684 9640 18690
rect 9588 18626 9640 18632
rect 9784 18672 9812 19034
rect 9876 18826 9904 19222
rect 10244 19098 10272 22176
rect 9956 19092 10008 19098
rect 9956 19034 10008 19040
rect 10232 19092 10284 19098
rect 10232 19034 10284 19040
rect 9864 18820 9916 18826
rect 9864 18762 9916 18768
rect 9864 18684 9916 18690
rect 9784 18644 9864 18672
rect 9496 18616 9548 18622
rect 9496 18558 9548 18564
rect 9600 18078 9628 18626
rect 9588 18072 9640 18078
rect 9588 18014 9640 18020
rect 9128 17392 9180 17398
rect 9128 17334 9180 17340
rect 9140 17058 9168 17334
rect 9128 17052 9180 17058
rect 9128 16994 9180 17000
rect 9140 16582 9168 16994
rect 9128 16576 9180 16582
rect 9128 16518 9180 16524
rect 9784 16514 9812 18644
rect 9864 18626 9916 18632
rect 9968 18622 9996 19034
rect 9956 18616 10008 18622
rect 9956 18558 10008 18564
rect 10600 18548 10652 18554
rect 10600 18490 10652 18496
rect 10416 17052 10468 17058
rect 10416 16994 10468 17000
rect 10140 16848 10192 16854
rect 10140 16790 10192 16796
rect 9772 16508 9824 16514
rect 9772 16450 9824 16456
rect 10152 15970 10180 16790
rect 10428 16582 10456 16994
rect 10416 16576 10468 16582
rect 10416 16518 10468 16524
rect 10140 15964 10192 15970
rect 10140 15906 10192 15912
rect 9036 15828 9088 15834
rect 9036 15770 9088 15776
rect 10048 15216 10100 15222
rect 10048 15158 10100 15164
rect 9956 14196 10008 14202
rect 9956 14138 10008 14144
rect 9968 13862 9996 14138
rect 9956 13856 10008 13862
rect 9956 13798 10008 13804
rect 10060 13318 10088 15158
rect 10232 14876 10284 14882
rect 10232 14818 10284 14824
rect 10244 14474 10272 14818
rect 10232 14468 10284 14474
rect 10232 14410 10284 14416
rect 10048 13312 10100 13318
rect 10048 13254 10100 13260
rect 10232 12564 10284 12570
rect 10232 12506 10284 12512
rect 8944 12292 8996 12298
rect 8944 12234 8996 12240
rect 8668 11952 8720 11958
rect 8668 11894 8720 11900
rect 8680 11618 8708 11894
rect 8668 11612 8720 11618
rect 8668 11554 8720 11560
rect 8576 11544 8628 11550
rect 8576 11486 8628 11492
rect 8300 11204 8352 11210
rect 8300 11146 8352 11152
rect 8484 11204 8536 11210
rect 8484 11146 8536 11152
rect 8588 11006 8616 11486
rect 8956 11142 8984 12234
rect 9772 12088 9824 12094
rect 9772 12030 9824 12036
rect 9784 11754 9812 12030
rect 10244 12026 10272 12506
rect 10416 12156 10468 12162
rect 10416 12098 10468 12104
rect 10232 12020 10284 12026
rect 10232 11962 10284 11968
rect 10428 11754 10456 12098
rect 9772 11748 9824 11754
rect 9772 11690 9824 11696
rect 10416 11748 10468 11754
rect 10416 11690 10468 11696
rect 8944 11136 8996 11142
rect 8944 11078 8996 11084
rect 10048 11068 10100 11074
rect 10048 11010 10100 11016
rect 8576 11000 8628 11006
rect 8576 10942 8628 10948
rect 8588 10598 8616 10942
rect 8576 10592 8628 10598
rect 8576 10534 8628 10540
rect 7196 10456 7248 10462
rect 7196 10398 7248 10404
rect 4388 9676 4684 9696
rect 4444 9674 4468 9676
rect 4524 9674 4548 9676
rect 4604 9674 4628 9676
rect 4466 9622 4468 9674
rect 4530 9622 4542 9674
rect 4604 9622 4606 9674
rect 4444 9620 4468 9622
rect 4524 9620 4548 9622
rect 4604 9620 4628 9622
rect 4388 9600 4684 9620
rect 7208 9374 7236 10398
rect 9312 10388 9364 10394
rect 9312 10330 9364 10336
rect 7820 10220 8116 10240
rect 7876 10218 7900 10220
rect 7956 10218 7980 10220
rect 8036 10218 8060 10220
rect 7898 10166 7900 10218
rect 7962 10166 7974 10218
rect 8036 10166 8038 10218
rect 7876 10164 7900 10166
rect 7956 10164 7980 10166
rect 8036 10164 8060 10166
rect 7820 10144 8116 10164
rect 9324 9850 9352 10330
rect 10060 10122 10088 11010
rect 10048 10116 10100 10122
rect 10048 10058 10100 10064
rect 10508 9912 10560 9918
rect 10508 9854 10560 9860
rect 9312 9844 9364 9850
rect 9312 9786 9364 9792
rect 9324 9510 9352 9786
rect 10520 9578 10548 9854
rect 10508 9572 10560 9578
rect 10508 9514 10560 9520
rect 9312 9504 9364 9510
rect 9312 9446 9364 9452
rect 7196 9368 7248 9374
rect 7196 9310 7248 9316
rect 8208 9232 8260 9238
rect 8208 9174 8260 9180
rect 7820 9132 8116 9152
rect 7876 9130 7900 9132
rect 7956 9130 7980 9132
rect 8036 9130 8060 9132
rect 7898 9078 7900 9130
rect 7962 9078 7974 9130
rect 8036 9078 8038 9130
rect 7876 9076 7900 9078
rect 7956 9076 7980 9078
rect 8036 9076 8060 9078
rect 7820 9056 8116 9076
rect 8220 8830 8248 9174
rect 8208 8824 8260 8830
rect 8208 8766 8260 8772
rect 4388 8588 4684 8608
rect 4444 8586 4468 8588
rect 4524 8586 4548 8588
rect 4604 8586 4628 8588
rect 4466 8534 4468 8586
rect 4530 8534 4542 8586
rect 4604 8534 4606 8586
rect 4444 8532 4468 8534
rect 4524 8532 4548 8534
rect 4604 8532 4628 8534
rect 4388 8512 4684 8532
rect 7820 8044 8116 8064
rect 7876 8042 7900 8044
rect 7956 8042 7980 8044
rect 8036 8042 8060 8044
rect 7898 7990 7900 8042
rect 7962 7990 7974 8042
rect 8036 7990 8038 8042
rect 7876 7988 7900 7990
rect 7956 7988 7980 7990
rect 8036 7988 8060 7990
rect 7820 7968 8116 7988
rect 4388 7500 4684 7520
rect 4444 7498 4468 7500
rect 4524 7498 4548 7500
rect 4604 7498 4628 7500
rect 4466 7446 4468 7498
rect 4530 7446 4542 7498
rect 4604 7446 4606 7498
rect 4444 7444 4468 7446
rect 4524 7444 4548 7446
rect 4604 7444 4628 7446
rect 4388 7424 4684 7444
rect 8220 7198 8248 8766
rect 7380 7192 7432 7198
rect 7380 7134 7432 7140
rect 8208 7192 8260 7198
rect 8208 7134 8260 7140
rect 4068 6716 4120 6722
rect 4068 6658 4120 6664
rect 4080 5673 4108 6658
rect 7392 6654 7420 7134
rect 9864 7124 9916 7130
rect 9864 7066 9916 7072
rect 7820 6956 8116 6976
rect 7876 6954 7900 6956
rect 7956 6954 7980 6956
rect 8036 6954 8060 6956
rect 7898 6902 7900 6954
rect 7962 6902 7974 6954
rect 8036 6902 8038 6954
rect 7876 6900 7900 6902
rect 7956 6900 7980 6902
rect 8036 6900 8060 6902
rect 7820 6880 8116 6900
rect 7380 6648 7432 6654
rect 7380 6590 7432 6596
rect 9876 6586 9904 7066
rect 10612 6722 10640 18490
rect 10796 17534 10824 22176
rect 11348 19658 11376 22176
rect 11348 19630 11652 19658
rect 11252 19468 11548 19488
rect 11308 19466 11332 19468
rect 11388 19466 11412 19468
rect 11468 19466 11492 19468
rect 11330 19414 11332 19466
rect 11394 19414 11406 19466
rect 11468 19414 11470 19466
rect 11308 19412 11332 19414
rect 11388 19412 11412 19414
rect 11468 19412 11492 19414
rect 11252 19392 11548 19412
rect 11060 19364 11112 19370
rect 11060 19306 11112 19312
rect 10968 19024 11020 19030
rect 10968 18966 11020 18972
rect 10784 17528 10836 17534
rect 10784 17470 10836 17476
rect 10980 16990 11008 18966
rect 11072 18758 11100 19306
rect 11152 19024 11204 19030
rect 11152 18966 11204 18972
rect 11060 18752 11112 18758
rect 11060 18694 11112 18700
rect 11164 18282 11192 18966
rect 11252 18380 11548 18400
rect 11308 18378 11332 18380
rect 11388 18378 11412 18380
rect 11468 18378 11492 18380
rect 11330 18326 11332 18378
rect 11394 18326 11406 18378
rect 11468 18326 11470 18378
rect 11308 18324 11332 18326
rect 11388 18324 11412 18326
rect 11468 18324 11492 18326
rect 11252 18304 11548 18324
rect 11152 18276 11204 18282
rect 11152 18218 11204 18224
rect 11252 17292 11548 17312
rect 11308 17290 11332 17292
rect 11388 17290 11412 17292
rect 11468 17290 11492 17292
rect 11330 17238 11332 17290
rect 11394 17238 11406 17290
rect 11468 17238 11470 17290
rect 11308 17236 11332 17238
rect 11388 17236 11412 17238
rect 11468 17236 11492 17238
rect 11252 17216 11548 17236
rect 10968 16984 11020 16990
rect 10968 16926 11020 16932
rect 11252 16204 11548 16224
rect 11308 16202 11332 16204
rect 11388 16202 11412 16204
rect 11468 16202 11492 16204
rect 11330 16150 11332 16202
rect 11394 16150 11406 16202
rect 11468 16150 11470 16202
rect 11308 16148 11332 16150
rect 11388 16148 11412 16150
rect 11468 16148 11492 16150
rect 11252 16128 11548 16148
rect 11060 15896 11112 15902
rect 10980 15844 11060 15850
rect 10980 15838 11112 15844
rect 10980 15822 11100 15838
rect 10980 14950 11008 15822
rect 11252 15116 11548 15136
rect 11308 15114 11332 15116
rect 11388 15114 11412 15116
rect 11468 15114 11492 15116
rect 11330 15062 11332 15114
rect 11394 15062 11406 15114
rect 11468 15062 11470 15114
rect 11308 15060 11332 15062
rect 11388 15060 11412 15062
rect 11468 15060 11492 15062
rect 11252 15040 11548 15060
rect 10968 14944 11020 14950
rect 10968 14886 11020 14892
rect 10980 13726 11008 14886
rect 11252 14028 11548 14048
rect 11308 14026 11332 14028
rect 11388 14026 11412 14028
rect 11468 14026 11492 14028
rect 11330 13974 11332 14026
rect 11394 13974 11406 14026
rect 11468 13974 11470 14026
rect 11308 13972 11332 13974
rect 11388 13972 11412 13974
rect 11468 13972 11492 13974
rect 11252 13952 11548 13972
rect 10876 13720 10928 13726
rect 10876 13662 10928 13668
rect 10968 13720 11020 13726
rect 10968 13662 11020 13668
rect 10888 13386 10916 13662
rect 11152 13652 11204 13658
rect 11152 13594 11204 13600
rect 10876 13380 10928 13386
rect 10876 13322 10928 13328
rect 11164 12842 11192 13594
rect 11252 12940 11548 12960
rect 11308 12938 11332 12940
rect 11388 12938 11412 12940
rect 11468 12938 11492 12940
rect 11330 12886 11332 12938
rect 11394 12886 11406 12938
rect 11468 12886 11470 12938
rect 11308 12884 11332 12886
rect 11388 12884 11412 12886
rect 11468 12884 11492 12886
rect 11252 12864 11548 12884
rect 11152 12836 11204 12842
rect 11152 12778 11204 12784
rect 11428 12632 11480 12638
rect 11428 12574 11480 12580
rect 11440 12298 11468 12574
rect 11428 12292 11480 12298
rect 11428 12234 11480 12240
rect 11252 11852 11548 11872
rect 11308 11850 11332 11852
rect 11388 11850 11412 11852
rect 11468 11850 11492 11852
rect 11330 11798 11332 11850
rect 11394 11798 11406 11850
rect 11468 11798 11470 11850
rect 11308 11796 11332 11798
rect 11388 11796 11412 11798
rect 11468 11796 11492 11798
rect 11252 11776 11548 11796
rect 11624 11482 11652 19630
rect 11704 19024 11756 19030
rect 11704 18966 11756 18972
rect 11796 19024 11848 19030
rect 11796 18966 11848 18972
rect 11716 18146 11744 18966
rect 11808 18486 11836 18966
rect 11796 18480 11848 18486
rect 11796 18422 11848 18428
rect 11704 18140 11756 18146
rect 11704 18082 11756 18088
rect 11888 18072 11940 18078
rect 11888 18014 11940 18020
rect 11704 17936 11756 17942
rect 11704 17878 11756 17884
rect 11716 14882 11744 17878
rect 11796 16644 11848 16650
rect 11796 16586 11848 16592
rect 11808 15902 11836 16586
rect 11796 15896 11848 15902
rect 11796 15838 11848 15844
rect 11900 15306 11928 18014
rect 11808 15278 11928 15306
rect 11704 14876 11756 14882
rect 11704 14818 11756 14824
rect 11704 14128 11756 14134
rect 11704 14070 11756 14076
rect 11716 13726 11744 14070
rect 11704 13720 11756 13726
rect 11704 13662 11756 13668
rect 11704 13176 11756 13182
rect 11704 13118 11756 13124
rect 11716 12706 11744 13118
rect 11704 12700 11756 12706
rect 11704 12642 11756 12648
rect 11808 11906 11836 15278
rect 11992 15170 12020 22176
rect 12440 18480 12492 18486
rect 12440 18422 12492 18428
rect 12452 18078 12480 18422
rect 12440 18072 12492 18078
rect 12440 18014 12492 18020
rect 12544 17942 12572 22176
rect 12624 19092 12676 19098
rect 12624 19034 12676 19040
rect 12636 18554 12664 19034
rect 12716 19024 12768 19030
rect 12716 18966 12768 18972
rect 12624 18548 12676 18554
rect 12624 18490 12676 18496
rect 12532 17936 12584 17942
rect 12532 17878 12584 17884
rect 12348 17732 12400 17738
rect 12348 17674 12400 17680
rect 12360 17398 12388 17674
rect 12348 17392 12400 17398
rect 12348 17334 12400 17340
rect 12348 17052 12400 17058
rect 12348 16994 12400 17000
rect 12360 16650 12388 16994
rect 12348 16644 12400 16650
rect 12348 16586 12400 16592
rect 12728 16446 12756 18966
rect 12808 18684 12860 18690
rect 12808 18626 12860 18632
rect 12820 16990 12848 18626
rect 12992 17936 13044 17942
rect 12992 17878 13044 17884
rect 12900 17052 12952 17058
rect 12900 16994 12952 17000
rect 12808 16984 12860 16990
rect 12808 16926 12860 16932
rect 12808 16848 12860 16854
rect 12808 16790 12860 16796
rect 12820 16650 12848 16790
rect 12808 16644 12860 16650
rect 12808 16586 12860 16592
rect 12912 16514 12940 16994
rect 12900 16508 12952 16514
rect 12900 16450 12952 16456
rect 12716 16440 12768 16446
rect 12716 16382 12768 16388
rect 11716 11878 11836 11906
rect 11900 15142 12020 15170
rect 11612 11476 11664 11482
rect 11612 11418 11664 11424
rect 11252 10764 11548 10784
rect 11308 10762 11332 10764
rect 11388 10762 11412 10764
rect 11468 10762 11492 10764
rect 11330 10710 11332 10762
rect 11394 10710 11406 10762
rect 11468 10710 11470 10762
rect 11308 10708 11332 10710
rect 11388 10708 11412 10710
rect 11468 10708 11492 10710
rect 11252 10688 11548 10708
rect 11716 10666 11744 11878
rect 11704 10660 11756 10666
rect 11704 10602 11756 10608
rect 11060 10320 11112 10326
rect 11060 10262 11112 10268
rect 11072 9306 11100 10262
rect 11612 10048 11664 10054
rect 11612 9990 11664 9996
rect 11152 9912 11204 9918
rect 11152 9854 11204 9860
rect 11164 9442 11192 9854
rect 11252 9676 11548 9696
rect 11308 9674 11332 9676
rect 11388 9674 11412 9676
rect 11468 9674 11492 9676
rect 11330 9622 11332 9674
rect 11394 9622 11406 9674
rect 11468 9622 11470 9674
rect 11308 9620 11332 9622
rect 11388 9620 11412 9622
rect 11468 9620 11492 9622
rect 11252 9600 11548 9620
rect 11624 9442 11652 9990
rect 11152 9436 11204 9442
rect 11152 9378 11204 9384
rect 11612 9436 11664 9442
rect 11612 9378 11664 9384
rect 11060 9300 11112 9306
rect 11060 9242 11112 9248
rect 10876 9232 10928 9238
rect 10876 9174 10928 9180
rect 10888 9034 10916 9174
rect 10876 9028 10928 9034
rect 10876 8970 10928 8976
rect 11164 8762 11192 9378
rect 11716 8966 11744 10602
rect 11796 10524 11848 10530
rect 11796 10466 11848 10472
rect 11808 9442 11836 10466
rect 11796 9436 11848 9442
rect 11796 9378 11848 9384
rect 11704 8960 11756 8966
rect 11704 8902 11756 8908
rect 11808 8898 11836 9378
rect 11796 8892 11848 8898
rect 11796 8834 11848 8840
rect 11152 8756 11204 8762
rect 11152 8698 11204 8704
rect 11252 8588 11548 8608
rect 11308 8586 11332 8588
rect 11388 8586 11412 8588
rect 11468 8586 11492 8588
rect 11330 8534 11332 8586
rect 11394 8534 11406 8586
rect 11468 8534 11470 8586
rect 11308 8532 11332 8534
rect 11388 8532 11412 8534
rect 11468 8532 11492 8534
rect 11252 8512 11548 8532
rect 11900 8490 11928 15142
rect 12728 14950 12756 16382
rect 12912 16106 12940 16450
rect 12900 16100 12952 16106
rect 12900 16042 12952 16048
rect 12716 14944 12768 14950
rect 12716 14886 12768 14892
rect 12164 14808 12216 14814
rect 12164 14750 12216 14756
rect 12348 14808 12400 14814
rect 12348 14750 12400 14756
rect 11980 14672 12032 14678
rect 11980 14614 12032 14620
rect 12072 14672 12124 14678
rect 12072 14614 12124 14620
rect 11992 14474 12020 14614
rect 11980 14468 12032 14474
rect 11980 14410 12032 14416
rect 11980 13788 12032 13794
rect 11980 13730 12032 13736
rect 11992 13658 12020 13730
rect 11980 13652 12032 13658
rect 11980 13594 12032 13600
rect 12084 10938 12112 14614
rect 12072 10932 12124 10938
rect 12072 10874 12124 10880
rect 12084 10462 12112 10874
rect 12072 10456 12124 10462
rect 12072 10398 12124 10404
rect 12176 9510 12204 14750
rect 12256 14400 12308 14406
rect 12256 14342 12308 14348
rect 12268 13930 12296 14342
rect 12256 13924 12308 13930
rect 12256 13866 12308 13872
rect 12360 13794 12388 14750
rect 12624 14332 12676 14338
rect 12624 14274 12676 14280
rect 12636 13930 12664 14274
rect 12624 13924 12676 13930
rect 12624 13866 12676 13872
rect 12348 13788 12400 13794
rect 12348 13730 12400 13736
rect 12624 13108 12676 13114
rect 12624 13050 12676 13056
rect 12636 12638 12664 13050
rect 12624 12632 12676 12638
rect 12624 12574 12676 12580
rect 12440 12088 12492 12094
rect 12440 12030 12492 12036
rect 12452 11754 12480 12030
rect 12440 11748 12492 11754
rect 12440 11690 12492 11696
rect 12452 10530 12480 11690
rect 12440 10524 12492 10530
rect 12440 10466 12492 10472
rect 12716 10524 12768 10530
rect 12716 10466 12768 10472
rect 12348 9980 12400 9986
rect 12348 9922 12400 9928
rect 12360 9578 12388 9922
rect 12348 9572 12400 9578
rect 12348 9514 12400 9520
rect 12728 9510 12756 10466
rect 12164 9504 12216 9510
rect 12164 9446 12216 9452
rect 12716 9504 12768 9510
rect 12716 9446 12768 9452
rect 12176 9034 12204 9446
rect 12164 9028 12216 9034
rect 12164 8970 12216 8976
rect 11888 8484 11940 8490
rect 11888 8426 11940 8432
rect 11336 8280 11388 8286
rect 11336 8222 11388 8228
rect 10692 8144 10744 8150
rect 10692 8086 10744 8092
rect 10704 7946 10732 8086
rect 10692 7940 10744 7946
rect 10692 7882 10744 7888
rect 11348 7878 11376 8222
rect 11336 7872 11388 7878
rect 11336 7814 11388 7820
rect 10876 7736 10928 7742
rect 10876 7678 10928 7684
rect 11060 7736 11112 7742
rect 11060 7678 11112 7684
rect 10888 6858 10916 7678
rect 11072 7402 11100 7678
rect 11252 7500 11548 7520
rect 11308 7498 11332 7500
rect 11388 7498 11412 7500
rect 11468 7498 11492 7500
rect 11330 7446 11332 7498
rect 11394 7446 11406 7498
rect 11468 7446 11470 7498
rect 11308 7444 11332 7446
rect 11388 7444 11412 7446
rect 11468 7444 11492 7446
rect 11252 7424 11548 7444
rect 11060 7396 11112 7402
rect 11060 7338 11112 7344
rect 12728 7198 12756 9446
rect 12900 9300 12952 9306
rect 12900 9242 12952 9248
rect 12912 8966 12940 9242
rect 12900 8960 12952 8966
rect 12900 8902 12952 8908
rect 12716 7192 12768 7198
rect 12716 7134 12768 7140
rect 10876 6852 10928 6858
rect 10876 6794 10928 6800
rect 10600 6716 10652 6722
rect 10600 6658 10652 6664
rect 9864 6580 9916 6586
rect 9864 6522 9916 6528
rect 4388 6412 4684 6432
rect 4444 6410 4468 6412
rect 4524 6410 4548 6412
rect 4604 6410 4628 6412
rect 4466 6358 4468 6410
rect 4530 6358 4542 6410
rect 4604 6358 4606 6410
rect 4444 6356 4468 6358
rect 4524 6356 4548 6358
rect 4604 6356 4628 6358
rect 4388 6336 4684 6356
rect 11252 6412 11548 6432
rect 11308 6410 11332 6412
rect 11388 6410 11412 6412
rect 11468 6410 11492 6412
rect 11330 6358 11332 6410
rect 11394 6358 11406 6410
rect 11468 6358 11470 6410
rect 11308 6356 11332 6358
rect 11388 6356 11412 6358
rect 11468 6356 11492 6358
rect 11252 6336 11548 6356
rect 7820 5868 8116 5888
rect 7876 5866 7900 5868
rect 7956 5866 7980 5868
rect 8036 5866 8060 5868
rect 7898 5814 7900 5866
rect 7962 5814 7974 5866
rect 8036 5814 8038 5866
rect 7876 5812 7900 5814
rect 7956 5812 7980 5814
rect 8036 5812 8060 5814
rect 7820 5792 8116 5812
rect 13004 5770 13032 17878
rect 13096 17210 13124 22176
rect 13452 19024 13504 19030
rect 13452 18966 13504 18972
rect 13464 18622 13492 18966
rect 13452 18616 13504 18622
rect 13452 18558 13504 18564
rect 13096 17182 13308 17210
rect 13176 16848 13228 16854
rect 13176 16790 13228 16796
rect 13188 15970 13216 16790
rect 13176 15964 13228 15970
rect 13176 15906 13228 15912
rect 13280 9034 13308 17182
rect 13360 14808 13412 14814
rect 13360 14750 13412 14756
rect 13372 12842 13400 14750
rect 13452 13040 13504 13046
rect 13452 12982 13504 12988
rect 13360 12836 13412 12842
rect 13360 12778 13412 12784
rect 13372 11550 13400 12778
rect 13464 12706 13492 12982
rect 13452 12700 13504 12706
rect 13452 12642 13504 12648
rect 13544 12700 13596 12706
rect 13544 12642 13596 12648
rect 13452 12496 13504 12502
rect 13452 12438 13504 12444
rect 13360 11544 13412 11550
rect 13360 11486 13412 11492
rect 13464 10870 13492 12438
rect 13556 12230 13584 12642
rect 13544 12224 13596 12230
rect 13544 12166 13596 12172
rect 13452 10864 13504 10870
rect 13452 10806 13504 10812
rect 13268 9028 13320 9034
rect 13268 8970 13320 8976
rect 13544 8892 13596 8898
rect 13544 8834 13596 8840
rect 13556 8354 13584 8834
rect 13544 8348 13596 8354
rect 13544 8290 13596 8296
rect 13360 8280 13412 8286
rect 13360 8222 13412 8228
rect 13372 7946 13400 8222
rect 13360 7940 13412 7946
rect 13360 7882 13412 7888
rect 13648 6586 13676 22176
rect 13728 19024 13780 19030
rect 13728 18966 13780 18972
rect 14004 19024 14056 19030
rect 14004 18966 14056 18972
rect 13740 18758 13768 18966
rect 13728 18752 13780 18758
rect 13728 18694 13780 18700
rect 13912 18752 13964 18758
rect 13912 18694 13964 18700
rect 13728 14740 13780 14746
rect 13728 14682 13780 14688
rect 13740 14354 13768 14682
rect 13740 14338 13860 14354
rect 13740 14332 13872 14338
rect 13740 14326 13820 14332
rect 13820 14274 13872 14280
rect 13820 12632 13872 12638
rect 13820 12574 13872 12580
rect 13832 11754 13860 12574
rect 13820 11748 13872 11754
rect 13820 11690 13872 11696
rect 13728 11408 13780 11414
rect 13728 11350 13780 11356
rect 13740 11210 13768 11350
rect 13728 11204 13780 11210
rect 13728 11146 13780 11152
rect 13924 7606 13952 18694
rect 14016 18010 14044 18966
rect 14096 18820 14148 18826
rect 14096 18762 14148 18768
rect 14108 18146 14136 18762
rect 14096 18140 14148 18146
rect 14096 18082 14148 18088
rect 14004 18004 14056 18010
rect 14004 17946 14056 17952
rect 14200 17942 14228 22176
rect 14752 20202 14780 22176
rect 14568 20174 14780 20202
rect 14568 18758 14596 20174
rect 14684 20012 14980 20032
rect 14740 20010 14764 20012
rect 14820 20010 14844 20012
rect 14900 20010 14924 20012
rect 14762 19958 14764 20010
rect 14826 19958 14838 20010
rect 14900 19958 14902 20010
rect 14740 19956 14764 19958
rect 14820 19956 14844 19958
rect 14900 19956 14924 19958
rect 14684 19936 14980 19956
rect 14684 18924 14980 18944
rect 14740 18922 14764 18924
rect 14820 18922 14844 18924
rect 14900 18922 14924 18924
rect 14762 18870 14764 18922
rect 14826 18870 14838 18922
rect 14900 18870 14902 18922
rect 14740 18868 14764 18870
rect 14820 18868 14844 18870
rect 14900 18868 14924 18870
rect 14684 18848 14980 18868
rect 14556 18752 14608 18758
rect 14556 18694 14608 18700
rect 15304 17942 15332 22176
rect 15384 19228 15436 19234
rect 15384 19170 15436 19176
rect 15396 18758 15424 19170
rect 15856 19030 15884 22176
rect 15568 19024 15620 19030
rect 15568 18966 15620 18972
rect 15752 19024 15804 19030
rect 15752 18966 15804 18972
rect 15844 19024 15896 19030
rect 15844 18966 15896 18972
rect 15580 18758 15608 18966
rect 15384 18752 15436 18758
rect 15384 18694 15436 18700
rect 15568 18752 15620 18758
rect 15568 18694 15620 18700
rect 14188 17936 14240 17942
rect 14188 17878 14240 17884
rect 15016 17936 15068 17942
rect 15016 17878 15068 17884
rect 15292 17936 15344 17942
rect 15292 17878 15344 17884
rect 14684 17836 14980 17856
rect 14740 17834 14764 17836
rect 14820 17834 14844 17836
rect 14900 17834 14924 17836
rect 14762 17782 14764 17834
rect 14826 17782 14838 17834
rect 14900 17782 14902 17834
rect 14740 17780 14764 17782
rect 14820 17780 14844 17782
rect 14900 17780 14924 17782
rect 14684 17760 14980 17780
rect 14188 16984 14240 16990
rect 14188 16926 14240 16932
rect 14200 12502 14228 16926
rect 14684 16748 14980 16768
rect 14740 16746 14764 16748
rect 14820 16746 14844 16748
rect 14900 16746 14924 16748
rect 14762 16694 14764 16746
rect 14826 16694 14838 16746
rect 14900 16694 14902 16746
rect 14740 16692 14764 16694
rect 14820 16692 14844 16694
rect 14900 16692 14924 16694
rect 14684 16672 14980 16692
rect 14372 16304 14424 16310
rect 14372 16246 14424 16252
rect 14384 15970 14412 16246
rect 14372 15964 14424 15970
rect 14372 15906 14424 15912
rect 14384 14814 14412 15906
rect 14464 15760 14516 15766
rect 14464 15702 14516 15708
rect 14476 15562 14504 15702
rect 14684 15660 14980 15680
rect 14740 15658 14764 15660
rect 14820 15658 14844 15660
rect 14900 15658 14924 15660
rect 14762 15606 14764 15658
rect 14826 15606 14838 15658
rect 14900 15606 14902 15658
rect 14740 15604 14764 15606
rect 14820 15604 14844 15606
rect 14900 15604 14924 15606
rect 14684 15584 14980 15604
rect 14464 15556 14516 15562
rect 14464 15498 14516 15504
rect 14372 14808 14424 14814
rect 14372 14750 14424 14756
rect 14476 14626 14504 15498
rect 14384 14598 14504 14626
rect 14004 12496 14056 12502
rect 14004 12438 14056 12444
rect 14188 12496 14240 12502
rect 14188 12438 14240 12444
rect 14016 12230 14044 12438
rect 14200 12298 14228 12438
rect 14188 12292 14240 12298
rect 14188 12234 14240 12240
rect 14004 12224 14056 12230
rect 14004 12166 14056 12172
rect 14200 11958 14228 12234
rect 14280 12020 14332 12026
rect 14280 11962 14332 11968
rect 14004 11952 14056 11958
rect 14004 11894 14056 11900
rect 14188 11952 14240 11958
rect 14188 11894 14240 11900
rect 14016 11618 14044 11894
rect 14004 11612 14056 11618
rect 14004 11554 14056 11560
rect 14096 11612 14148 11618
rect 14096 11554 14148 11560
rect 14108 10666 14136 11554
rect 14188 11204 14240 11210
rect 14188 11146 14240 11152
rect 14200 11006 14228 11146
rect 14292 11006 14320 11962
rect 14384 11686 14412 14598
rect 14684 14572 14980 14592
rect 14740 14570 14764 14572
rect 14820 14570 14844 14572
rect 14900 14570 14924 14572
rect 14762 14518 14764 14570
rect 14826 14518 14838 14570
rect 14900 14518 14902 14570
rect 14740 14516 14764 14518
rect 14820 14516 14844 14518
rect 14900 14516 14924 14518
rect 14684 14496 14980 14516
rect 14684 13484 14980 13504
rect 14740 13482 14764 13484
rect 14820 13482 14844 13484
rect 14900 13482 14924 13484
rect 14762 13430 14764 13482
rect 14826 13430 14838 13482
rect 14900 13430 14902 13482
rect 14740 13428 14764 13430
rect 14820 13428 14844 13430
rect 14900 13428 14924 13430
rect 14684 13408 14980 13428
rect 14464 13244 14516 13250
rect 14464 13186 14516 13192
rect 14476 12570 14504 13186
rect 14556 12768 14608 12774
rect 14556 12710 14608 12716
rect 14464 12564 14516 12570
rect 14464 12506 14516 12512
rect 14372 11680 14424 11686
rect 14372 11622 14424 11628
rect 14384 11210 14412 11622
rect 14372 11204 14424 11210
rect 14372 11146 14424 11152
rect 14188 11000 14240 11006
rect 14188 10942 14240 10948
rect 14280 11000 14332 11006
rect 14280 10942 14332 10948
rect 14096 10660 14148 10666
rect 14096 10602 14148 10608
rect 14108 9374 14136 10602
rect 14200 9560 14228 10942
rect 14292 10462 14320 10942
rect 14280 10456 14332 10462
rect 14280 10398 14332 10404
rect 14200 9532 14320 9560
rect 14096 9368 14148 9374
rect 14096 9310 14148 9316
rect 14188 7736 14240 7742
rect 14188 7678 14240 7684
rect 13912 7600 13964 7606
rect 13912 7542 13964 7548
rect 14200 6858 14228 7678
rect 14188 6852 14240 6858
rect 14188 6794 14240 6800
rect 13636 6580 13688 6586
rect 13636 6522 13688 6528
rect 12992 5764 13044 5770
rect 12992 5706 13044 5712
rect 4066 5664 4122 5673
rect 4066 5599 4122 5608
rect 4388 5324 4684 5344
rect 4444 5322 4468 5324
rect 4524 5322 4548 5324
rect 4604 5322 4628 5324
rect 4466 5270 4468 5322
rect 4530 5270 4542 5322
rect 4604 5270 4606 5322
rect 4444 5268 4468 5270
rect 4524 5268 4548 5270
rect 4604 5268 4628 5270
rect 4388 5248 4684 5268
rect 11252 5324 11548 5344
rect 11308 5322 11332 5324
rect 11388 5322 11412 5324
rect 11468 5322 11492 5324
rect 11330 5270 11332 5322
rect 11394 5270 11406 5322
rect 11468 5270 11470 5322
rect 11308 5268 11332 5270
rect 11388 5268 11412 5270
rect 11468 5268 11492 5270
rect 11252 5248 11548 5268
rect 7820 4780 8116 4800
rect 7876 4778 7900 4780
rect 7956 4778 7980 4780
rect 8036 4778 8060 4780
rect 7898 4726 7900 4778
rect 7962 4726 7974 4778
rect 8036 4726 8038 4778
rect 7876 4724 7900 4726
rect 7956 4724 7980 4726
rect 8036 4724 8060 4726
rect 7820 4704 8116 4724
rect 4388 4236 4684 4256
rect 4444 4234 4468 4236
rect 4524 4234 4548 4236
rect 4604 4234 4628 4236
rect 4466 4182 4468 4234
rect 4530 4182 4542 4234
rect 4604 4182 4606 4234
rect 4444 4180 4468 4182
rect 4524 4180 4548 4182
rect 4604 4180 4628 4182
rect 4388 4160 4684 4180
rect 11252 4236 11548 4256
rect 11308 4234 11332 4236
rect 11388 4234 11412 4236
rect 11468 4234 11492 4236
rect 11330 4182 11332 4234
rect 11394 4182 11406 4234
rect 11468 4182 11470 4234
rect 11308 4180 11332 4182
rect 11388 4180 11412 4182
rect 11468 4180 11492 4182
rect 11252 4160 11548 4180
rect 14292 4002 14320 9532
rect 14372 7736 14424 7742
rect 14372 7678 14424 7684
rect 14384 7334 14412 7678
rect 14372 7328 14424 7334
rect 14372 7270 14424 7276
rect 14280 3996 14332 4002
rect 14280 3938 14332 3944
rect 7820 3692 8116 3712
rect 7876 3690 7900 3692
rect 7956 3690 7980 3692
rect 8036 3690 8060 3692
rect 7898 3638 7900 3690
rect 7962 3638 7974 3690
rect 8036 3638 8038 3690
rect 7876 3636 7900 3638
rect 7956 3636 7980 3638
rect 8036 3636 8060 3638
rect 7820 3616 8116 3636
rect 4388 3148 4684 3168
rect 4444 3146 4468 3148
rect 4524 3146 4548 3148
rect 4604 3146 4628 3148
rect 4466 3094 4468 3146
rect 4530 3094 4542 3146
rect 4604 3094 4606 3146
rect 4444 3092 4468 3094
rect 4524 3092 4548 3094
rect 4604 3092 4628 3094
rect 4388 3072 4684 3092
rect 11252 3148 11548 3168
rect 11308 3146 11332 3148
rect 11388 3146 11412 3148
rect 11468 3146 11492 3148
rect 11330 3094 11332 3146
rect 11394 3094 11406 3146
rect 11468 3094 11470 3146
rect 11308 3092 11332 3094
rect 11388 3092 11412 3094
rect 11468 3092 11492 3094
rect 11252 3072 11548 3092
rect 7820 2604 8116 2624
rect 7876 2602 7900 2604
rect 7956 2602 7980 2604
rect 8036 2602 8060 2604
rect 7898 2550 7900 2602
rect 7962 2550 7974 2602
rect 8036 2550 8038 2602
rect 7876 2548 7900 2550
rect 7956 2548 7980 2550
rect 8036 2548 8060 2550
rect 7820 2528 8116 2548
rect 14476 2506 14504 12506
rect 14568 12298 14596 12710
rect 14684 12396 14980 12416
rect 14740 12394 14764 12396
rect 14820 12394 14844 12396
rect 14900 12394 14924 12396
rect 14762 12342 14764 12394
rect 14826 12342 14838 12394
rect 14900 12342 14902 12394
rect 14740 12340 14764 12342
rect 14820 12340 14844 12342
rect 14900 12340 14924 12342
rect 14684 12320 14980 12340
rect 14556 12292 14608 12298
rect 14556 12234 14608 12240
rect 14556 11476 14608 11482
rect 14556 11418 14608 11424
rect 14568 11006 14596 11418
rect 14684 11308 14980 11328
rect 14740 11306 14764 11308
rect 14820 11306 14844 11308
rect 14900 11306 14924 11308
rect 14762 11254 14764 11306
rect 14826 11254 14838 11306
rect 14900 11254 14902 11306
rect 14740 11252 14764 11254
rect 14820 11252 14844 11254
rect 14900 11252 14924 11254
rect 14684 11232 14980 11252
rect 14556 11000 14608 11006
rect 14556 10942 14608 10948
rect 14684 10220 14980 10240
rect 14740 10218 14764 10220
rect 14820 10218 14844 10220
rect 14900 10218 14924 10220
rect 14762 10166 14764 10218
rect 14826 10166 14838 10218
rect 14900 10166 14902 10218
rect 14740 10164 14764 10166
rect 14820 10164 14844 10166
rect 14900 10164 14924 10166
rect 14684 10144 14980 10164
rect 15028 9510 15056 17878
rect 15764 17194 15792 18966
rect 16408 18554 16436 22176
rect 16764 19160 16816 19166
rect 16764 19102 16816 19108
rect 16776 18826 16804 19102
rect 16960 18826 16988 22176
rect 16764 18820 16816 18826
rect 16764 18762 16816 18768
rect 16948 18820 17000 18826
rect 16948 18762 17000 18768
rect 16580 18684 16632 18690
rect 16580 18626 16632 18632
rect 16488 18616 16540 18622
rect 16488 18558 16540 18564
rect 16396 18548 16448 18554
rect 16396 18490 16448 18496
rect 16500 18486 16528 18558
rect 16488 18480 16540 18486
rect 16488 18422 16540 18428
rect 16396 17936 16448 17942
rect 16396 17878 16448 17884
rect 15752 17188 15804 17194
rect 15752 17130 15804 17136
rect 15568 16984 15620 16990
rect 15568 16926 15620 16932
rect 15580 16582 15608 16926
rect 15568 16576 15620 16582
rect 15568 16518 15620 16524
rect 15476 16508 15528 16514
rect 15476 16450 15528 16456
rect 15488 15902 15516 16450
rect 15476 15896 15528 15902
rect 15476 15838 15528 15844
rect 15108 15420 15160 15426
rect 15108 15362 15160 15368
rect 15120 15018 15148 15362
rect 15108 15012 15160 15018
rect 15108 14954 15160 14960
rect 15200 14944 15252 14950
rect 15200 14886 15252 14892
rect 15212 14406 15240 14886
rect 15200 14400 15252 14406
rect 15200 14342 15252 14348
rect 15108 12700 15160 12706
rect 15108 12642 15160 12648
rect 15200 12700 15252 12706
rect 15200 12642 15252 12648
rect 15120 12298 15148 12642
rect 15108 12292 15160 12298
rect 15108 12234 15160 12240
rect 15212 12162 15240 12642
rect 15200 12156 15252 12162
rect 15200 12098 15252 12104
rect 15212 9986 15240 12098
rect 15764 11550 15792 17130
rect 15844 15964 15896 15970
rect 15844 15906 15896 15912
rect 15856 14950 15884 15906
rect 15844 14944 15896 14950
rect 15844 14886 15896 14892
rect 15752 11544 15804 11550
rect 15752 11486 15804 11492
rect 15200 9980 15252 9986
rect 15200 9922 15252 9928
rect 15016 9504 15068 9510
rect 15016 9446 15068 9452
rect 15292 9368 15344 9374
rect 15292 9310 15344 9316
rect 14684 9132 14980 9152
rect 14740 9130 14764 9132
rect 14820 9130 14844 9132
rect 14900 9130 14924 9132
rect 14762 9078 14764 9130
rect 14826 9078 14838 9130
rect 14900 9078 14902 9130
rect 14740 9076 14764 9078
rect 14820 9076 14844 9078
rect 14900 9076 14924 9078
rect 14684 9056 14980 9076
rect 15304 8966 15332 9310
rect 15764 9238 15792 11486
rect 15936 9980 15988 9986
rect 15936 9922 15988 9928
rect 15752 9232 15804 9238
rect 15752 9174 15804 9180
rect 15292 8960 15344 8966
rect 15292 8902 15344 8908
rect 14684 8044 14980 8064
rect 14740 8042 14764 8044
rect 14820 8042 14844 8044
rect 14900 8042 14924 8044
rect 14762 7990 14764 8042
rect 14826 7990 14838 8042
rect 14900 7990 14902 8042
rect 14740 7988 14764 7990
rect 14820 7988 14844 7990
rect 14900 7988 14924 7990
rect 14684 7968 14980 7988
rect 15948 7810 15976 9922
rect 16304 8892 16356 8898
rect 16304 8834 16356 8840
rect 16316 8490 16344 8834
rect 16304 8484 16356 8490
rect 16304 8426 16356 8432
rect 16408 8234 16436 17878
rect 16500 16582 16528 18422
rect 16592 18146 16620 18626
rect 17512 18486 17540 22176
rect 17958 21440 18014 21449
rect 17958 21375 18014 21384
rect 17972 19914 18000 21375
rect 17960 19908 18012 19914
rect 17960 19850 18012 19856
rect 17684 19772 17736 19778
rect 17684 19714 17736 19720
rect 17696 19234 17724 19714
rect 18064 19658 18092 22176
rect 18512 19772 18564 19778
rect 18512 19714 18564 19720
rect 17972 19630 18092 19658
rect 17684 19228 17736 19234
rect 17684 19170 17736 19176
rect 17972 18826 18000 19630
rect 18116 19468 18412 19488
rect 18172 19466 18196 19468
rect 18252 19466 18276 19468
rect 18332 19466 18356 19468
rect 18194 19414 18196 19466
rect 18258 19414 18270 19466
rect 18332 19414 18334 19466
rect 18172 19412 18196 19414
rect 18252 19412 18276 19414
rect 18332 19412 18356 19414
rect 18116 19392 18412 19412
rect 17960 18820 18012 18826
rect 17960 18762 18012 18768
rect 18524 18758 18552 19714
rect 18512 18752 18564 18758
rect 18512 18694 18564 18700
rect 17960 18684 18012 18690
rect 17960 18626 18012 18632
rect 17500 18480 17552 18486
rect 17500 18422 17552 18428
rect 16580 18140 16632 18146
rect 16580 18082 16632 18088
rect 16856 18072 16908 18078
rect 16856 18014 16908 18020
rect 16488 16576 16540 16582
rect 16488 16518 16540 16524
rect 16868 13794 16896 18014
rect 17040 17528 17092 17534
rect 17040 17470 17092 17476
rect 16948 16916 17000 16922
rect 16948 16858 17000 16864
rect 16960 16650 16988 16858
rect 16948 16644 17000 16650
rect 16948 16586 17000 16592
rect 16960 15970 16988 16586
rect 16948 15964 17000 15970
rect 16948 15906 17000 15912
rect 17052 15902 17080 17470
rect 17868 17392 17920 17398
rect 17868 17334 17920 17340
rect 17880 17194 17908 17334
rect 17972 17194 18000 18626
rect 18116 18380 18412 18400
rect 18172 18378 18196 18380
rect 18252 18378 18276 18380
rect 18332 18378 18356 18380
rect 18194 18326 18196 18378
rect 18258 18326 18270 18378
rect 18332 18326 18334 18378
rect 18172 18324 18196 18326
rect 18252 18324 18276 18326
rect 18332 18324 18356 18326
rect 18116 18304 18412 18324
rect 18116 17292 18412 17312
rect 18172 17290 18196 17292
rect 18252 17290 18276 17292
rect 18332 17290 18356 17292
rect 18194 17238 18196 17290
rect 18258 17238 18270 17290
rect 18332 17238 18334 17290
rect 18172 17236 18196 17238
rect 18252 17236 18276 17238
rect 18332 17236 18356 17238
rect 18116 17216 18412 17236
rect 17868 17188 17920 17194
rect 17868 17130 17920 17136
rect 17960 17188 18012 17194
rect 17960 17130 18012 17136
rect 17960 16916 18012 16922
rect 17960 16858 18012 16864
rect 17972 16106 18000 16858
rect 18052 16848 18104 16854
rect 18052 16790 18104 16796
rect 18064 16650 18092 16790
rect 18052 16644 18104 16650
rect 18052 16586 18104 16592
rect 18116 16204 18412 16224
rect 18172 16202 18196 16204
rect 18252 16202 18276 16204
rect 18332 16202 18356 16204
rect 18194 16150 18196 16202
rect 18258 16150 18270 16202
rect 18332 16150 18334 16202
rect 18172 16148 18196 16150
rect 18252 16148 18276 16150
rect 18332 16148 18356 16150
rect 18116 16128 18412 16148
rect 17960 16100 18012 16106
rect 17960 16042 18012 16048
rect 17040 15896 17092 15902
rect 17040 15838 17092 15844
rect 16948 15760 17000 15766
rect 16948 15702 17000 15708
rect 16960 15562 16988 15702
rect 16948 15556 17000 15562
rect 16948 15498 17000 15504
rect 18116 15116 18412 15136
rect 18172 15114 18196 15116
rect 18252 15114 18276 15116
rect 18332 15114 18356 15116
rect 18194 15062 18196 15114
rect 18258 15062 18270 15114
rect 18332 15062 18334 15114
rect 18172 15060 18196 15062
rect 18252 15060 18276 15062
rect 18332 15060 18356 15062
rect 18116 15040 18412 15060
rect 17040 14876 17092 14882
rect 17040 14818 17092 14824
rect 16948 14672 17000 14678
rect 16948 14614 17000 14620
rect 16960 13862 16988 14614
rect 17052 14474 17080 14818
rect 17408 14740 17460 14746
rect 17408 14682 17460 14688
rect 17040 14468 17092 14474
rect 17040 14410 17092 14416
rect 17040 14332 17092 14338
rect 17040 14274 17092 14280
rect 17132 14332 17184 14338
rect 17132 14274 17184 14280
rect 16948 13856 17000 13862
rect 16948 13798 17000 13804
rect 17052 13794 17080 14274
rect 16856 13788 16908 13794
rect 16856 13730 16908 13736
rect 17040 13788 17092 13794
rect 17040 13730 17092 13736
rect 17144 13726 17172 14274
rect 17420 13930 17448 14682
rect 17776 14264 17828 14270
rect 17776 14206 17828 14212
rect 17408 13924 17460 13930
rect 17408 13866 17460 13872
rect 17132 13720 17184 13726
rect 17132 13662 17184 13668
rect 17788 13658 17816 14206
rect 18116 14028 18412 14048
rect 18172 14026 18196 14028
rect 18252 14026 18276 14028
rect 18332 14026 18356 14028
rect 18194 13974 18196 14026
rect 18258 13974 18270 14026
rect 18332 13974 18334 14026
rect 18172 13972 18196 13974
rect 18252 13972 18276 13974
rect 18332 13972 18356 13974
rect 18116 13952 18412 13972
rect 18616 13930 18644 22176
rect 18694 21984 18750 21993
rect 18694 21919 18750 21928
rect 18708 19914 18736 21919
rect 18696 19908 18748 19914
rect 18696 19850 18748 19856
rect 18892 19166 18920 22327
rect 19154 22176 19210 22656
rect 19706 22176 19762 22656
rect 20258 22176 20314 22656
rect 20810 22176 20866 22656
rect 21362 22176 21418 22656
rect 21914 22176 21970 22656
rect 22466 22176 22522 22656
rect 18880 19160 18932 19166
rect 18880 19102 18932 19108
rect 18788 19092 18840 19098
rect 18788 19034 18840 19040
rect 18696 17460 18748 17466
rect 18696 17402 18748 17408
rect 18708 16514 18736 17402
rect 18696 16508 18748 16514
rect 18696 16450 18748 16456
rect 18800 15222 18828 19034
rect 19168 18146 19196 22176
rect 19246 21032 19302 21041
rect 19246 20967 19302 20976
rect 19260 19030 19288 20967
rect 19720 19930 19748 22176
rect 19720 19902 20116 19930
rect 19432 19772 19484 19778
rect 19432 19714 19484 19720
rect 19708 19772 19760 19778
rect 19708 19714 19760 19720
rect 19248 19024 19300 19030
rect 19248 18966 19300 18972
rect 19340 18820 19392 18826
rect 19340 18762 19392 18768
rect 19246 18720 19302 18729
rect 19246 18655 19302 18664
rect 19156 18140 19208 18146
rect 19156 18082 19208 18088
rect 18880 15896 18932 15902
rect 18880 15838 18932 15844
rect 18892 15494 18920 15838
rect 19260 15562 19288 18655
rect 19248 15556 19300 15562
rect 19248 15498 19300 15504
rect 18880 15488 18932 15494
rect 18880 15430 18932 15436
rect 18788 15216 18840 15222
rect 18788 15158 18840 15164
rect 18604 13924 18656 13930
rect 18604 13866 18656 13872
rect 17868 13856 17920 13862
rect 17868 13798 17920 13804
rect 17880 13726 17908 13798
rect 17868 13720 17920 13726
rect 17868 13662 17920 13668
rect 18420 13720 18472 13726
rect 18420 13662 18472 13668
rect 17776 13652 17828 13658
rect 17776 13594 17828 13600
rect 16764 13584 16816 13590
rect 16764 13526 16816 13532
rect 16776 11074 16804 13526
rect 17500 12564 17552 12570
rect 17500 12506 17552 12512
rect 16948 12088 17000 12094
rect 16948 12030 17000 12036
rect 16764 11068 16816 11074
rect 16764 11010 16816 11016
rect 16960 10938 16988 12030
rect 17512 11618 17540 12506
rect 17500 11612 17552 11618
rect 17500 11554 17552 11560
rect 17132 11068 17184 11074
rect 17132 11010 17184 11016
rect 17316 11068 17368 11074
rect 17316 11010 17368 11016
rect 16488 10932 16540 10938
rect 16488 10874 16540 10880
rect 16948 10932 17000 10938
rect 16948 10874 17000 10880
rect 16500 10598 16528 10874
rect 16488 10592 16540 10598
rect 16488 10534 16540 10540
rect 17144 10546 17172 11010
rect 17328 10666 17356 11010
rect 17512 11006 17540 11554
rect 17880 11074 17908 13662
rect 18432 13318 18460 13662
rect 18420 13312 18472 13318
rect 18420 13254 18472 13260
rect 18696 13244 18748 13250
rect 18696 13186 18748 13192
rect 19248 13244 19300 13250
rect 19248 13186 19300 13192
rect 18116 12940 18412 12960
rect 18172 12938 18196 12940
rect 18252 12938 18276 12940
rect 18332 12938 18356 12940
rect 18194 12886 18196 12938
rect 18258 12886 18270 12938
rect 18332 12886 18334 12938
rect 18172 12884 18196 12886
rect 18252 12884 18276 12886
rect 18332 12884 18356 12886
rect 18116 12864 18412 12884
rect 17960 12496 18012 12502
rect 17960 12438 18012 12444
rect 17972 12298 18000 12438
rect 17960 12292 18012 12298
rect 17960 12234 18012 12240
rect 17960 12156 18012 12162
rect 17960 12098 18012 12104
rect 17972 11754 18000 12098
rect 18604 11952 18656 11958
rect 18604 11894 18656 11900
rect 18116 11852 18412 11872
rect 18172 11850 18196 11852
rect 18252 11850 18276 11852
rect 18332 11850 18356 11852
rect 18194 11798 18196 11850
rect 18258 11798 18270 11850
rect 18332 11798 18334 11850
rect 18172 11796 18196 11798
rect 18252 11796 18276 11798
rect 18332 11796 18356 11798
rect 18116 11776 18412 11796
rect 17960 11748 18012 11754
rect 17960 11690 18012 11696
rect 17868 11068 17920 11074
rect 17868 11010 17920 11016
rect 17500 11000 17552 11006
rect 17500 10942 17552 10948
rect 17316 10660 17368 10666
rect 17316 10602 17368 10608
rect 16500 10054 16528 10534
rect 17144 10518 17356 10546
rect 17040 10320 17092 10326
rect 17040 10262 17092 10268
rect 16488 10048 16540 10054
rect 16488 9990 16540 9996
rect 17052 9578 17080 10262
rect 17040 9572 17092 9578
rect 17040 9514 17092 9520
rect 16408 8206 16896 8234
rect 16764 8144 16816 8150
rect 16764 8086 16816 8092
rect 16672 7940 16724 7946
rect 16672 7882 16724 7888
rect 14648 7804 14700 7810
rect 14648 7746 14700 7752
rect 15936 7804 15988 7810
rect 15936 7746 15988 7752
rect 14660 7266 14688 7746
rect 14648 7260 14700 7266
rect 14648 7202 14700 7208
rect 15948 7198 15976 7746
rect 16684 7402 16712 7882
rect 16776 7402 16804 8086
rect 16868 7878 16896 8206
rect 16856 7872 16908 7878
rect 16856 7814 16908 7820
rect 16672 7396 16724 7402
rect 16672 7338 16724 7344
rect 16764 7396 16816 7402
rect 16764 7338 16816 7344
rect 14556 7192 14608 7198
rect 14556 7134 14608 7140
rect 15936 7192 15988 7198
rect 15936 7134 15988 7140
rect 14568 6738 14596 7134
rect 14684 6956 14980 6976
rect 14740 6954 14764 6956
rect 14820 6954 14844 6956
rect 14900 6954 14924 6956
rect 14762 6902 14764 6954
rect 14826 6902 14838 6954
rect 14900 6902 14902 6954
rect 14740 6900 14764 6902
rect 14820 6900 14844 6902
rect 14900 6900 14924 6902
rect 14684 6880 14980 6900
rect 16488 6852 16540 6858
rect 16488 6794 16540 6800
rect 14568 6710 14688 6738
rect 14660 6654 14688 6710
rect 14648 6648 14700 6654
rect 14648 6590 14700 6596
rect 14684 5868 14980 5888
rect 14740 5866 14764 5868
rect 14820 5866 14844 5868
rect 14900 5866 14924 5868
rect 14762 5814 14764 5866
rect 14826 5814 14838 5866
rect 14900 5814 14902 5866
rect 14740 5812 14764 5814
rect 14820 5812 14844 5814
rect 14900 5812 14924 5814
rect 14684 5792 14980 5812
rect 16500 5226 16528 6794
rect 16488 5220 16540 5226
rect 16488 5162 16540 5168
rect 14684 4780 14980 4800
rect 14740 4778 14764 4780
rect 14820 4778 14844 4780
rect 14900 4778 14924 4780
rect 14762 4726 14764 4778
rect 14826 4726 14838 4778
rect 14900 4726 14902 4778
rect 14740 4724 14764 4726
rect 14820 4724 14844 4726
rect 14900 4724 14924 4726
rect 14684 4704 14980 4724
rect 14684 3692 14980 3712
rect 14740 3690 14764 3692
rect 14820 3690 14844 3692
rect 14900 3690 14924 3692
rect 14762 3638 14764 3690
rect 14826 3638 14838 3690
rect 14900 3638 14902 3690
rect 14740 3636 14764 3638
rect 14820 3636 14844 3638
rect 14900 3636 14924 3638
rect 14684 3616 14980 3636
rect 14684 2604 14980 2624
rect 14740 2602 14764 2604
rect 14820 2602 14844 2604
rect 14900 2602 14924 2604
rect 14762 2550 14764 2602
rect 14826 2550 14838 2602
rect 14900 2550 14902 2602
rect 14740 2548 14764 2550
rect 14820 2548 14844 2550
rect 14900 2548 14924 2550
rect 14684 2528 14980 2548
rect 14464 2500 14516 2506
rect 14464 2442 14516 2448
rect 4388 2060 4684 2080
rect 4444 2058 4468 2060
rect 4524 2058 4548 2060
rect 4604 2058 4628 2060
rect 4466 2006 4468 2058
rect 4530 2006 4542 2058
rect 4604 2006 4606 2058
rect 4444 2004 4468 2006
rect 4524 2004 4548 2006
rect 4604 2004 4628 2006
rect 4388 1984 4684 2004
rect 11252 2060 11548 2080
rect 11308 2058 11332 2060
rect 11388 2058 11412 2060
rect 11468 2058 11492 2060
rect 11330 2006 11332 2058
rect 11394 2006 11406 2058
rect 11468 2006 11470 2058
rect 11308 2004 11332 2006
rect 11388 2004 11412 2006
rect 11468 2004 11492 2006
rect 11252 1984 11548 2004
rect 17052 1214 17080 9514
rect 17040 1208 17092 1214
rect 17040 1150 17092 1156
rect 17328 97 17356 10518
rect 17512 10122 17540 10942
rect 17500 10116 17552 10122
rect 17500 10058 17552 10064
rect 17880 9034 17908 11010
rect 18512 10864 18564 10870
rect 18512 10806 18564 10812
rect 18116 10764 18412 10784
rect 18172 10762 18196 10764
rect 18252 10762 18276 10764
rect 18332 10762 18356 10764
rect 18194 10710 18196 10762
rect 18258 10710 18270 10762
rect 18332 10710 18334 10762
rect 18172 10708 18196 10710
rect 18252 10708 18276 10710
rect 18332 10708 18356 10710
rect 18116 10688 18412 10708
rect 17960 9912 18012 9918
rect 17960 9854 18012 9860
rect 17868 9028 17920 9034
rect 17868 8970 17920 8976
rect 17684 8348 17736 8354
rect 17684 8290 17736 8296
rect 17696 7946 17724 8290
rect 17684 7940 17736 7946
rect 17684 7882 17736 7888
rect 17408 7192 17460 7198
rect 17408 7134 17460 7140
rect 17420 6654 17448 7134
rect 17408 6648 17460 6654
rect 17408 6590 17460 6596
rect 17880 3633 17908 8970
rect 17972 8830 18000 9854
rect 18116 9676 18412 9696
rect 18172 9674 18196 9676
rect 18252 9674 18276 9676
rect 18332 9674 18356 9676
rect 18194 9622 18196 9674
rect 18258 9622 18270 9674
rect 18332 9622 18334 9674
rect 18172 9620 18196 9622
rect 18252 9620 18276 9622
rect 18332 9620 18356 9622
rect 18116 9600 18412 9620
rect 17960 8824 18012 8830
rect 17960 8766 18012 8772
rect 17972 7742 18000 8766
rect 18116 8588 18412 8608
rect 18172 8586 18196 8588
rect 18252 8586 18276 8588
rect 18332 8586 18356 8588
rect 18194 8534 18196 8586
rect 18258 8534 18270 8586
rect 18332 8534 18334 8586
rect 18172 8532 18196 8534
rect 18252 8532 18276 8534
rect 18332 8532 18356 8534
rect 18116 8512 18412 8532
rect 17960 7736 18012 7742
rect 17960 7678 18012 7684
rect 18116 7500 18412 7520
rect 18172 7498 18196 7500
rect 18252 7498 18276 7500
rect 18332 7498 18356 7500
rect 18194 7446 18196 7498
rect 18258 7446 18270 7498
rect 18332 7446 18334 7498
rect 18172 7444 18196 7446
rect 18252 7444 18276 7446
rect 18332 7444 18356 7446
rect 18116 7424 18412 7444
rect 18524 7418 18552 10806
rect 18616 10546 18644 11894
rect 18708 10666 18736 13186
rect 19156 12632 19208 12638
rect 19156 12574 19208 12580
rect 19168 12298 19196 12574
rect 19260 12337 19288 13186
rect 19246 12328 19302 12337
rect 19156 12292 19208 12298
rect 19246 12263 19302 12272
rect 19156 12234 19208 12240
rect 19156 11544 19208 11550
rect 19156 11486 19208 11492
rect 18788 11408 18840 11414
rect 18788 11350 18840 11356
rect 18800 11210 18828 11350
rect 18788 11204 18840 11210
rect 18788 11146 18840 11152
rect 19168 10938 19196 11486
rect 19156 10932 19208 10938
rect 19156 10874 19208 10880
rect 18696 10660 18748 10666
rect 18696 10602 18748 10608
rect 18616 10518 18828 10546
rect 18524 7390 18736 7418
rect 18512 7124 18564 7130
rect 18512 7066 18564 7072
rect 18524 6489 18552 7066
rect 18604 6716 18656 6722
rect 18604 6658 18656 6664
rect 18510 6480 18566 6489
rect 18116 6412 18412 6432
rect 18510 6415 18566 6424
rect 18172 6410 18196 6412
rect 18252 6410 18276 6412
rect 18332 6410 18356 6412
rect 18194 6358 18196 6410
rect 18258 6358 18270 6410
rect 18332 6358 18334 6410
rect 18172 6356 18196 6358
rect 18252 6356 18276 6358
rect 18332 6356 18356 6358
rect 18116 6336 18412 6356
rect 18616 5537 18644 6658
rect 18602 5528 18658 5537
rect 18602 5463 18658 5472
rect 18116 5324 18412 5344
rect 18172 5322 18196 5324
rect 18252 5322 18276 5324
rect 18332 5322 18356 5324
rect 18194 5270 18196 5322
rect 18258 5270 18270 5322
rect 18332 5270 18334 5322
rect 18172 5268 18196 5270
rect 18252 5268 18276 5270
rect 18332 5268 18356 5270
rect 18116 5248 18412 5268
rect 17960 5220 18012 5226
rect 17960 5162 18012 5168
rect 17972 4585 18000 5162
rect 17958 4576 18014 4585
rect 17958 4511 18014 4520
rect 18116 4236 18412 4256
rect 18172 4234 18196 4236
rect 18252 4234 18276 4236
rect 18332 4234 18356 4236
rect 18194 4182 18196 4234
rect 18258 4182 18270 4234
rect 18332 4182 18334 4234
rect 18172 4180 18196 4182
rect 18252 4180 18276 4182
rect 18332 4180 18356 4182
rect 18116 4160 18412 4180
rect 18512 3996 18564 4002
rect 18512 3938 18564 3944
rect 17866 3624 17922 3633
rect 17866 3559 17922 3568
rect 18524 3225 18552 3938
rect 18510 3216 18566 3225
rect 18116 3148 18412 3168
rect 18510 3151 18566 3160
rect 18172 3146 18196 3148
rect 18252 3146 18276 3148
rect 18332 3146 18356 3148
rect 18194 3094 18196 3146
rect 18258 3094 18270 3146
rect 18332 3094 18334 3146
rect 18172 3092 18196 3094
rect 18252 3092 18276 3094
rect 18332 3092 18356 3094
rect 18116 3072 18412 3092
rect 18604 2500 18656 2506
rect 18604 2442 18656 2448
rect 18116 2060 18412 2080
rect 18172 2058 18196 2060
rect 18252 2058 18276 2060
rect 18332 2058 18356 2060
rect 18194 2006 18196 2058
rect 18258 2006 18270 2058
rect 18332 2006 18334 2058
rect 18172 2004 18196 2006
rect 18252 2004 18276 2006
rect 18332 2004 18356 2006
rect 18116 1984 18412 2004
rect 18616 1457 18644 2442
rect 18602 1448 18658 1457
rect 18602 1383 18658 1392
rect 18708 505 18736 7390
rect 18800 2273 18828 10518
rect 18972 10456 19024 10462
rect 18972 10398 19024 10404
rect 18880 10320 18932 10326
rect 18880 10262 18932 10268
rect 18892 9578 18920 10262
rect 18880 9572 18932 9578
rect 18880 9514 18932 9520
rect 18984 9481 19012 10398
rect 19062 10016 19118 10025
rect 19168 10002 19196 10874
rect 19248 10864 19300 10870
rect 19248 10806 19300 10812
rect 19260 10598 19288 10806
rect 19352 10666 19380 18762
rect 19444 18010 19472 19714
rect 19524 19160 19576 19166
rect 19524 19102 19576 19108
rect 19536 18214 19564 19102
rect 19616 19092 19668 19098
rect 19616 19034 19668 19040
rect 19524 18208 19576 18214
rect 19524 18150 19576 18156
rect 19524 18072 19576 18078
rect 19524 18014 19576 18020
rect 19628 18026 19656 19034
rect 19720 18622 19748 19714
rect 19800 19704 19852 19710
rect 19800 19646 19852 19652
rect 19982 19672 20038 19681
rect 19812 18826 19840 19646
rect 19982 19607 20038 19616
rect 19800 18820 19852 18826
rect 19800 18762 19852 18768
rect 19708 18616 19760 18622
rect 19708 18558 19760 18564
rect 19892 18616 19944 18622
rect 19892 18558 19944 18564
rect 19904 18214 19932 18558
rect 19996 18282 20024 19607
rect 19984 18276 20036 18282
rect 19984 18218 20036 18224
rect 19892 18208 19944 18214
rect 19892 18150 19944 18156
rect 19800 18072 19852 18078
rect 19432 18004 19484 18010
rect 19432 17946 19484 17952
rect 19536 16582 19564 18014
rect 19628 17998 19748 18026
rect 19800 18014 19852 18020
rect 19616 17936 19668 17942
rect 19616 17878 19668 17884
rect 19524 16576 19576 16582
rect 19524 16518 19576 16524
rect 19524 15216 19576 15222
rect 19524 15158 19576 15164
rect 19536 13386 19564 15158
rect 19524 13380 19576 13386
rect 19524 13322 19576 13328
rect 19628 12026 19656 17878
rect 19720 14898 19748 17998
rect 19812 15222 19840 18014
rect 19892 17392 19944 17398
rect 19892 17334 19944 17340
rect 19904 16961 19932 17334
rect 19984 16984 20036 16990
rect 19890 16952 19946 16961
rect 19984 16926 20036 16932
rect 19890 16887 19946 16896
rect 19996 15902 20024 16926
rect 19984 15896 20036 15902
rect 19984 15838 20036 15844
rect 19984 15420 20036 15426
rect 19984 15362 20036 15368
rect 19800 15216 19852 15222
rect 19800 15158 19852 15164
rect 19890 15048 19946 15057
rect 19890 14983 19892 14992
rect 19944 14983 19946 14992
rect 19892 14954 19944 14960
rect 19720 14870 19840 14898
rect 19996 14882 20024 15362
rect 19708 14808 19760 14814
rect 19708 14750 19760 14756
rect 19720 14270 19748 14750
rect 19708 14264 19760 14270
rect 19708 14206 19760 14212
rect 19616 12020 19668 12026
rect 19616 11962 19668 11968
rect 19340 10660 19392 10666
rect 19340 10602 19392 10608
rect 19248 10592 19300 10598
rect 19248 10534 19300 10540
rect 19260 10122 19288 10534
rect 19340 10524 19392 10530
rect 19340 10466 19392 10472
rect 19248 10116 19300 10122
rect 19248 10058 19300 10064
rect 19168 9974 19288 10002
rect 19352 9986 19380 10466
rect 19708 10388 19760 10394
rect 19708 10330 19760 10336
rect 19062 9951 19118 9960
rect 18970 9472 19026 9481
rect 18970 9407 19026 9416
rect 19076 9374 19104 9951
rect 19064 9368 19116 9374
rect 19064 9310 19116 9316
rect 19156 9232 19208 9238
rect 19156 9174 19208 9180
rect 19168 7198 19196 9174
rect 19156 7192 19208 7198
rect 19156 7134 19208 7140
rect 19260 2817 19288 9974
rect 19340 9980 19392 9986
rect 19340 9922 19392 9928
rect 19352 9034 19380 9922
rect 19720 9442 19748 10330
rect 19432 9436 19484 9442
rect 19432 9378 19484 9384
rect 19708 9436 19760 9442
rect 19708 9378 19760 9384
rect 19340 9028 19392 9034
rect 19340 8970 19392 8976
rect 19444 8898 19472 9378
rect 19432 8892 19484 8898
rect 19432 8834 19484 8840
rect 19444 7946 19472 8834
rect 19812 8490 19840 14870
rect 19984 14876 20036 14882
rect 19984 14818 20036 14824
rect 19984 12156 20036 12162
rect 19984 12098 20036 12104
rect 19996 11929 20024 12098
rect 19982 11920 20038 11929
rect 19982 11855 20038 11864
rect 20088 11754 20116 19902
rect 20168 18140 20220 18146
rect 20168 18082 20220 18088
rect 20180 15986 20208 18082
rect 20272 17942 20300 22176
rect 20626 20624 20682 20633
rect 20626 20559 20682 20568
rect 20640 19914 20668 20559
rect 20718 20080 20774 20089
rect 20718 20015 20774 20024
rect 20628 19908 20680 19914
rect 20628 19850 20680 19856
rect 20732 18826 20760 20015
rect 20720 18820 20772 18826
rect 20720 18762 20772 18768
rect 20536 18548 20588 18554
rect 20536 18490 20588 18496
rect 20442 18312 20498 18321
rect 20442 18247 20498 18256
rect 20260 17936 20312 17942
rect 20260 17878 20312 17884
rect 20456 17738 20484 18247
rect 20444 17732 20496 17738
rect 20444 17674 20496 17680
rect 20260 17596 20312 17602
rect 20260 17538 20312 17544
rect 20352 17596 20404 17602
rect 20352 17538 20404 17544
rect 20272 17058 20300 17538
rect 20260 17052 20312 17058
rect 20260 16994 20312 17000
rect 20364 16582 20392 17538
rect 20548 17040 20576 18490
rect 20628 17936 20680 17942
rect 20628 17878 20680 17884
rect 20456 17012 20576 17040
rect 20352 16576 20404 16582
rect 20352 16518 20404 16524
rect 20456 16394 20484 17012
rect 20536 16916 20588 16922
rect 20536 16858 20588 16864
rect 20548 16514 20576 16858
rect 20536 16508 20588 16514
rect 20536 16450 20588 16456
rect 20456 16366 20576 16394
rect 20442 16272 20498 16281
rect 20442 16207 20498 16216
rect 20456 16106 20484 16207
rect 20444 16100 20496 16106
rect 20444 16042 20496 16048
rect 20442 16000 20498 16009
rect 20180 15958 20392 15986
rect 20168 15828 20220 15834
rect 20168 15770 20220 15776
rect 20180 14814 20208 15770
rect 20168 14808 20220 14814
rect 20168 14750 20220 14756
rect 20166 14640 20222 14649
rect 20166 14575 20222 14584
rect 20180 13386 20208 14575
rect 20364 13794 20392 15958
rect 20442 15935 20498 15944
rect 20456 15018 20484 15935
rect 20444 15012 20496 15018
rect 20444 14954 20496 14960
rect 20352 13788 20404 13794
rect 20352 13730 20404 13736
rect 20260 13720 20312 13726
rect 20548 13674 20576 16366
rect 20640 13930 20668 17878
rect 20824 16938 20852 22176
rect 21270 19264 21326 19273
rect 21270 19199 21326 19208
rect 21180 18480 21232 18486
rect 21180 18422 21232 18428
rect 21088 18004 21140 18010
rect 21088 17946 21140 17952
rect 20994 17904 21050 17913
rect 20994 17839 21050 17848
rect 21008 17738 21036 17839
rect 20996 17732 21048 17738
rect 20996 17674 21048 17680
rect 20824 16910 21036 16938
rect 20902 15592 20958 15601
rect 20902 15527 20958 15536
rect 20916 14474 20944 15527
rect 20904 14468 20956 14474
rect 20904 14410 20956 14416
rect 20810 14232 20866 14241
rect 20810 14167 20866 14176
rect 20628 13924 20680 13930
rect 20628 13866 20680 13872
rect 20628 13788 20680 13794
rect 20628 13730 20680 13736
rect 20260 13662 20312 13668
rect 20168 13380 20220 13386
rect 20168 13322 20220 13328
rect 20166 13280 20222 13289
rect 20166 13215 20222 13224
rect 20180 12842 20208 13215
rect 20272 12881 20300 13662
rect 20364 13646 20576 13674
rect 20258 12872 20314 12881
rect 20168 12836 20220 12842
rect 20258 12807 20314 12816
rect 20168 12778 20220 12784
rect 20076 11748 20128 11754
rect 20076 11690 20128 11696
rect 20260 11544 20312 11550
rect 20260 11486 20312 11492
rect 19984 11068 20036 11074
rect 19984 11010 20036 11016
rect 19996 10569 20024 11010
rect 20272 10977 20300 11486
rect 20258 10968 20314 10977
rect 20258 10903 20314 10912
rect 19982 10560 20038 10569
rect 19982 10495 20038 10504
rect 20260 10456 20312 10462
rect 20260 10398 20312 10404
rect 20272 9617 20300 10398
rect 20258 9608 20314 9617
rect 20258 9543 20314 9552
rect 20364 9034 20392 13646
rect 20536 13244 20588 13250
rect 20536 13186 20588 13192
rect 20548 12706 20576 13186
rect 20536 12700 20588 12706
rect 20536 12642 20588 12648
rect 20536 12156 20588 12162
rect 20536 12098 20588 12104
rect 20548 11521 20576 12098
rect 20534 11512 20590 11521
rect 20534 11447 20590 11456
rect 20640 11210 20668 13730
rect 20718 13688 20774 13697
rect 20718 13623 20774 13632
rect 20732 13386 20760 13623
rect 20720 13380 20772 13386
rect 20720 13322 20772 13328
rect 20824 11210 20852 14167
rect 21008 12298 21036 16910
rect 20996 12292 21048 12298
rect 20996 12234 21048 12240
rect 20628 11204 20680 11210
rect 20628 11146 20680 11152
rect 20812 11204 20864 11210
rect 20812 11146 20864 11152
rect 20536 9980 20588 9986
rect 20536 9922 20588 9928
rect 20548 9209 20576 9922
rect 20534 9200 20590 9209
rect 20534 9135 20590 9144
rect 20352 9028 20404 9034
rect 20352 8970 20404 8976
rect 19984 8892 20036 8898
rect 19984 8834 20036 8840
rect 20536 8892 20588 8898
rect 20536 8834 20588 8840
rect 19800 8484 19852 8490
rect 19800 8426 19852 8432
rect 19996 8257 20024 8834
rect 20548 8665 20576 8834
rect 20534 8656 20590 8665
rect 20534 8591 20590 8600
rect 20260 8280 20312 8286
rect 19982 8248 20038 8257
rect 20260 8222 20312 8228
rect 19982 8183 20038 8192
rect 19432 7940 19484 7946
rect 19432 7882 19484 7888
rect 20272 7849 20300 8222
rect 20258 7840 20314 7849
rect 19984 7804 20036 7810
rect 20258 7775 20314 7784
rect 20536 7804 20588 7810
rect 19984 7746 20036 7752
rect 20536 7746 20588 7752
rect 19996 6897 20024 7746
rect 20548 7305 20576 7746
rect 20534 7296 20590 7305
rect 20534 7231 20590 7240
rect 19982 6888 20038 6897
rect 19982 6823 20038 6832
rect 20536 6716 20588 6722
rect 20536 6658 20588 6664
rect 20548 5945 20576 6658
rect 20534 5936 20590 5945
rect 20534 5871 20590 5880
rect 20536 5628 20588 5634
rect 20536 5570 20588 5576
rect 20548 4993 20576 5570
rect 20534 4984 20590 4993
rect 20534 4919 20590 4928
rect 21100 4682 21128 17946
rect 21192 10122 21220 18422
rect 21284 15562 21312 19199
rect 21376 18078 21404 22176
rect 21456 18752 21508 18758
rect 21456 18694 21508 18700
rect 21364 18072 21416 18078
rect 21364 18014 21416 18020
rect 21272 15556 21324 15562
rect 21272 15498 21324 15504
rect 21180 10116 21232 10122
rect 21180 10058 21232 10064
rect 21468 9034 21496 18694
rect 21928 17942 21956 22176
rect 22480 18010 22508 22176
rect 22468 18004 22520 18010
rect 22468 17946 22520 17952
rect 21916 17936 21968 17942
rect 21916 17878 21968 17884
rect 21730 17360 21786 17369
rect 21730 17295 21732 17304
rect 21784 17295 21786 17304
rect 21732 17266 21784 17272
rect 21456 9028 21508 9034
rect 21456 8970 21508 8976
rect 21088 4676 21140 4682
rect 21088 4618 21140 4624
rect 20536 4540 20588 4546
rect 20536 4482 20588 4488
rect 20548 4177 20576 4482
rect 20534 4168 20590 4177
rect 20534 4103 20590 4112
rect 19246 2808 19302 2817
rect 19246 2743 19302 2752
rect 18786 2264 18842 2273
rect 18786 2199 18842 2208
rect 19064 1208 19116 1214
rect 19064 1150 19116 1156
rect 19076 913 19104 1150
rect 19062 904 19118 913
rect 19062 839 19118 848
rect 18694 496 18750 505
rect 18694 431 18750 440
rect 17314 88 17370 97
rect 17314 23 17370 32
<< via2 >>
rect 18878 22336 18934 22392
rect 4066 17032 4122 17088
rect 4388 19466 4444 19468
rect 4468 19466 4524 19468
rect 4548 19466 4604 19468
rect 4628 19466 4684 19468
rect 4388 19414 4414 19466
rect 4414 19414 4444 19466
rect 4468 19414 4478 19466
rect 4478 19414 4524 19466
rect 4548 19414 4594 19466
rect 4594 19414 4604 19466
rect 4628 19414 4658 19466
rect 4658 19414 4684 19466
rect 4388 19412 4444 19414
rect 4468 19412 4524 19414
rect 4548 19412 4604 19414
rect 4628 19412 4684 19414
rect 4388 18378 4444 18380
rect 4468 18378 4524 18380
rect 4548 18378 4604 18380
rect 4628 18378 4684 18380
rect 4388 18326 4414 18378
rect 4414 18326 4444 18378
rect 4468 18326 4478 18378
rect 4478 18326 4524 18378
rect 4548 18326 4594 18378
rect 4594 18326 4604 18378
rect 4628 18326 4658 18378
rect 4658 18326 4684 18378
rect 4388 18324 4444 18326
rect 4468 18324 4524 18326
rect 4548 18324 4604 18326
rect 4628 18324 4684 18326
rect 4388 17290 4444 17292
rect 4468 17290 4524 17292
rect 4548 17290 4604 17292
rect 4628 17290 4684 17292
rect 4388 17238 4414 17290
rect 4414 17238 4444 17290
rect 4468 17238 4478 17290
rect 4478 17238 4524 17290
rect 4548 17238 4594 17290
rect 4594 17238 4604 17290
rect 4628 17238 4658 17290
rect 4658 17238 4684 17290
rect 4388 17236 4444 17238
rect 4468 17236 4524 17238
rect 4548 17236 4604 17238
rect 4628 17236 4684 17238
rect 4388 16202 4444 16204
rect 4468 16202 4524 16204
rect 4548 16202 4604 16204
rect 4628 16202 4684 16204
rect 4388 16150 4414 16202
rect 4414 16150 4444 16202
rect 4468 16150 4478 16202
rect 4478 16150 4524 16202
rect 4548 16150 4594 16202
rect 4594 16150 4604 16202
rect 4628 16150 4658 16202
rect 4658 16150 4684 16202
rect 4388 16148 4444 16150
rect 4468 16148 4524 16150
rect 4548 16148 4604 16150
rect 4628 16148 4684 16150
rect 4388 15114 4444 15116
rect 4468 15114 4524 15116
rect 4548 15114 4604 15116
rect 4628 15114 4684 15116
rect 4388 15062 4414 15114
rect 4414 15062 4444 15114
rect 4468 15062 4478 15114
rect 4478 15062 4524 15114
rect 4548 15062 4594 15114
rect 4594 15062 4604 15114
rect 4628 15062 4658 15114
rect 4658 15062 4684 15114
rect 4388 15060 4444 15062
rect 4468 15060 4524 15062
rect 4548 15060 4604 15062
rect 4628 15060 4684 15062
rect 4388 14026 4444 14028
rect 4468 14026 4524 14028
rect 4548 14026 4604 14028
rect 4628 14026 4684 14028
rect 4388 13974 4414 14026
rect 4414 13974 4444 14026
rect 4468 13974 4478 14026
rect 4478 13974 4524 14026
rect 4548 13974 4594 14026
rect 4594 13974 4604 14026
rect 4628 13974 4658 14026
rect 4658 13974 4684 14026
rect 4388 13972 4444 13974
rect 4468 13972 4524 13974
rect 4548 13972 4604 13974
rect 4628 13972 4684 13974
rect 7820 20010 7876 20012
rect 7900 20010 7956 20012
rect 7980 20010 8036 20012
rect 8060 20010 8116 20012
rect 7820 19958 7846 20010
rect 7846 19958 7876 20010
rect 7900 19958 7910 20010
rect 7910 19958 7956 20010
rect 7980 19958 8026 20010
rect 8026 19958 8036 20010
rect 8060 19958 8090 20010
rect 8090 19958 8116 20010
rect 7820 19956 7876 19958
rect 7900 19956 7956 19958
rect 7980 19956 8036 19958
rect 8060 19956 8116 19958
rect 7820 18922 7876 18924
rect 7900 18922 7956 18924
rect 7980 18922 8036 18924
rect 8060 18922 8116 18924
rect 7820 18870 7846 18922
rect 7846 18870 7876 18922
rect 7900 18870 7910 18922
rect 7910 18870 7956 18922
rect 7980 18870 8026 18922
rect 8026 18870 8036 18922
rect 8060 18870 8090 18922
rect 8090 18870 8116 18922
rect 7820 18868 7876 18870
rect 7900 18868 7956 18870
rect 7980 18868 8036 18870
rect 8060 18868 8116 18870
rect 7820 17834 7876 17836
rect 7900 17834 7956 17836
rect 7980 17834 8036 17836
rect 8060 17834 8116 17836
rect 7820 17782 7846 17834
rect 7846 17782 7876 17834
rect 7900 17782 7910 17834
rect 7910 17782 7956 17834
rect 7980 17782 8026 17834
rect 8026 17782 8036 17834
rect 8060 17782 8090 17834
rect 8090 17782 8116 17834
rect 7820 17780 7876 17782
rect 7900 17780 7956 17782
rect 7980 17780 8036 17782
rect 8060 17780 8116 17782
rect 7820 16746 7876 16748
rect 7900 16746 7956 16748
rect 7980 16746 8036 16748
rect 8060 16746 8116 16748
rect 7820 16694 7846 16746
rect 7846 16694 7876 16746
rect 7900 16694 7910 16746
rect 7910 16694 7956 16746
rect 7980 16694 8026 16746
rect 8026 16694 8036 16746
rect 8060 16694 8090 16746
rect 8090 16694 8116 16746
rect 7820 16692 7876 16694
rect 7900 16692 7956 16694
rect 7980 16692 8036 16694
rect 8060 16692 8116 16694
rect 7820 15658 7876 15660
rect 7900 15658 7956 15660
rect 7980 15658 8036 15660
rect 8060 15658 8116 15660
rect 7820 15606 7846 15658
rect 7846 15606 7876 15658
rect 7900 15606 7910 15658
rect 7910 15606 7956 15658
rect 7980 15606 8026 15658
rect 8026 15606 8036 15658
rect 8060 15606 8090 15658
rect 8090 15606 8116 15658
rect 7820 15604 7876 15606
rect 7900 15604 7956 15606
rect 7980 15604 8036 15606
rect 8060 15604 8116 15606
rect 7820 14570 7876 14572
rect 7900 14570 7956 14572
rect 7980 14570 8036 14572
rect 8060 14570 8116 14572
rect 7820 14518 7846 14570
rect 7846 14518 7876 14570
rect 7900 14518 7910 14570
rect 7910 14518 7956 14570
rect 7980 14518 8026 14570
rect 8026 14518 8036 14570
rect 8060 14518 8090 14570
rect 8090 14518 8116 14570
rect 7820 14516 7876 14518
rect 7900 14516 7956 14518
rect 7980 14516 8036 14518
rect 8060 14516 8116 14518
rect 4388 12938 4444 12940
rect 4468 12938 4524 12940
rect 4548 12938 4604 12940
rect 4628 12938 4684 12940
rect 4388 12886 4414 12938
rect 4414 12886 4444 12938
rect 4468 12886 4478 12938
rect 4478 12886 4524 12938
rect 4548 12886 4594 12938
rect 4594 12886 4604 12938
rect 4628 12886 4658 12938
rect 4658 12886 4684 12938
rect 4388 12884 4444 12886
rect 4468 12884 4524 12886
rect 4548 12884 4604 12886
rect 4628 12884 4684 12886
rect 4388 11850 4444 11852
rect 4468 11850 4524 11852
rect 4548 11850 4604 11852
rect 4628 11850 4684 11852
rect 4388 11798 4414 11850
rect 4414 11798 4444 11850
rect 4468 11798 4478 11850
rect 4478 11798 4524 11850
rect 4548 11798 4594 11850
rect 4594 11798 4604 11850
rect 4628 11798 4658 11850
rect 4658 11798 4684 11850
rect 4388 11796 4444 11798
rect 4468 11796 4524 11798
rect 4548 11796 4604 11798
rect 4628 11796 4684 11798
rect 7820 13482 7876 13484
rect 7900 13482 7956 13484
rect 7980 13482 8036 13484
rect 8060 13482 8116 13484
rect 7820 13430 7846 13482
rect 7846 13430 7876 13482
rect 7900 13430 7910 13482
rect 7910 13430 7956 13482
rect 7980 13430 8026 13482
rect 8026 13430 8036 13482
rect 8060 13430 8090 13482
rect 8090 13430 8116 13482
rect 7820 13428 7876 13430
rect 7900 13428 7956 13430
rect 7980 13428 8036 13430
rect 8060 13428 8116 13430
rect 7820 12394 7876 12396
rect 7900 12394 7956 12396
rect 7980 12394 8036 12396
rect 8060 12394 8116 12396
rect 7820 12342 7846 12394
rect 7846 12342 7876 12394
rect 7900 12342 7910 12394
rect 7910 12342 7956 12394
rect 7980 12342 8026 12394
rect 8026 12342 8036 12394
rect 8060 12342 8090 12394
rect 8090 12342 8116 12394
rect 7820 12340 7876 12342
rect 7900 12340 7956 12342
rect 7980 12340 8036 12342
rect 8060 12340 8116 12342
rect 4388 10762 4444 10764
rect 4468 10762 4524 10764
rect 4548 10762 4604 10764
rect 4628 10762 4684 10764
rect 4388 10710 4414 10762
rect 4414 10710 4444 10762
rect 4468 10710 4478 10762
rect 4478 10710 4524 10762
rect 4548 10710 4594 10762
rect 4594 10710 4604 10762
rect 4628 10710 4658 10762
rect 4658 10710 4684 10762
rect 4388 10708 4444 10710
rect 4468 10708 4524 10710
rect 4548 10708 4604 10710
rect 4628 10708 4684 10710
rect 7820 11306 7876 11308
rect 7900 11306 7956 11308
rect 7980 11306 8036 11308
rect 8060 11306 8116 11308
rect 7820 11254 7846 11306
rect 7846 11254 7876 11306
rect 7900 11254 7910 11306
rect 7910 11254 7956 11306
rect 7980 11254 8026 11306
rect 8026 11254 8036 11306
rect 8060 11254 8090 11306
rect 8090 11254 8116 11306
rect 7820 11252 7876 11254
rect 7900 11252 7956 11254
rect 7980 11252 8036 11254
rect 8060 11252 8116 11254
rect 4388 9674 4444 9676
rect 4468 9674 4524 9676
rect 4548 9674 4604 9676
rect 4628 9674 4684 9676
rect 4388 9622 4414 9674
rect 4414 9622 4444 9674
rect 4468 9622 4478 9674
rect 4478 9622 4524 9674
rect 4548 9622 4594 9674
rect 4594 9622 4604 9674
rect 4628 9622 4658 9674
rect 4658 9622 4684 9674
rect 4388 9620 4444 9622
rect 4468 9620 4524 9622
rect 4548 9620 4604 9622
rect 4628 9620 4684 9622
rect 7820 10218 7876 10220
rect 7900 10218 7956 10220
rect 7980 10218 8036 10220
rect 8060 10218 8116 10220
rect 7820 10166 7846 10218
rect 7846 10166 7876 10218
rect 7900 10166 7910 10218
rect 7910 10166 7956 10218
rect 7980 10166 8026 10218
rect 8026 10166 8036 10218
rect 8060 10166 8090 10218
rect 8090 10166 8116 10218
rect 7820 10164 7876 10166
rect 7900 10164 7956 10166
rect 7980 10164 8036 10166
rect 8060 10164 8116 10166
rect 7820 9130 7876 9132
rect 7900 9130 7956 9132
rect 7980 9130 8036 9132
rect 8060 9130 8116 9132
rect 7820 9078 7846 9130
rect 7846 9078 7876 9130
rect 7900 9078 7910 9130
rect 7910 9078 7956 9130
rect 7980 9078 8026 9130
rect 8026 9078 8036 9130
rect 8060 9078 8090 9130
rect 8090 9078 8116 9130
rect 7820 9076 7876 9078
rect 7900 9076 7956 9078
rect 7980 9076 8036 9078
rect 8060 9076 8116 9078
rect 4388 8586 4444 8588
rect 4468 8586 4524 8588
rect 4548 8586 4604 8588
rect 4628 8586 4684 8588
rect 4388 8534 4414 8586
rect 4414 8534 4444 8586
rect 4468 8534 4478 8586
rect 4478 8534 4524 8586
rect 4548 8534 4594 8586
rect 4594 8534 4604 8586
rect 4628 8534 4658 8586
rect 4658 8534 4684 8586
rect 4388 8532 4444 8534
rect 4468 8532 4524 8534
rect 4548 8532 4604 8534
rect 4628 8532 4684 8534
rect 7820 8042 7876 8044
rect 7900 8042 7956 8044
rect 7980 8042 8036 8044
rect 8060 8042 8116 8044
rect 7820 7990 7846 8042
rect 7846 7990 7876 8042
rect 7900 7990 7910 8042
rect 7910 7990 7956 8042
rect 7980 7990 8026 8042
rect 8026 7990 8036 8042
rect 8060 7990 8090 8042
rect 8090 7990 8116 8042
rect 7820 7988 7876 7990
rect 7900 7988 7956 7990
rect 7980 7988 8036 7990
rect 8060 7988 8116 7990
rect 4388 7498 4444 7500
rect 4468 7498 4524 7500
rect 4548 7498 4604 7500
rect 4628 7498 4684 7500
rect 4388 7446 4414 7498
rect 4414 7446 4444 7498
rect 4468 7446 4478 7498
rect 4478 7446 4524 7498
rect 4548 7446 4594 7498
rect 4594 7446 4604 7498
rect 4628 7446 4658 7498
rect 4658 7446 4684 7498
rect 4388 7444 4444 7446
rect 4468 7444 4524 7446
rect 4548 7444 4604 7446
rect 4628 7444 4684 7446
rect 7820 6954 7876 6956
rect 7900 6954 7956 6956
rect 7980 6954 8036 6956
rect 8060 6954 8116 6956
rect 7820 6902 7846 6954
rect 7846 6902 7876 6954
rect 7900 6902 7910 6954
rect 7910 6902 7956 6954
rect 7980 6902 8026 6954
rect 8026 6902 8036 6954
rect 8060 6902 8090 6954
rect 8090 6902 8116 6954
rect 7820 6900 7876 6902
rect 7900 6900 7956 6902
rect 7980 6900 8036 6902
rect 8060 6900 8116 6902
rect 11252 19466 11308 19468
rect 11332 19466 11388 19468
rect 11412 19466 11468 19468
rect 11492 19466 11548 19468
rect 11252 19414 11278 19466
rect 11278 19414 11308 19466
rect 11332 19414 11342 19466
rect 11342 19414 11388 19466
rect 11412 19414 11458 19466
rect 11458 19414 11468 19466
rect 11492 19414 11522 19466
rect 11522 19414 11548 19466
rect 11252 19412 11308 19414
rect 11332 19412 11388 19414
rect 11412 19412 11468 19414
rect 11492 19412 11548 19414
rect 11252 18378 11308 18380
rect 11332 18378 11388 18380
rect 11412 18378 11468 18380
rect 11492 18378 11548 18380
rect 11252 18326 11278 18378
rect 11278 18326 11308 18378
rect 11332 18326 11342 18378
rect 11342 18326 11388 18378
rect 11412 18326 11458 18378
rect 11458 18326 11468 18378
rect 11492 18326 11522 18378
rect 11522 18326 11548 18378
rect 11252 18324 11308 18326
rect 11332 18324 11388 18326
rect 11412 18324 11468 18326
rect 11492 18324 11548 18326
rect 11252 17290 11308 17292
rect 11332 17290 11388 17292
rect 11412 17290 11468 17292
rect 11492 17290 11548 17292
rect 11252 17238 11278 17290
rect 11278 17238 11308 17290
rect 11332 17238 11342 17290
rect 11342 17238 11388 17290
rect 11412 17238 11458 17290
rect 11458 17238 11468 17290
rect 11492 17238 11522 17290
rect 11522 17238 11548 17290
rect 11252 17236 11308 17238
rect 11332 17236 11388 17238
rect 11412 17236 11468 17238
rect 11492 17236 11548 17238
rect 11252 16202 11308 16204
rect 11332 16202 11388 16204
rect 11412 16202 11468 16204
rect 11492 16202 11548 16204
rect 11252 16150 11278 16202
rect 11278 16150 11308 16202
rect 11332 16150 11342 16202
rect 11342 16150 11388 16202
rect 11412 16150 11458 16202
rect 11458 16150 11468 16202
rect 11492 16150 11522 16202
rect 11522 16150 11548 16202
rect 11252 16148 11308 16150
rect 11332 16148 11388 16150
rect 11412 16148 11468 16150
rect 11492 16148 11548 16150
rect 11252 15114 11308 15116
rect 11332 15114 11388 15116
rect 11412 15114 11468 15116
rect 11492 15114 11548 15116
rect 11252 15062 11278 15114
rect 11278 15062 11308 15114
rect 11332 15062 11342 15114
rect 11342 15062 11388 15114
rect 11412 15062 11458 15114
rect 11458 15062 11468 15114
rect 11492 15062 11522 15114
rect 11522 15062 11548 15114
rect 11252 15060 11308 15062
rect 11332 15060 11388 15062
rect 11412 15060 11468 15062
rect 11492 15060 11548 15062
rect 11252 14026 11308 14028
rect 11332 14026 11388 14028
rect 11412 14026 11468 14028
rect 11492 14026 11548 14028
rect 11252 13974 11278 14026
rect 11278 13974 11308 14026
rect 11332 13974 11342 14026
rect 11342 13974 11388 14026
rect 11412 13974 11458 14026
rect 11458 13974 11468 14026
rect 11492 13974 11522 14026
rect 11522 13974 11548 14026
rect 11252 13972 11308 13974
rect 11332 13972 11388 13974
rect 11412 13972 11468 13974
rect 11492 13972 11548 13974
rect 11252 12938 11308 12940
rect 11332 12938 11388 12940
rect 11412 12938 11468 12940
rect 11492 12938 11548 12940
rect 11252 12886 11278 12938
rect 11278 12886 11308 12938
rect 11332 12886 11342 12938
rect 11342 12886 11388 12938
rect 11412 12886 11458 12938
rect 11458 12886 11468 12938
rect 11492 12886 11522 12938
rect 11522 12886 11548 12938
rect 11252 12884 11308 12886
rect 11332 12884 11388 12886
rect 11412 12884 11468 12886
rect 11492 12884 11548 12886
rect 11252 11850 11308 11852
rect 11332 11850 11388 11852
rect 11412 11850 11468 11852
rect 11492 11850 11548 11852
rect 11252 11798 11278 11850
rect 11278 11798 11308 11850
rect 11332 11798 11342 11850
rect 11342 11798 11388 11850
rect 11412 11798 11458 11850
rect 11458 11798 11468 11850
rect 11492 11798 11522 11850
rect 11522 11798 11548 11850
rect 11252 11796 11308 11798
rect 11332 11796 11388 11798
rect 11412 11796 11468 11798
rect 11492 11796 11548 11798
rect 11252 10762 11308 10764
rect 11332 10762 11388 10764
rect 11412 10762 11468 10764
rect 11492 10762 11548 10764
rect 11252 10710 11278 10762
rect 11278 10710 11308 10762
rect 11332 10710 11342 10762
rect 11342 10710 11388 10762
rect 11412 10710 11458 10762
rect 11458 10710 11468 10762
rect 11492 10710 11522 10762
rect 11522 10710 11548 10762
rect 11252 10708 11308 10710
rect 11332 10708 11388 10710
rect 11412 10708 11468 10710
rect 11492 10708 11548 10710
rect 11252 9674 11308 9676
rect 11332 9674 11388 9676
rect 11412 9674 11468 9676
rect 11492 9674 11548 9676
rect 11252 9622 11278 9674
rect 11278 9622 11308 9674
rect 11332 9622 11342 9674
rect 11342 9622 11388 9674
rect 11412 9622 11458 9674
rect 11458 9622 11468 9674
rect 11492 9622 11522 9674
rect 11522 9622 11548 9674
rect 11252 9620 11308 9622
rect 11332 9620 11388 9622
rect 11412 9620 11468 9622
rect 11492 9620 11548 9622
rect 11252 8586 11308 8588
rect 11332 8586 11388 8588
rect 11412 8586 11468 8588
rect 11492 8586 11548 8588
rect 11252 8534 11278 8586
rect 11278 8534 11308 8586
rect 11332 8534 11342 8586
rect 11342 8534 11388 8586
rect 11412 8534 11458 8586
rect 11458 8534 11468 8586
rect 11492 8534 11522 8586
rect 11522 8534 11548 8586
rect 11252 8532 11308 8534
rect 11332 8532 11388 8534
rect 11412 8532 11468 8534
rect 11492 8532 11548 8534
rect 11252 7498 11308 7500
rect 11332 7498 11388 7500
rect 11412 7498 11468 7500
rect 11492 7498 11548 7500
rect 11252 7446 11278 7498
rect 11278 7446 11308 7498
rect 11332 7446 11342 7498
rect 11342 7446 11388 7498
rect 11412 7446 11458 7498
rect 11458 7446 11468 7498
rect 11492 7446 11522 7498
rect 11522 7446 11548 7498
rect 11252 7444 11308 7446
rect 11332 7444 11388 7446
rect 11412 7444 11468 7446
rect 11492 7444 11548 7446
rect 4388 6410 4444 6412
rect 4468 6410 4524 6412
rect 4548 6410 4604 6412
rect 4628 6410 4684 6412
rect 4388 6358 4414 6410
rect 4414 6358 4444 6410
rect 4468 6358 4478 6410
rect 4478 6358 4524 6410
rect 4548 6358 4594 6410
rect 4594 6358 4604 6410
rect 4628 6358 4658 6410
rect 4658 6358 4684 6410
rect 4388 6356 4444 6358
rect 4468 6356 4524 6358
rect 4548 6356 4604 6358
rect 4628 6356 4684 6358
rect 11252 6410 11308 6412
rect 11332 6410 11388 6412
rect 11412 6410 11468 6412
rect 11492 6410 11548 6412
rect 11252 6358 11278 6410
rect 11278 6358 11308 6410
rect 11332 6358 11342 6410
rect 11342 6358 11388 6410
rect 11412 6358 11458 6410
rect 11458 6358 11468 6410
rect 11492 6358 11522 6410
rect 11522 6358 11548 6410
rect 11252 6356 11308 6358
rect 11332 6356 11388 6358
rect 11412 6356 11468 6358
rect 11492 6356 11548 6358
rect 7820 5866 7876 5868
rect 7900 5866 7956 5868
rect 7980 5866 8036 5868
rect 8060 5866 8116 5868
rect 7820 5814 7846 5866
rect 7846 5814 7876 5866
rect 7900 5814 7910 5866
rect 7910 5814 7956 5866
rect 7980 5814 8026 5866
rect 8026 5814 8036 5866
rect 8060 5814 8090 5866
rect 8090 5814 8116 5866
rect 7820 5812 7876 5814
rect 7900 5812 7956 5814
rect 7980 5812 8036 5814
rect 8060 5812 8116 5814
rect 14684 20010 14740 20012
rect 14764 20010 14820 20012
rect 14844 20010 14900 20012
rect 14924 20010 14980 20012
rect 14684 19958 14710 20010
rect 14710 19958 14740 20010
rect 14764 19958 14774 20010
rect 14774 19958 14820 20010
rect 14844 19958 14890 20010
rect 14890 19958 14900 20010
rect 14924 19958 14954 20010
rect 14954 19958 14980 20010
rect 14684 19956 14740 19958
rect 14764 19956 14820 19958
rect 14844 19956 14900 19958
rect 14924 19956 14980 19958
rect 14684 18922 14740 18924
rect 14764 18922 14820 18924
rect 14844 18922 14900 18924
rect 14924 18922 14980 18924
rect 14684 18870 14710 18922
rect 14710 18870 14740 18922
rect 14764 18870 14774 18922
rect 14774 18870 14820 18922
rect 14844 18870 14890 18922
rect 14890 18870 14900 18922
rect 14924 18870 14954 18922
rect 14954 18870 14980 18922
rect 14684 18868 14740 18870
rect 14764 18868 14820 18870
rect 14844 18868 14900 18870
rect 14924 18868 14980 18870
rect 14684 17834 14740 17836
rect 14764 17834 14820 17836
rect 14844 17834 14900 17836
rect 14924 17834 14980 17836
rect 14684 17782 14710 17834
rect 14710 17782 14740 17834
rect 14764 17782 14774 17834
rect 14774 17782 14820 17834
rect 14844 17782 14890 17834
rect 14890 17782 14900 17834
rect 14924 17782 14954 17834
rect 14954 17782 14980 17834
rect 14684 17780 14740 17782
rect 14764 17780 14820 17782
rect 14844 17780 14900 17782
rect 14924 17780 14980 17782
rect 14684 16746 14740 16748
rect 14764 16746 14820 16748
rect 14844 16746 14900 16748
rect 14924 16746 14980 16748
rect 14684 16694 14710 16746
rect 14710 16694 14740 16746
rect 14764 16694 14774 16746
rect 14774 16694 14820 16746
rect 14844 16694 14890 16746
rect 14890 16694 14900 16746
rect 14924 16694 14954 16746
rect 14954 16694 14980 16746
rect 14684 16692 14740 16694
rect 14764 16692 14820 16694
rect 14844 16692 14900 16694
rect 14924 16692 14980 16694
rect 14684 15658 14740 15660
rect 14764 15658 14820 15660
rect 14844 15658 14900 15660
rect 14924 15658 14980 15660
rect 14684 15606 14710 15658
rect 14710 15606 14740 15658
rect 14764 15606 14774 15658
rect 14774 15606 14820 15658
rect 14844 15606 14890 15658
rect 14890 15606 14900 15658
rect 14924 15606 14954 15658
rect 14954 15606 14980 15658
rect 14684 15604 14740 15606
rect 14764 15604 14820 15606
rect 14844 15604 14900 15606
rect 14924 15604 14980 15606
rect 14684 14570 14740 14572
rect 14764 14570 14820 14572
rect 14844 14570 14900 14572
rect 14924 14570 14980 14572
rect 14684 14518 14710 14570
rect 14710 14518 14740 14570
rect 14764 14518 14774 14570
rect 14774 14518 14820 14570
rect 14844 14518 14890 14570
rect 14890 14518 14900 14570
rect 14924 14518 14954 14570
rect 14954 14518 14980 14570
rect 14684 14516 14740 14518
rect 14764 14516 14820 14518
rect 14844 14516 14900 14518
rect 14924 14516 14980 14518
rect 14684 13482 14740 13484
rect 14764 13482 14820 13484
rect 14844 13482 14900 13484
rect 14924 13482 14980 13484
rect 14684 13430 14710 13482
rect 14710 13430 14740 13482
rect 14764 13430 14774 13482
rect 14774 13430 14820 13482
rect 14844 13430 14890 13482
rect 14890 13430 14900 13482
rect 14924 13430 14954 13482
rect 14954 13430 14980 13482
rect 14684 13428 14740 13430
rect 14764 13428 14820 13430
rect 14844 13428 14900 13430
rect 14924 13428 14980 13430
rect 4066 5608 4122 5664
rect 4388 5322 4444 5324
rect 4468 5322 4524 5324
rect 4548 5322 4604 5324
rect 4628 5322 4684 5324
rect 4388 5270 4414 5322
rect 4414 5270 4444 5322
rect 4468 5270 4478 5322
rect 4478 5270 4524 5322
rect 4548 5270 4594 5322
rect 4594 5270 4604 5322
rect 4628 5270 4658 5322
rect 4658 5270 4684 5322
rect 4388 5268 4444 5270
rect 4468 5268 4524 5270
rect 4548 5268 4604 5270
rect 4628 5268 4684 5270
rect 11252 5322 11308 5324
rect 11332 5322 11388 5324
rect 11412 5322 11468 5324
rect 11492 5322 11548 5324
rect 11252 5270 11278 5322
rect 11278 5270 11308 5322
rect 11332 5270 11342 5322
rect 11342 5270 11388 5322
rect 11412 5270 11458 5322
rect 11458 5270 11468 5322
rect 11492 5270 11522 5322
rect 11522 5270 11548 5322
rect 11252 5268 11308 5270
rect 11332 5268 11388 5270
rect 11412 5268 11468 5270
rect 11492 5268 11548 5270
rect 7820 4778 7876 4780
rect 7900 4778 7956 4780
rect 7980 4778 8036 4780
rect 8060 4778 8116 4780
rect 7820 4726 7846 4778
rect 7846 4726 7876 4778
rect 7900 4726 7910 4778
rect 7910 4726 7956 4778
rect 7980 4726 8026 4778
rect 8026 4726 8036 4778
rect 8060 4726 8090 4778
rect 8090 4726 8116 4778
rect 7820 4724 7876 4726
rect 7900 4724 7956 4726
rect 7980 4724 8036 4726
rect 8060 4724 8116 4726
rect 4388 4234 4444 4236
rect 4468 4234 4524 4236
rect 4548 4234 4604 4236
rect 4628 4234 4684 4236
rect 4388 4182 4414 4234
rect 4414 4182 4444 4234
rect 4468 4182 4478 4234
rect 4478 4182 4524 4234
rect 4548 4182 4594 4234
rect 4594 4182 4604 4234
rect 4628 4182 4658 4234
rect 4658 4182 4684 4234
rect 4388 4180 4444 4182
rect 4468 4180 4524 4182
rect 4548 4180 4604 4182
rect 4628 4180 4684 4182
rect 11252 4234 11308 4236
rect 11332 4234 11388 4236
rect 11412 4234 11468 4236
rect 11492 4234 11548 4236
rect 11252 4182 11278 4234
rect 11278 4182 11308 4234
rect 11332 4182 11342 4234
rect 11342 4182 11388 4234
rect 11412 4182 11458 4234
rect 11458 4182 11468 4234
rect 11492 4182 11522 4234
rect 11522 4182 11548 4234
rect 11252 4180 11308 4182
rect 11332 4180 11388 4182
rect 11412 4180 11468 4182
rect 11492 4180 11548 4182
rect 7820 3690 7876 3692
rect 7900 3690 7956 3692
rect 7980 3690 8036 3692
rect 8060 3690 8116 3692
rect 7820 3638 7846 3690
rect 7846 3638 7876 3690
rect 7900 3638 7910 3690
rect 7910 3638 7956 3690
rect 7980 3638 8026 3690
rect 8026 3638 8036 3690
rect 8060 3638 8090 3690
rect 8090 3638 8116 3690
rect 7820 3636 7876 3638
rect 7900 3636 7956 3638
rect 7980 3636 8036 3638
rect 8060 3636 8116 3638
rect 4388 3146 4444 3148
rect 4468 3146 4524 3148
rect 4548 3146 4604 3148
rect 4628 3146 4684 3148
rect 4388 3094 4414 3146
rect 4414 3094 4444 3146
rect 4468 3094 4478 3146
rect 4478 3094 4524 3146
rect 4548 3094 4594 3146
rect 4594 3094 4604 3146
rect 4628 3094 4658 3146
rect 4658 3094 4684 3146
rect 4388 3092 4444 3094
rect 4468 3092 4524 3094
rect 4548 3092 4604 3094
rect 4628 3092 4684 3094
rect 11252 3146 11308 3148
rect 11332 3146 11388 3148
rect 11412 3146 11468 3148
rect 11492 3146 11548 3148
rect 11252 3094 11278 3146
rect 11278 3094 11308 3146
rect 11332 3094 11342 3146
rect 11342 3094 11388 3146
rect 11412 3094 11458 3146
rect 11458 3094 11468 3146
rect 11492 3094 11522 3146
rect 11522 3094 11548 3146
rect 11252 3092 11308 3094
rect 11332 3092 11388 3094
rect 11412 3092 11468 3094
rect 11492 3092 11548 3094
rect 7820 2602 7876 2604
rect 7900 2602 7956 2604
rect 7980 2602 8036 2604
rect 8060 2602 8116 2604
rect 7820 2550 7846 2602
rect 7846 2550 7876 2602
rect 7900 2550 7910 2602
rect 7910 2550 7956 2602
rect 7980 2550 8026 2602
rect 8026 2550 8036 2602
rect 8060 2550 8090 2602
rect 8090 2550 8116 2602
rect 7820 2548 7876 2550
rect 7900 2548 7956 2550
rect 7980 2548 8036 2550
rect 8060 2548 8116 2550
rect 14684 12394 14740 12396
rect 14764 12394 14820 12396
rect 14844 12394 14900 12396
rect 14924 12394 14980 12396
rect 14684 12342 14710 12394
rect 14710 12342 14740 12394
rect 14764 12342 14774 12394
rect 14774 12342 14820 12394
rect 14844 12342 14890 12394
rect 14890 12342 14900 12394
rect 14924 12342 14954 12394
rect 14954 12342 14980 12394
rect 14684 12340 14740 12342
rect 14764 12340 14820 12342
rect 14844 12340 14900 12342
rect 14924 12340 14980 12342
rect 14684 11306 14740 11308
rect 14764 11306 14820 11308
rect 14844 11306 14900 11308
rect 14924 11306 14980 11308
rect 14684 11254 14710 11306
rect 14710 11254 14740 11306
rect 14764 11254 14774 11306
rect 14774 11254 14820 11306
rect 14844 11254 14890 11306
rect 14890 11254 14900 11306
rect 14924 11254 14954 11306
rect 14954 11254 14980 11306
rect 14684 11252 14740 11254
rect 14764 11252 14820 11254
rect 14844 11252 14900 11254
rect 14924 11252 14980 11254
rect 14684 10218 14740 10220
rect 14764 10218 14820 10220
rect 14844 10218 14900 10220
rect 14924 10218 14980 10220
rect 14684 10166 14710 10218
rect 14710 10166 14740 10218
rect 14764 10166 14774 10218
rect 14774 10166 14820 10218
rect 14844 10166 14890 10218
rect 14890 10166 14900 10218
rect 14924 10166 14954 10218
rect 14954 10166 14980 10218
rect 14684 10164 14740 10166
rect 14764 10164 14820 10166
rect 14844 10164 14900 10166
rect 14924 10164 14980 10166
rect 14684 9130 14740 9132
rect 14764 9130 14820 9132
rect 14844 9130 14900 9132
rect 14924 9130 14980 9132
rect 14684 9078 14710 9130
rect 14710 9078 14740 9130
rect 14764 9078 14774 9130
rect 14774 9078 14820 9130
rect 14844 9078 14890 9130
rect 14890 9078 14900 9130
rect 14924 9078 14954 9130
rect 14954 9078 14980 9130
rect 14684 9076 14740 9078
rect 14764 9076 14820 9078
rect 14844 9076 14900 9078
rect 14924 9076 14980 9078
rect 14684 8042 14740 8044
rect 14764 8042 14820 8044
rect 14844 8042 14900 8044
rect 14924 8042 14980 8044
rect 14684 7990 14710 8042
rect 14710 7990 14740 8042
rect 14764 7990 14774 8042
rect 14774 7990 14820 8042
rect 14844 7990 14890 8042
rect 14890 7990 14900 8042
rect 14924 7990 14954 8042
rect 14954 7990 14980 8042
rect 14684 7988 14740 7990
rect 14764 7988 14820 7990
rect 14844 7988 14900 7990
rect 14924 7988 14980 7990
rect 17958 21384 18014 21440
rect 18116 19466 18172 19468
rect 18196 19466 18252 19468
rect 18276 19466 18332 19468
rect 18356 19466 18412 19468
rect 18116 19414 18142 19466
rect 18142 19414 18172 19466
rect 18196 19414 18206 19466
rect 18206 19414 18252 19466
rect 18276 19414 18322 19466
rect 18322 19414 18332 19466
rect 18356 19414 18386 19466
rect 18386 19414 18412 19466
rect 18116 19412 18172 19414
rect 18196 19412 18252 19414
rect 18276 19412 18332 19414
rect 18356 19412 18412 19414
rect 18116 18378 18172 18380
rect 18196 18378 18252 18380
rect 18276 18378 18332 18380
rect 18356 18378 18412 18380
rect 18116 18326 18142 18378
rect 18142 18326 18172 18378
rect 18196 18326 18206 18378
rect 18206 18326 18252 18378
rect 18276 18326 18322 18378
rect 18322 18326 18332 18378
rect 18356 18326 18386 18378
rect 18386 18326 18412 18378
rect 18116 18324 18172 18326
rect 18196 18324 18252 18326
rect 18276 18324 18332 18326
rect 18356 18324 18412 18326
rect 18116 17290 18172 17292
rect 18196 17290 18252 17292
rect 18276 17290 18332 17292
rect 18356 17290 18412 17292
rect 18116 17238 18142 17290
rect 18142 17238 18172 17290
rect 18196 17238 18206 17290
rect 18206 17238 18252 17290
rect 18276 17238 18322 17290
rect 18322 17238 18332 17290
rect 18356 17238 18386 17290
rect 18386 17238 18412 17290
rect 18116 17236 18172 17238
rect 18196 17236 18252 17238
rect 18276 17236 18332 17238
rect 18356 17236 18412 17238
rect 18116 16202 18172 16204
rect 18196 16202 18252 16204
rect 18276 16202 18332 16204
rect 18356 16202 18412 16204
rect 18116 16150 18142 16202
rect 18142 16150 18172 16202
rect 18196 16150 18206 16202
rect 18206 16150 18252 16202
rect 18276 16150 18322 16202
rect 18322 16150 18332 16202
rect 18356 16150 18386 16202
rect 18386 16150 18412 16202
rect 18116 16148 18172 16150
rect 18196 16148 18252 16150
rect 18276 16148 18332 16150
rect 18356 16148 18412 16150
rect 18116 15114 18172 15116
rect 18196 15114 18252 15116
rect 18276 15114 18332 15116
rect 18356 15114 18412 15116
rect 18116 15062 18142 15114
rect 18142 15062 18172 15114
rect 18196 15062 18206 15114
rect 18206 15062 18252 15114
rect 18276 15062 18322 15114
rect 18322 15062 18332 15114
rect 18356 15062 18386 15114
rect 18386 15062 18412 15114
rect 18116 15060 18172 15062
rect 18196 15060 18252 15062
rect 18276 15060 18332 15062
rect 18356 15060 18412 15062
rect 18116 14026 18172 14028
rect 18196 14026 18252 14028
rect 18276 14026 18332 14028
rect 18356 14026 18412 14028
rect 18116 13974 18142 14026
rect 18142 13974 18172 14026
rect 18196 13974 18206 14026
rect 18206 13974 18252 14026
rect 18276 13974 18322 14026
rect 18322 13974 18332 14026
rect 18356 13974 18386 14026
rect 18386 13974 18412 14026
rect 18116 13972 18172 13974
rect 18196 13972 18252 13974
rect 18276 13972 18332 13974
rect 18356 13972 18412 13974
rect 18694 21928 18750 21984
rect 19246 20976 19302 21032
rect 19246 18664 19302 18720
rect 18116 12938 18172 12940
rect 18196 12938 18252 12940
rect 18276 12938 18332 12940
rect 18356 12938 18412 12940
rect 18116 12886 18142 12938
rect 18142 12886 18172 12938
rect 18196 12886 18206 12938
rect 18206 12886 18252 12938
rect 18276 12886 18322 12938
rect 18322 12886 18332 12938
rect 18356 12886 18386 12938
rect 18386 12886 18412 12938
rect 18116 12884 18172 12886
rect 18196 12884 18252 12886
rect 18276 12884 18332 12886
rect 18356 12884 18412 12886
rect 18116 11850 18172 11852
rect 18196 11850 18252 11852
rect 18276 11850 18332 11852
rect 18356 11850 18412 11852
rect 18116 11798 18142 11850
rect 18142 11798 18172 11850
rect 18196 11798 18206 11850
rect 18206 11798 18252 11850
rect 18276 11798 18322 11850
rect 18322 11798 18332 11850
rect 18356 11798 18386 11850
rect 18386 11798 18412 11850
rect 18116 11796 18172 11798
rect 18196 11796 18252 11798
rect 18276 11796 18332 11798
rect 18356 11796 18412 11798
rect 14684 6954 14740 6956
rect 14764 6954 14820 6956
rect 14844 6954 14900 6956
rect 14924 6954 14980 6956
rect 14684 6902 14710 6954
rect 14710 6902 14740 6954
rect 14764 6902 14774 6954
rect 14774 6902 14820 6954
rect 14844 6902 14890 6954
rect 14890 6902 14900 6954
rect 14924 6902 14954 6954
rect 14954 6902 14980 6954
rect 14684 6900 14740 6902
rect 14764 6900 14820 6902
rect 14844 6900 14900 6902
rect 14924 6900 14980 6902
rect 14684 5866 14740 5868
rect 14764 5866 14820 5868
rect 14844 5866 14900 5868
rect 14924 5866 14980 5868
rect 14684 5814 14710 5866
rect 14710 5814 14740 5866
rect 14764 5814 14774 5866
rect 14774 5814 14820 5866
rect 14844 5814 14890 5866
rect 14890 5814 14900 5866
rect 14924 5814 14954 5866
rect 14954 5814 14980 5866
rect 14684 5812 14740 5814
rect 14764 5812 14820 5814
rect 14844 5812 14900 5814
rect 14924 5812 14980 5814
rect 14684 4778 14740 4780
rect 14764 4778 14820 4780
rect 14844 4778 14900 4780
rect 14924 4778 14980 4780
rect 14684 4726 14710 4778
rect 14710 4726 14740 4778
rect 14764 4726 14774 4778
rect 14774 4726 14820 4778
rect 14844 4726 14890 4778
rect 14890 4726 14900 4778
rect 14924 4726 14954 4778
rect 14954 4726 14980 4778
rect 14684 4724 14740 4726
rect 14764 4724 14820 4726
rect 14844 4724 14900 4726
rect 14924 4724 14980 4726
rect 14684 3690 14740 3692
rect 14764 3690 14820 3692
rect 14844 3690 14900 3692
rect 14924 3690 14980 3692
rect 14684 3638 14710 3690
rect 14710 3638 14740 3690
rect 14764 3638 14774 3690
rect 14774 3638 14820 3690
rect 14844 3638 14890 3690
rect 14890 3638 14900 3690
rect 14924 3638 14954 3690
rect 14954 3638 14980 3690
rect 14684 3636 14740 3638
rect 14764 3636 14820 3638
rect 14844 3636 14900 3638
rect 14924 3636 14980 3638
rect 14684 2602 14740 2604
rect 14764 2602 14820 2604
rect 14844 2602 14900 2604
rect 14924 2602 14980 2604
rect 14684 2550 14710 2602
rect 14710 2550 14740 2602
rect 14764 2550 14774 2602
rect 14774 2550 14820 2602
rect 14844 2550 14890 2602
rect 14890 2550 14900 2602
rect 14924 2550 14954 2602
rect 14954 2550 14980 2602
rect 14684 2548 14740 2550
rect 14764 2548 14820 2550
rect 14844 2548 14900 2550
rect 14924 2548 14980 2550
rect 4388 2058 4444 2060
rect 4468 2058 4524 2060
rect 4548 2058 4604 2060
rect 4628 2058 4684 2060
rect 4388 2006 4414 2058
rect 4414 2006 4444 2058
rect 4468 2006 4478 2058
rect 4478 2006 4524 2058
rect 4548 2006 4594 2058
rect 4594 2006 4604 2058
rect 4628 2006 4658 2058
rect 4658 2006 4684 2058
rect 4388 2004 4444 2006
rect 4468 2004 4524 2006
rect 4548 2004 4604 2006
rect 4628 2004 4684 2006
rect 11252 2058 11308 2060
rect 11332 2058 11388 2060
rect 11412 2058 11468 2060
rect 11492 2058 11548 2060
rect 11252 2006 11278 2058
rect 11278 2006 11308 2058
rect 11332 2006 11342 2058
rect 11342 2006 11388 2058
rect 11412 2006 11458 2058
rect 11458 2006 11468 2058
rect 11492 2006 11522 2058
rect 11522 2006 11548 2058
rect 11252 2004 11308 2006
rect 11332 2004 11388 2006
rect 11412 2004 11468 2006
rect 11492 2004 11548 2006
rect 18116 10762 18172 10764
rect 18196 10762 18252 10764
rect 18276 10762 18332 10764
rect 18356 10762 18412 10764
rect 18116 10710 18142 10762
rect 18142 10710 18172 10762
rect 18196 10710 18206 10762
rect 18206 10710 18252 10762
rect 18276 10710 18322 10762
rect 18322 10710 18332 10762
rect 18356 10710 18386 10762
rect 18386 10710 18412 10762
rect 18116 10708 18172 10710
rect 18196 10708 18252 10710
rect 18276 10708 18332 10710
rect 18356 10708 18412 10710
rect 18116 9674 18172 9676
rect 18196 9674 18252 9676
rect 18276 9674 18332 9676
rect 18356 9674 18412 9676
rect 18116 9622 18142 9674
rect 18142 9622 18172 9674
rect 18196 9622 18206 9674
rect 18206 9622 18252 9674
rect 18276 9622 18322 9674
rect 18322 9622 18332 9674
rect 18356 9622 18386 9674
rect 18386 9622 18412 9674
rect 18116 9620 18172 9622
rect 18196 9620 18252 9622
rect 18276 9620 18332 9622
rect 18356 9620 18412 9622
rect 18116 8586 18172 8588
rect 18196 8586 18252 8588
rect 18276 8586 18332 8588
rect 18356 8586 18412 8588
rect 18116 8534 18142 8586
rect 18142 8534 18172 8586
rect 18196 8534 18206 8586
rect 18206 8534 18252 8586
rect 18276 8534 18322 8586
rect 18322 8534 18332 8586
rect 18356 8534 18386 8586
rect 18386 8534 18412 8586
rect 18116 8532 18172 8534
rect 18196 8532 18252 8534
rect 18276 8532 18332 8534
rect 18356 8532 18412 8534
rect 18116 7498 18172 7500
rect 18196 7498 18252 7500
rect 18276 7498 18332 7500
rect 18356 7498 18412 7500
rect 18116 7446 18142 7498
rect 18142 7446 18172 7498
rect 18196 7446 18206 7498
rect 18206 7446 18252 7498
rect 18276 7446 18322 7498
rect 18322 7446 18332 7498
rect 18356 7446 18386 7498
rect 18386 7446 18412 7498
rect 18116 7444 18172 7446
rect 18196 7444 18252 7446
rect 18276 7444 18332 7446
rect 18356 7444 18412 7446
rect 19246 12272 19302 12328
rect 18510 6424 18566 6480
rect 18116 6410 18172 6412
rect 18196 6410 18252 6412
rect 18276 6410 18332 6412
rect 18356 6410 18412 6412
rect 18116 6358 18142 6410
rect 18142 6358 18172 6410
rect 18196 6358 18206 6410
rect 18206 6358 18252 6410
rect 18276 6358 18322 6410
rect 18322 6358 18332 6410
rect 18356 6358 18386 6410
rect 18386 6358 18412 6410
rect 18116 6356 18172 6358
rect 18196 6356 18252 6358
rect 18276 6356 18332 6358
rect 18356 6356 18412 6358
rect 18602 5472 18658 5528
rect 18116 5322 18172 5324
rect 18196 5322 18252 5324
rect 18276 5322 18332 5324
rect 18356 5322 18412 5324
rect 18116 5270 18142 5322
rect 18142 5270 18172 5322
rect 18196 5270 18206 5322
rect 18206 5270 18252 5322
rect 18276 5270 18322 5322
rect 18322 5270 18332 5322
rect 18356 5270 18386 5322
rect 18386 5270 18412 5322
rect 18116 5268 18172 5270
rect 18196 5268 18252 5270
rect 18276 5268 18332 5270
rect 18356 5268 18412 5270
rect 17958 4520 18014 4576
rect 18116 4234 18172 4236
rect 18196 4234 18252 4236
rect 18276 4234 18332 4236
rect 18356 4234 18412 4236
rect 18116 4182 18142 4234
rect 18142 4182 18172 4234
rect 18196 4182 18206 4234
rect 18206 4182 18252 4234
rect 18276 4182 18322 4234
rect 18322 4182 18332 4234
rect 18356 4182 18386 4234
rect 18386 4182 18412 4234
rect 18116 4180 18172 4182
rect 18196 4180 18252 4182
rect 18276 4180 18332 4182
rect 18356 4180 18412 4182
rect 17866 3568 17922 3624
rect 18510 3160 18566 3216
rect 18116 3146 18172 3148
rect 18196 3146 18252 3148
rect 18276 3146 18332 3148
rect 18356 3146 18412 3148
rect 18116 3094 18142 3146
rect 18142 3094 18172 3146
rect 18196 3094 18206 3146
rect 18206 3094 18252 3146
rect 18276 3094 18322 3146
rect 18322 3094 18332 3146
rect 18356 3094 18386 3146
rect 18386 3094 18412 3146
rect 18116 3092 18172 3094
rect 18196 3092 18252 3094
rect 18276 3092 18332 3094
rect 18356 3092 18412 3094
rect 18116 2058 18172 2060
rect 18196 2058 18252 2060
rect 18276 2058 18332 2060
rect 18356 2058 18412 2060
rect 18116 2006 18142 2058
rect 18142 2006 18172 2058
rect 18196 2006 18206 2058
rect 18206 2006 18252 2058
rect 18276 2006 18322 2058
rect 18322 2006 18332 2058
rect 18356 2006 18386 2058
rect 18386 2006 18412 2058
rect 18116 2004 18172 2006
rect 18196 2004 18252 2006
rect 18276 2004 18332 2006
rect 18356 2004 18412 2006
rect 18602 1392 18658 1448
rect 19062 9960 19118 10016
rect 19982 19616 20038 19672
rect 19890 16896 19946 16952
rect 19890 15012 19946 15048
rect 19890 14992 19892 15012
rect 19892 14992 19944 15012
rect 19944 14992 19946 15012
rect 18970 9416 19026 9472
rect 19982 11864 20038 11920
rect 20626 20568 20682 20624
rect 20718 20024 20774 20080
rect 20442 18256 20498 18312
rect 20442 16216 20498 16272
rect 20166 14584 20222 14640
rect 20442 15944 20498 16000
rect 21270 19208 21326 19264
rect 20994 17848 21050 17904
rect 20902 15536 20958 15592
rect 20810 14176 20866 14232
rect 20166 13224 20222 13280
rect 20258 12816 20314 12872
rect 20258 10912 20314 10968
rect 19982 10504 20038 10560
rect 20258 9552 20314 9608
rect 20534 11456 20590 11512
rect 20718 13632 20774 13688
rect 20534 9144 20590 9200
rect 20534 8600 20590 8656
rect 19982 8192 20038 8248
rect 20258 7784 20314 7840
rect 20534 7240 20590 7296
rect 19982 6832 20038 6888
rect 20534 5880 20590 5936
rect 20534 4928 20590 4984
rect 21730 17324 21786 17360
rect 21730 17304 21732 17324
rect 21732 17304 21784 17324
rect 21784 17304 21786 17324
rect 20534 4112 20590 4168
rect 19246 2752 19302 2808
rect 18786 2208 18842 2264
rect 19062 848 19118 904
rect 18694 440 18750 496
rect 17314 32 17370 88
<< metal3 >>
rect 18873 22394 18939 22397
rect 22320 22394 22800 22424
rect 18873 22392 22800 22394
rect 18873 22336 18878 22392
rect 18934 22336 22800 22392
rect 18873 22334 22800 22336
rect 18873 22331 18939 22334
rect 22320 22304 22800 22334
rect 18689 21986 18755 21989
rect 22320 21986 22800 22016
rect 18689 21984 22800 21986
rect 18689 21928 18694 21984
rect 18750 21928 22800 21984
rect 18689 21926 22800 21928
rect 18689 21923 18755 21926
rect 22320 21896 22800 21926
rect 17953 21442 18019 21445
rect 22320 21442 22800 21472
rect 17953 21440 22800 21442
rect 17953 21384 17958 21440
rect 18014 21384 22800 21440
rect 17953 21382 22800 21384
rect 17953 21379 18019 21382
rect 22320 21352 22800 21382
rect 19241 21034 19307 21037
rect 22320 21034 22800 21064
rect 19241 21032 22800 21034
rect 19241 20976 19246 21032
rect 19302 20976 22800 21032
rect 19241 20974 22800 20976
rect 19241 20971 19307 20974
rect 22320 20944 22800 20974
rect 20621 20626 20687 20629
rect 22320 20626 22800 20656
rect 20621 20624 22800 20626
rect 20621 20568 20626 20624
rect 20682 20568 22800 20624
rect 20621 20566 22800 20568
rect 20621 20563 20687 20566
rect 22320 20536 22800 20566
rect 20713 20082 20779 20085
rect 22320 20082 22800 20112
rect 20713 20080 22800 20082
rect 20713 20024 20718 20080
rect 20774 20024 22800 20080
rect 20713 20022 22800 20024
rect 20713 20019 20779 20022
rect 7808 20016 8128 20017
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 19951 8128 19952
rect 14672 20016 14992 20017
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 22320 19992 22800 20022
rect 14672 19951 14992 19952
rect 19977 19674 20043 19677
rect 22320 19674 22800 19704
rect 19977 19672 22800 19674
rect 19977 19616 19982 19672
rect 20038 19616 22800 19672
rect 19977 19614 22800 19616
rect 19977 19611 20043 19614
rect 22320 19584 22800 19614
rect 4376 19472 4696 19473
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 19407 4696 19408
rect 11240 19472 11560 19473
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 19407 11560 19408
rect 18104 19472 18424 19473
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 19407 18424 19408
rect 21265 19266 21331 19269
rect 22320 19266 22800 19296
rect 21265 19264 22800 19266
rect 21265 19208 21270 19264
rect 21326 19208 22800 19264
rect 21265 19206 22800 19208
rect 21265 19203 21331 19206
rect 22320 19176 22800 19206
rect 7808 18928 8128 18929
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 18863 8128 18864
rect 14672 18928 14992 18929
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 18863 14992 18864
rect 19241 18722 19307 18725
rect 22320 18722 22800 18752
rect 19241 18720 22800 18722
rect 19241 18664 19246 18720
rect 19302 18664 22800 18720
rect 19241 18662 22800 18664
rect 19241 18659 19307 18662
rect 22320 18632 22800 18662
rect 4376 18384 4696 18385
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 18319 4696 18320
rect 11240 18384 11560 18385
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 18319 11560 18320
rect 18104 18384 18424 18385
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 18319 18424 18320
rect 20437 18314 20503 18317
rect 22320 18314 22800 18344
rect 20437 18312 22800 18314
rect 20437 18256 20442 18312
rect 20498 18256 22800 18312
rect 20437 18254 22800 18256
rect 20437 18251 20503 18254
rect 22320 18224 22800 18254
rect 20989 17906 21055 17909
rect 22320 17906 22800 17936
rect 20989 17904 22800 17906
rect 20989 17848 20994 17904
rect 21050 17848 22800 17904
rect 20989 17846 22800 17848
rect 20989 17843 21055 17846
rect 7808 17840 8128 17841
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 17775 8128 17776
rect 14672 17840 14992 17841
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 22320 17816 22800 17846
rect 14672 17775 14992 17776
rect 21725 17362 21791 17365
rect 22320 17362 22800 17392
rect 21725 17360 22800 17362
rect 21725 17304 21730 17360
rect 21786 17304 22800 17360
rect 21725 17302 22800 17304
rect 21725 17299 21791 17302
rect 4376 17296 4696 17297
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 17231 4696 17232
rect 11240 17296 11560 17297
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 17231 11560 17232
rect 18104 17296 18424 17297
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 22320 17272 22800 17302
rect 18104 17231 18424 17232
rect 0 17090 480 17120
rect 4061 17090 4127 17093
rect 0 17088 4127 17090
rect 0 17032 4066 17088
rect 4122 17032 4127 17088
rect 0 17030 4127 17032
rect 0 17000 480 17030
rect 4061 17027 4127 17030
rect 19885 16954 19951 16957
rect 22320 16954 22800 16984
rect 19885 16952 22800 16954
rect 19885 16896 19890 16952
rect 19946 16896 22800 16952
rect 19885 16894 22800 16896
rect 19885 16891 19951 16894
rect 22320 16864 22800 16894
rect 7808 16752 8128 16753
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 16687 8128 16688
rect 14672 16752 14992 16753
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 16687 14992 16688
rect 22320 16410 22800 16440
rect 20486 16350 22800 16410
rect 20486 16277 20546 16350
rect 22320 16320 22800 16350
rect 20437 16272 20546 16277
rect 20437 16216 20442 16272
rect 20498 16216 20546 16272
rect 20437 16214 20546 16216
rect 20437 16211 20503 16214
rect 4376 16208 4696 16209
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 16143 4696 16144
rect 11240 16208 11560 16209
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 16143 11560 16144
rect 18104 16208 18424 16209
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 16143 18424 16144
rect 20437 16002 20503 16005
rect 22320 16002 22800 16032
rect 20437 16000 22800 16002
rect 20437 15944 20442 16000
rect 20498 15944 22800 16000
rect 20437 15942 22800 15944
rect 20437 15939 20503 15942
rect 22320 15912 22800 15942
rect 7808 15664 8128 15665
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 15599 8128 15600
rect 14672 15664 14992 15665
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 15599 14992 15600
rect 20897 15594 20963 15597
rect 22320 15594 22800 15624
rect 20897 15592 22800 15594
rect 20897 15536 20902 15592
rect 20958 15536 22800 15592
rect 20897 15534 22800 15536
rect 20897 15531 20963 15534
rect 22320 15504 22800 15534
rect 4376 15120 4696 15121
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 15055 4696 15056
rect 11240 15120 11560 15121
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 15055 11560 15056
rect 18104 15120 18424 15121
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 15055 18424 15056
rect 19885 15050 19951 15053
rect 22320 15050 22800 15080
rect 19885 15048 22800 15050
rect 19885 14992 19890 15048
rect 19946 14992 22800 15048
rect 19885 14990 22800 14992
rect 19885 14987 19951 14990
rect 22320 14960 22800 14990
rect 20161 14642 20227 14645
rect 22320 14642 22800 14672
rect 20161 14640 22800 14642
rect 20161 14584 20166 14640
rect 20222 14584 22800 14640
rect 20161 14582 22800 14584
rect 20161 14579 20227 14582
rect 7808 14576 8128 14577
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 14511 8128 14512
rect 14672 14576 14992 14577
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 22320 14552 22800 14582
rect 14672 14511 14992 14512
rect 20805 14234 20871 14237
rect 22320 14234 22800 14264
rect 20805 14232 22800 14234
rect 20805 14176 20810 14232
rect 20866 14176 22800 14232
rect 20805 14174 22800 14176
rect 20805 14171 20871 14174
rect 22320 14144 22800 14174
rect 4376 14032 4696 14033
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 13967 4696 13968
rect 11240 14032 11560 14033
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 13967 11560 13968
rect 18104 14032 18424 14033
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 13967 18424 13968
rect 20713 13690 20779 13693
rect 22320 13690 22800 13720
rect 20713 13688 22800 13690
rect 20713 13632 20718 13688
rect 20774 13632 22800 13688
rect 20713 13630 22800 13632
rect 20713 13627 20779 13630
rect 22320 13600 22800 13630
rect 7808 13488 8128 13489
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 13423 8128 13424
rect 14672 13488 14992 13489
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 13423 14992 13424
rect 20161 13282 20227 13285
rect 22320 13282 22800 13312
rect 20161 13280 22800 13282
rect 20161 13224 20166 13280
rect 20222 13224 22800 13280
rect 20161 13222 22800 13224
rect 20161 13219 20227 13222
rect 22320 13192 22800 13222
rect 4376 12944 4696 12945
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 12879 4696 12880
rect 11240 12944 11560 12945
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 12879 11560 12880
rect 18104 12944 18424 12945
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 12879 18424 12880
rect 20253 12874 20319 12877
rect 22320 12874 22800 12904
rect 20253 12872 22800 12874
rect 20253 12816 20258 12872
rect 20314 12816 22800 12872
rect 20253 12814 22800 12816
rect 20253 12811 20319 12814
rect 22320 12784 22800 12814
rect 7808 12400 8128 12401
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 12335 8128 12336
rect 14672 12400 14992 12401
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 12335 14992 12336
rect 19241 12330 19307 12333
rect 22320 12330 22800 12360
rect 19241 12328 22800 12330
rect 19241 12272 19246 12328
rect 19302 12272 22800 12328
rect 19241 12270 22800 12272
rect 19241 12267 19307 12270
rect 22320 12240 22800 12270
rect 19977 11922 20043 11925
rect 22320 11922 22800 11952
rect 19977 11920 22800 11922
rect 19977 11864 19982 11920
rect 20038 11864 22800 11920
rect 19977 11862 22800 11864
rect 19977 11859 20043 11862
rect 4376 11856 4696 11857
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 11791 4696 11792
rect 11240 11856 11560 11857
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 11791 11560 11792
rect 18104 11856 18424 11857
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 22320 11832 22800 11862
rect 18104 11791 18424 11792
rect 20529 11514 20595 11517
rect 22320 11514 22800 11544
rect 20529 11512 22800 11514
rect 20529 11456 20534 11512
rect 20590 11456 22800 11512
rect 20529 11454 22800 11456
rect 20529 11451 20595 11454
rect 22320 11424 22800 11454
rect 7808 11312 8128 11313
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 11247 8128 11248
rect 14672 11312 14992 11313
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 11247 14992 11248
rect 20253 10970 20319 10973
rect 22320 10970 22800 11000
rect 20253 10968 22800 10970
rect 20253 10912 20258 10968
rect 20314 10912 22800 10968
rect 20253 10910 22800 10912
rect 20253 10907 20319 10910
rect 22320 10880 22800 10910
rect 4376 10768 4696 10769
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 10703 4696 10704
rect 11240 10768 11560 10769
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 10703 11560 10704
rect 18104 10768 18424 10769
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 10703 18424 10704
rect 19977 10562 20043 10565
rect 22320 10562 22800 10592
rect 19977 10560 22800 10562
rect 19977 10504 19982 10560
rect 20038 10504 22800 10560
rect 19977 10502 22800 10504
rect 19977 10499 20043 10502
rect 22320 10472 22800 10502
rect 7808 10224 8128 10225
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 10159 8128 10160
rect 14672 10224 14992 10225
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 10159 14992 10160
rect 19057 10018 19123 10021
rect 22320 10018 22800 10048
rect 19057 10016 22800 10018
rect 19057 9960 19062 10016
rect 19118 9960 22800 10016
rect 19057 9958 22800 9960
rect 19057 9955 19123 9958
rect 22320 9928 22800 9958
rect 4376 9680 4696 9681
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 9615 4696 9616
rect 11240 9680 11560 9681
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 9615 11560 9616
rect 18104 9680 18424 9681
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 9615 18424 9616
rect 20253 9610 20319 9613
rect 22320 9610 22800 9640
rect 20253 9608 22800 9610
rect 20253 9552 20258 9608
rect 20314 9552 22800 9608
rect 20253 9550 22800 9552
rect 20253 9547 20319 9550
rect 22320 9520 22800 9550
rect 18822 9412 18828 9476
rect 18892 9474 18898 9476
rect 18965 9474 19031 9477
rect 18892 9472 19031 9474
rect 18892 9416 18970 9472
rect 19026 9416 19031 9472
rect 18892 9414 19031 9416
rect 18892 9412 18898 9414
rect 18965 9411 19031 9414
rect 20529 9202 20595 9205
rect 22320 9202 22800 9232
rect 20529 9200 22800 9202
rect 20529 9144 20534 9200
rect 20590 9144 22800 9200
rect 20529 9142 22800 9144
rect 20529 9139 20595 9142
rect 7808 9136 8128 9137
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 9071 8128 9072
rect 14672 9136 14992 9137
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 22320 9112 22800 9142
rect 14672 9071 14992 9072
rect 20529 8658 20595 8661
rect 22320 8658 22800 8688
rect 20529 8656 22800 8658
rect 20529 8600 20534 8656
rect 20590 8600 22800 8656
rect 20529 8598 22800 8600
rect 20529 8595 20595 8598
rect 4376 8592 4696 8593
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 8527 4696 8528
rect 11240 8592 11560 8593
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 8527 11560 8528
rect 18104 8592 18424 8593
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 22320 8568 22800 8598
rect 18104 8527 18424 8528
rect 19977 8250 20043 8253
rect 22320 8250 22800 8280
rect 19977 8248 22800 8250
rect 19977 8192 19982 8248
rect 20038 8192 22800 8248
rect 19977 8190 22800 8192
rect 19977 8187 20043 8190
rect 22320 8160 22800 8190
rect 7808 8048 8128 8049
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 7983 8128 7984
rect 14672 8048 14992 8049
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 7983 14992 7984
rect 20253 7842 20319 7845
rect 22320 7842 22800 7872
rect 20253 7840 22800 7842
rect 20253 7784 20258 7840
rect 20314 7784 22800 7840
rect 20253 7782 22800 7784
rect 20253 7779 20319 7782
rect 22320 7752 22800 7782
rect 4376 7504 4696 7505
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 7439 4696 7440
rect 11240 7504 11560 7505
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 7439 11560 7440
rect 18104 7504 18424 7505
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 7439 18424 7440
rect 20529 7298 20595 7301
rect 22320 7298 22800 7328
rect 20529 7296 22800 7298
rect 20529 7240 20534 7296
rect 20590 7240 22800 7296
rect 20529 7238 22800 7240
rect 20529 7235 20595 7238
rect 22320 7208 22800 7238
rect 7808 6960 8128 6961
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 6895 8128 6896
rect 14672 6960 14992 6961
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 6895 14992 6896
rect 19977 6890 20043 6893
rect 22320 6890 22800 6920
rect 19977 6888 22800 6890
rect 19977 6832 19982 6888
rect 20038 6832 22800 6888
rect 19977 6830 22800 6832
rect 19977 6827 20043 6830
rect 22320 6800 22800 6830
rect 18505 6482 18571 6485
rect 22320 6482 22800 6512
rect 18505 6480 22800 6482
rect 18505 6424 18510 6480
rect 18566 6424 22800 6480
rect 18505 6422 22800 6424
rect 18505 6419 18571 6422
rect 4376 6416 4696 6417
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 6351 4696 6352
rect 11240 6416 11560 6417
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 6351 11560 6352
rect 18104 6416 18424 6417
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 22320 6392 22800 6422
rect 18104 6351 18424 6352
rect 20529 5938 20595 5941
rect 22320 5938 22800 5968
rect 20529 5936 22800 5938
rect 20529 5880 20534 5936
rect 20590 5880 22800 5936
rect 20529 5878 22800 5880
rect 20529 5875 20595 5878
rect 7808 5872 8128 5873
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 5807 8128 5808
rect 14672 5872 14992 5873
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 22320 5848 22800 5878
rect 14672 5807 14992 5808
rect 0 5666 480 5696
rect 4061 5666 4127 5669
rect 0 5664 4127 5666
rect 0 5608 4066 5664
rect 4122 5608 4127 5664
rect 0 5606 4127 5608
rect 0 5576 480 5606
rect 4061 5603 4127 5606
rect 18597 5530 18663 5533
rect 22320 5530 22800 5560
rect 18597 5528 22800 5530
rect 18597 5472 18602 5528
rect 18658 5472 22800 5528
rect 18597 5470 22800 5472
rect 18597 5467 18663 5470
rect 22320 5440 22800 5470
rect 4376 5328 4696 5329
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 5263 4696 5264
rect 11240 5328 11560 5329
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 5263 11560 5264
rect 18104 5328 18424 5329
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 5263 18424 5264
rect 20529 4986 20595 4989
rect 22320 4986 22800 5016
rect 20529 4984 22800 4986
rect 20529 4928 20534 4984
rect 20590 4928 22800 4984
rect 20529 4926 22800 4928
rect 20529 4923 20595 4926
rect 22320 4896 22800 4926
rect 7808 4784 8128 4785
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 4719 8128 4720
rect 14672 4784 14992 4785
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 4719 14992 4720
rect 17953 4578 18019 4581
rect 22320 4578 22800 4608
rect 17953 4576 22800 4578
rect 17953 4520 17958 4576
rect 18014 4520 22800 4576
rect 17953 4518 22800 4520
rect 17953 4515 18019 4518
rect 22320 4488 22800 4518
rect 4376 4240 4696 4241
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 4175 4696 4176
rect 11240 4240 11560 4241
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 4175 11560 4176
rect 18104 4240 18424 4241
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 4175 18424 4176
rect 20529 4170 20595 4173
rect 22320 4170 22800 4200
rect 20529 4168 22800 4170
rect 20529 4112 20534 4168
rect 20590 4112 22800 4168
rect 20529 4110 22800 4112
rect 20529 4107 20595 4110
rect 22320 4080 22800 4110
rect 7808 3696 8128 3697
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 3631 8128 3632
rect 14672 3696 14992 3697
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 3631 14992 3632
rect 17861 3626 17927 3629
rect 22320 3626 22800 3656
rect 17861 3624 22800 3626
rect 17861 3568 17866 3624
rect 17922 3568 22800 3624
rect 17861 3566 22800 3568
rect 17861 3563 17927 3566
rect 22320 3536 22800 3566
rect 18505 3218 18571 3221
rect 22320 3218 22800 3248
rect 18505 3216 22800 3218
rect 18505 3160 18510 3216
rect 18566 3160 22800 3216
rect 18505 3158 22800 3160
rect 18505 3155 18571 3158
rect 4376 3152 4696 3153
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 3087 4696 3088
rect 11240 3152 11560 3153
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 3087 11560 3088
rect 18104 3152 18424 3153
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 22320 3128 22800 3158
rect 18104 3087 18424 3088
rect 19241 2810 19307 2813
rect 22320 2810 22800 2840
rect 19241 2808 22800 2810
rect 19241 2752 19246 2808
rect 19302 2752 22800 2808
rect 19241 2750 22800 2752
rect 19241 2747 19307 2750
rect 22320 2720 22800 2750
rect 7808 2608 8128 2609
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 2543 8128 2544
rect 14672 2608 14992 2609
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 2543 14992 2544
rect 18781 2266 18847 2269
rect 22320 2266 22800 2296
rect 18781 2264 22800 2266
rect 18781 2208 18786 2264
rect 18842 2208 22800 2264
rect 18781 2206 22800 2208
rect 18781 2203 18847 2206
rect 22320 2176 22800 2206
rect 4376 2064 4696 2065
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1999 4696 2000
rect 11240 2064 11560 2065
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1999 11560 2000
rect 18104 2064 18424 2065
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1999 18424 2000
rect 18822 1796 18828 1860
rect 18892 1858 18898 1860
rect 22320 1858 22800 1888
rect 18892 1798 22800 1858
rect 18892 1796 18898 1798
rect 22320 1768 22800 1798
rect 18597 1450 18663 1453
rect 22320 1450 22800 1480
rect 18597 1448 22800 1450
rect 18597 1392 18602 1448
rect 18658 1392 22800 1448
rect 18597 1390 22800 1392
rect 18597 1387 18663 1390
rect 22320 1360 22800 1390
rect 19057 906 19123 909
rect 22320 906 22800 936
rect 19057 904 22800 906
rect 19057 848 19062 904
rect 19118 848 22800 904
rect 19057 846 22800 848
rect 19057 843 19123 846
rect 22320 816 22800 846
rect 18689 498 18755 501
rect 22320 498 22800 528
rect 18689 496 22800 498
rect 18689 440 18694 496
rect 18750 440 22800 496
rect 18689 438 22800 440
rect 18689 435 18755 438
rect 22320 408 22800 438
rect 17309 90 17375 93
rect 22320 90 22800 120
rect 17309 88 22800 90
rect 17309 32 17314 88
rect 17370 32 22800 88
rect 17309 30 22800 32
rect 17309 27 17375 30
rect 22320 0 22800 30
<< via3 >>
rect 7816 20012 7880 20016
rect 7816 19956 7820 20012
rect 7820 19956 7876 20012
rect 7876 19956 7880 20012
rect 7816 19952 7880 19956
rect 7896 20012 7960 20016
rect 7896 19956 7900 20012
rect 7900 19956 7956 20012
rect 7956 19956 7960 20012
rect 7896 19952 7960 19956
rect 7976 20012 8040 20016
rect 7976 19956 7980 20012
rect 7980 19956 8036 20012
rect 8036 19956 8040 20012
rect 7976 19952 8040 19956
rect 8056 20012 8120 20016
rect 8056 19956 8060 20012
rect 8060 19956 8116 20012
rect 8116 19956 8120 20012
rect 8056 19952 8120 19956
rect 14680 20012 14744 20016
rect 14680 19956 14684 20012
rect 14684 19956 14740 20012
rect 14740 19956 14744 20012
rect 14680 19952 14744 19956
rect 14760 20012 14824 20016
rect 14760 19956 14764 20012
rect 14764 19956 14820 20012
rect 14820 19956 14824 20012
rect 14760 19952 14824 19956
rect 14840 20012 14904 20016
rect 14840 19956 14844 20012
rect 14844 19956 14900 20012
rect 14900 19956 14904 20012
rect 14840 19952 14904 19956
rect 14920 20012 14984 20016
rect 14920 19956 14924 20012
rect 14924 19956 14980 20012
rect 14980 19956 14984 20012
rect 14920 19952 14984 19956
rect 4384 19468 4448 19472
rect 4384 19412 4388 19468
rect 4388 19412 4444 19468
rect 4444 19412 4448 19468
rect 4384 19408 4448 19412
rect 4464 19468 4528 19472
rect 4464 19412 4468 19468
rect 4468 19412 4524 19468
rect 4524 19412 4528 19468
rect 4464 19408 4528 19412
rect 4544 19468 4608 19472
rect 4544 19412 4548 19468
rect 4548 19412 4604 19468
rect 4604 19412 4608 19468
rect 4544 19408 4608 19412
rect 4624 19468 4688 19472
rect 4624 19412 4628 19468
rect 4628 19412 4684 19468
rect 4684 19412 4688 19468
rect 4624 19408 4688 19412
rect 11248 19468 11312 19472
rect 11248 19412 11252 19468
rect 11252 19412 11308 19468
rect 11308 19412 11312 19468
rect 11248 19408 11312 19412
rect 11328 19468 11392 19472
rect 11328 19412 11332 19468
rect 11332 19412 11388 19468
rect 11388 19412 11392 19468
rect 11328 19408 11392 19412
rect 11408 19468 11472 19472
rect 11408 19412 11412 19468
rect 11412 19412 11468 19468
rect 11468 19412 11472 19468
rect 11408 19408 11472 19412
rect 11488 19468 11552 19472
rect 11488 19412 11492 19468
rect 11492 19412 11548 19468
rect 11548 19412 11552 19468
rect 11488 19408 11552 19412
rect 18112 19468 18176 19472
rect 18112 19412 18116 19468
rect 18116 19412 18172 19468
rect 18172 19412 18176 19468
rect 18112 19408 18176 19412
rect 18192 19468 18256 19472
rect 18192 19412 18196 19468
rect 18196 19412 18252 19468
rect 18252 19412 18256 19468
rect 18192 19408 18256 19412
rect 18272 19468 18336 19472
rect 18272 19412 18276 19468
rect 18276 19412 18332 19468
rect 18332 19412 18336 19468
rect 18272 19408 18336 19412
rect 18352 19468 18416 19472
rect 18352 19412 18356 19468
rect 18356 19412 18412 19468
rect 18412 19412 18416 19468
rect 18352 19408 18416 19412
rect 7816 18924 7880 18928
rect 7816 18868 7820 18924
rect 7820 18868 7876 18924
rect 7876 18868 7880 18924
rect 7816 18864 7880 18868
rect 7896 18924 7960 18928
rect 7896 18868 7900 18924
rect 7900 18868 7956 18924
rect 7956 18868 7960 18924
rect 7896 18864 7960 18868
rect 7976 18924 8040 18928
rect 7976 18868 7980 18924
rect 7980 18868 8036 18924
rect 8036 18868 8040 18924
rect 7976 18864 8040 18868
rect 8056 18924 8120 18928
rect 8056 18868 8060 18924
rect 8060 18868 8116 18924
rect 8116 18868 8120 18924
rect 8056 18864 8120 18868
rect 14680 18924 14744 18928
rect 14680 18868 14684 18924
rect 14684 18868 14740 18924
rect 14740 18868 14744 18924
rect 14680 18864 14744 18868
rect 14760 18924 14824 18928
rect 14760 18868 14764 18924
rect 14764 18868 14820 18924
rect 14820 18868 14824 18924
rect 14760 18864 14824 18868
rect 14840 18924 14904 18928
rect 14840 18868 14844 18924
rect 14844 18868 14900 18924
rect 14900 18868 14904 18924
rect 14840 18864 14904 18868
rect 14920 18924 14984 18928
rect 14920 18868 14924 18924
rect 14924 18868 14980 18924
rect 14980 18868 14984 18924
rect 14920 18864 14984 18868
rect 4384 18380 4448 18384
rect 4384 18324 4388 18380
rect 4388 18324 4444 18380
rect 4444 18324 4448 18380
rect 4384 18320 4448 18324
rect 4464 18380 4528 18384
rect 4464 18324 4468 18380
rect 4468 18324 4524 18380
rect 4524 18324 4528 18380
rect 4464 18320 4528 18324
rect 4544 18380 4608 18384
rect 4544 18324 4548 18380
rect 4548 18324 4604 18380
rect 4604 18324 4608 18380
rect 4544 18320 4608 18324
rect 4624 18380 4688 18384
rect 4624 18324 4628 18380
rect 4628 18324 4684 18380
rect 4684 18324 4688 18380
rect 4624 18320 4688 18324
rect 11248 18380 11312 18384
rect 11248 18324 11252 18380
rect 11252 18324 11308 18380
rect 11308 18324 11312 18380
rect 11248 18320 11312 18324
rect 11328 18380 11392 18384
rect 11328 18324 11332 18380
rect 11332 18324 11388 18380
rect 11388 18324 11392 18380
rect 11328 18320 11392 18324
rect 11408 18380 11472 18384
rect 11408 18324 11412 18380
rect 11412 18324 11468 18380
rect 11468 18324 11472 18380
rect 11408 18320 11472 18324
rect 11488 18380 11552 18384
rect 11488 18324 11492 18380
rect 11492 18324 11548 18380
rect 11548 18324 11552 18380
rect 11488 18320 11552 18324
rect 18112 18380 18176 18384
rect 18112 18324 18116 18380
rect 18116 18324 18172 18380
rect 18172 18324 18176 18380
rect 18112 18320 18176 18324
rect 18192 18380 18256 18384
rect 18192 18324 18196 18380
rect 18196 18324 18252 18380
rect 18252 18324 18256 18380
rect 18192 18320 18256 18324
rect 18272 18380 18336 18384
rect 18272 18324 18276 18380
rect 18276 18324 18332 18380
rect 18332 18324 18336 18380
rect 18272 18320 18336 18324
rect 18352 18380 18416 18384
rect 18352 18324 18356 18380
rect 18356 18324 18412 18380
rect 18412 18324 18416 18380
rect 18352 18320 18416 18324
rect 7816 17836 7880 17840
rect 7816 17780 7820 17836
rect 7820 17780 7876 17836
rect 7876 17780 7880 17836
rect 7816 17776 7880 17780
rect 7896 17836 7960 17840
rect 7896 17780 7900 17836
rect 7900 17780 7956 17836
rect 7956 17780 7960 17836
rect 7896 17776 7960 17780
rect 7976 17836 8040 17840
rect 7976 17780 7980 17836
rect 7980 17780 8036 17836
rect 8036 17780 8040 17836
rect 7976 17776 8040 17780
rect 8056 17836 8120 17840
rect 8056 17780 8060 17836
rect 8060 17780 8116 17836
rect 8116 17780 8120 17836
rect 8056 17776 8120 17780
rect 14680 17836 14744 17840
rect 14680 17780 14684 17836
rect 14684 17780 14740 17836
rect 14740 17780 14744 17836
rect 14680 17776 14744 17780
rect 14760 17836 14824 17840
rect 14760 17780 14764 17836
rect 14764 17780 14820 17836
rect 14820 17780 14824 17836
rect 14760 17776 14824 17780
rect 14840 17836 14904 17840
rect 14840 17780 14844 17836
rect 14844 17780 14900 17836
rect 14900 17780 14904 17836
rect 14840 17776 14904 17780
rect 14920 17836 14984 17840
rect 14920 17780 14924 17836
rect 14924 17780 14980 17836
rect 14980 17780 14984 17836
rect 14920 17776 14984 17780
rect 4384 17292 4448 17296
rect 4384 17236 4388 17292
rect 4388 17236 4444 17292
rect 4444 17236 4448 17292
rect 4384 17232 4448 17236
rect 4464 17292 4528 17296
rect 4464 17236 4468 17292
rect 4468 17236 4524 17292
rect 4524 17236 4528 17292
rect 4464 17232 4528 17236
rect 4544 17292 4608 17296
rect 4544 17236 4548 17292
rect 4548 17236 4604 17292
rect 4604 17236 4608 17292
rect 4544 17232 4608 17236
rect 4624 17292 4688 17296
rect 4624 17236 4628 17292
rect 4628 17236 4684 17292
rect 4684 17236 4688 17292
rect 4624 17232 4688 17236
rect 11248 17292 11312 17296
rect 11248 17236 11252 17292
rect 11252 17236 11308 17292
rect 11308 17236 11312 17292
rect 11248 17232 11312 17236
rect 11328 17292 11392 17296
rect 11328 17236 11332 17292
rect 11332 17236 11388 17292
rect 11388 17236 11392 17292
rect 11328 17232 11392 17236
rect 11408 17292 11472 17296
rect 11408 17236 11412 17292
rect 11412 17236 11468 17292
rect 11468 17236 11472 17292
rect 11408 17232 11472 17236
rect 11488 17292 11552 17296
rect 11488 17236 11492 17292
rect 11492 17236 11548 17292
rect 11548 17236 11552 17292
rect 11488 17232 11552 17236
rect 18112 17292 18176 17296
rect 18112 17236 18116 17292
rect 18116 17236 18172 17292
rect 18172 17236 18176 17292
rect 18112 17232 18176 17236
rect 18192 17292 18256 17296
rect 18192 17236 18196 17292
rect 18196 17236 18252 17292
rect 18252 17236 18256 17292
rect 18192 17232 18256 17236
rect 18272 17292 18336 17296
rect 18272 17236 18276 17292
rect 18276 17236 18332 17292
rect 18332 17236 18336 17292
rect 18272 17232 18336 17236
rect 18352 17292 18416 17296
rect 18352 17236 18356 17292
rect 18356 17236 18412 17292
rect 18412 17236 18416 17292
rect 18352 17232 18416 17236
rect 7816 16748 7880 16752
rect 7816 16692 7820 16748
rect 7820 16692 7876 16748
rect 7876 16692 7880 16748
rect 7816 16688 7880 16692
rect 7896 16748 7960 16752
rect 7896 16692 7900 16748
rect 7900 16692 7956 16748
rect 7956 16692 7960 16748
rect 7896 16688 7960 16692
rect 7976 16748 8040 16752
rect 7976 16692 7980 16748
rect 7980 16692 8036 16748
rect 8036 16692 8040 16748
rect 7976 16688 8040 16692
rect 8056 16748 8120 16752
rect 8056 16692 8060 16748
rect 8060 16692 8116 16748
rect 8116 16692 8120 16748
rect 8056 16688 8120 16692
rect 14680 16748 14744 16752
rect 14680 16692 14684 16748
rect 14684 16692 14740 16748
rect 14740 16692 14744 16748
rect 14680 16688 14744 16692
rect 14760 16748 14824 16752
rect 14760 16692 14764 16748
rect 14764 16692 14820 16748
rect 14820 16692 14824 16748
rect 14760 16688 14824 16692
rect 14840 16748 14904 16752
rect 14840 16692 14844 16748
rect 14844 16692 14900 16748
rect 14900 16692 14904 16748
rect 14840 16688 14904 16692
rect 14920 16748 14984 16752
rect 14920 16692 14924 16748
rect 14924 16692 14980 16748
rect 14980 16692 14984 16748
rect 14920 16688 14984 16692
rect 4384 16204 4448 16208
rect 4384 16148 4388 16204
rect 4388 16148 4444 16204
rect 4444 16148 4448 16204
rect 4384 16144 4448 16148
rect 4464 16204 4528 16208
rect 4464 16148 4468 16204
rect 4468 16148 4524 16204
rect 4524 16148 4528 16204
rect 4464 16144 4528 16148
rect 4544 16204 4608 16208
rect 4544 16148 4548 16204
rect 4548 16148 4604 16204
rect 4604 16148 4608 16204
rect 4544 16144 4608 16148
rect 4624 16204 4688 16208
rect 4624 16148 4628 16204
rect 4628 16148 4684 16204
rect 4684 16148 4688 16204
rect 4624 16144 4688 16148
rect 11248 16204 11312 16208
rect 11248 16148 11252 16204
rect 11252 16148 11308 16204
rect 11308 16148 11312 16204
rect 11248 16144 11312 16148
rect 11328 16204 11392 16208
rect 11328 16148 11332 16204
rect 11332 16148 11388 16204
rect 11388 16148 11392 16204
rect 11328 16144 11392 16148
rect 11408 16204 11472 16208
rect 11408 16148 11412 16204
rect 11412 16148 11468 16204
rect 11468 16148 11472 16204
rect 11408 16144 11472 16148
rect 11488 16204 11552 16208
rect 11488 16148 11492 16204
rect 11492 16148 11548 16204
rect 11548 16148 11552 16204
rect 11488 16144 11552 16148
rect 18112 16204 18176 16208
rect 18112 16148 18116 16204
rect 18116 16148 18172 16204
rect 18172 16148 18176 16204
rect 18112 16144 18176 16148
rect 18192 16204 18256 16208
rect 18192 16148 18196 16204
rect 18196 16148 18252 16204
rect 18252 16148 18256 16204
rect 18192 16144 18256 16148
rect 18272 16204 18336 16208
rect 18272 16148 18276 16204
rect 18276 16148 18332 16204
rect 18332 16148 18336 16204
rect 18272 16144 18336 16148
rect 18352 16204 18416 16208
rect 18352 16148 18356 16204
rect 18356 16148 18412 16204
rect 18412 16148 18416 16204
rect 18352 16144 18416 16148
rect 7816 15660 7880 15664
rect 7816 15604 7820 15660
rect 7820 15604 7876 15660
rect 7876 15604 7880 15660
rect 7816 15600 7880 15604
rect 7896 15660 7960 15664
rect 7896 15604 7900 15660
rect 7900 15604 7956 15660
rect 7956 15604 7960 15660
rect 7896 15600 7960 15604
rect 7976 15660 8040 15664
rect 7976 15604 7980 15660
rect 7980 15604 8036 15660
rect 8036 15604 8040 15660
rect 7976 15600 8040 15604
rect 8056 15660 8120 15664
rect 8056 15604 8060 15660
rect 8060 15604 8116 15660
rect 8116 15604 8120 15660
rect 8056 15600 8120 15604
rect 14680 15660 14744 15664
rect 14680 15604 14684 15660
rect 14684 15604 14740 15660
rect 14740 15604 14744 15660
rect 14680 15600 14744 15604
rect 14760 15660 14824 15664
rect 14760 15604 14764 15660
rect 14764 15604 14820 15660
rect 14820 15604 14824 15660
rect 14760 15600 14824 15604
rect 14840 15660 14904 15664
rect 14840 15604 14844 15660
rect 14844 15604 14900 15660
rect 14900 15604 14904 15660
rect 14840 15600 14904 15604
rect 14920 15660 14984 15664
rect 14920 15604 14924 15660
rect 14924 15604 14980 15660
rect 14980 15604 14984 15660
rect 14920 15600 14984 15604
rect 4384 15116 4448 15120
rect 4384 15060 4388 15116
rect 4388 15060 4444 15116
rect 4444 15060 4448 15116
rect 4384 15056 4448 15060
rect 4464 15116 4528 15120
rect 4464 15060 4468 15116
rect 4468 15060 4524 15116
rect 4524 15060 4528 15116
rect 4464 15056 4528 15060
rect 4544 15116 4608 15120
rect 4544 15060 4548 15116
rect 4548 15060 4604 15116
rect 4604 15060 4608 15116
rect 4544 15056 4608 15060
rect 4624 15116 4688 15120
rect 4624 15060 4628 15116
rect 4628 15060 4684 15116
rect 4684 15060 4688 15116
rect 4624 15056 4688 15060
rect 11248 15116 11312 15120
rect 11248 15060 11252 15116
rect 11252 15060 11308 15116
rect 11308 15060 11312 15116
rect 11248 15056 11312 15060
rect 11328 15116 11392 15120
rect 11328 15060 11332 15116
rect 11332 15060 11388 15116
rect 11388 15060 11392 15116
rect 11328 15056 11392 15060
rect 11408 15116 11472 15120
rect 11408 15060 11412 15116
rect 11412 15060 11468 15116
rect 11468 15060 11472 15116
rect 11408 15056 11472 15060
rect 11488 15116 11552 15120
rect 11488 15060 11492 15116
rect 11492 15060 11548 15116
rect 11548 15060 11552 15116
rect 11488 15056 11552 15060
rect 18112 15116 18176 15120
rect 18112 15060 18116 15116
rect 18116 15060 18172 15116
rect 18172 15060 18176 15116
rect 18112 15056 18176 15060
rect 18192 15116 18256 15120
rect 18192 15060 18196 15116
rect 18196 15060 18252 15116
rect 18252 15060 18256 15116
rect 18192 15056 18256 15060
rect 18272 15116 18336 15120
rect 18272 15060 18276 15116
rect 18276 15060 18332 15116
rect 18332 15060 18336 15116
rect 18272 15056 18336 15060
rect 18352 15116 18416 15120
rect 18352 15060 18356 15116
rect 18356 15060 18412 15116
rect 18412 15060 18416 15116
rect 18352 15056 18416 15060
rect 7816 14572 7880 14576
rect 7816 14516 7820 14572
rect 7820 14516 7876 14572
rect 7876 14516 7880 14572
rect 7816 14512 7880 14516
rect 7896 14572 7960 14576
rect 7896 14516 7900 14572
rect 7900 14516 7956 14572
rect 7956 14516 7960 14572
rect 7896 14512 7960 14516
rect 7976 14572 8040 14576
rect 7976 14516 7980 14572
rect 7980 14516 8036 14572
rect 8036 14516 8040 14572
rect 7976 14512 8040 14516
rect 8056 14572 8120 14576
rect 8056 14516 8060 14572
rect 8060 14516 8116 14572
rect 8116 14516 8120 14572
rect 8056 14512 8120 14516
rect 14680 14572 14744 14576
rect 14680 14516 14684 14572
rect 14684 14516 14740 14572
rect 14740 14516 14744 14572
rect 14680 14512 14744 14516
rect 14760 14572 14824 14576
rect 14760 14516 14764 14572
rect 14764 14516 14820 14572
rect 14820 14516 14824 14572
rect 14760 14512 14824 14516
rect 14840 14572 14904 14576
rect 14840 14516 14844 14572
rect 14844 14516 14900 14572
rect 14900 14516 14904 14572
rect 14840 14512 14904 14516
rect 14920 14572 14984 14576
rect 14920 14516 14924 14572
rect 14924 14516 14980 14572
rect 14980 14516 14984 14572
rect 14920 14512 14984 14516
rect 4384 14028 4448 14032
rect 4384 13972 4388 14028
rect 4388 13972 4444 14028
rect 4444 13972 4448 14028
rect 4384 13968 4448 13972
rect 4464 14028 4528 14032
rect 4464 13972 4468 14028
rect 4468 13972 4524 14028
rect 4524 13972 4528 14028
rect 4464 13968 4528 13972
rect 4544 14028 4608 14032
rect 4544 13972 4548 14028
rect 4548 13972 4604 14028
rect 4604 13972 4608 14028
rect 4544 13968 4608 13972
rect 4624 14028 4688 14032
rect 4624 13972 4628 14028
rect 4628 13972 4684 14028
rect 4684 13972 4688 14028
rect 4624 13968 4688 13972
rect 11248 14028 11312 14032
rect 11248 13972 11252 14028
rect 11252 13972 11308 14028
rect 11308 13972 11312 14028
rect 11248 13968 11312 13972
rect 11328 14028 11392 14032
rect 11328 13972 11332 14028
rect 11332 13972 11388 14028
rect 11388 13972 11392 14028
rect 11328 13968 11392 13972
rect 11408 14028 11472 14032
rect 11408 13972 11412 14028
rect 11412 13972 11468 14028
rect 11468 13972 11472 14028
rect 11408 13968 11472 13972
rect 11488 14028 11552 14032
rect 11488 13972 11492 14028
rect 11492 13972 11548 14028
rect 11548 13972 11552 14028
rect 11488 13968 11552 13972
rect 18112 14028 18176 14032
rect 18112 13972 18116 14028
rect 18116 13972 18172 14028
rect 18172 13972 18176 14028
rect 18112 13968 18176 13972
rect 18192 14028 18256 14032
rect 18192 13972 18196 14028
rect 18196 13972 18252 14028
rect 18252 13972 18256 14028
rect 18192 13968 18256 13972
rect 18272 14028 18336 14032
rect 18272 13972 18276 14028
rect 18276 13972 18332 14028
rect 18332 13972 18336 14028
rect 18272 13968 18336 13972
rect 18352 14028 18416 14032
rect 18352 13972 18356 14028
rect 18356 13972 18412 14028
rect 18412 13972 18416 14028
rect 18352 13968 18416 13972
rect 7816 13484 7880 13488
rect 7816 13428 7820 13484
rect 7820 13428 7876 13484
rect 7876 13428 7880 13484
rect 7816 13424 7880 13428
rect 7896 13484 7960 13488
rect 7896 13428 7900 13484
rect 7900 13428 7956 13484
rect 7956 13428 7960 13484
rect 7896 13424 7960 13428
rect 7976 13484 8040 13488
rect 7976 13428 7980 13484
rect 7980 13428 8036 13484
rect 8036 13428 8040 13484
rect 7976 13424 8040 13428
rect 8056 13484 8120 13488
rect 8056 13428 8060 13484
rect 8060 13428 8116 13484
rect 8116 13428 8120 13484
rect 8056 13424 8120 13428
rect 14680 13484 14744 13488
rect 14680 13428 14684 13484
rect 14684 13428 14740 13484
rect 14740 13428 14744 13484
rect 14680 13424 14744 13428
rect 14760 13484 14824 13488
rect 14760 13428 14764 13484
rect 14764 13428 14820 13484
rect 14820 13428 14824 13484
rect 14760 13424 14824 13428
rect 14840 13484 14904 13488
rect 14840 13428 14844 13484
rect 14844 13428 14900 13484
rect 14900 13428 14904 13484
rect 14840 13424 14904 13428
rect 14920 13484 14984 13488
rect 14920 13428 14924 13484
rect 14924 13428 14980 13484
rect 14980 13428 14984 13484
rect 14920 13424 14984 13428
rect 4384 12940 4448 12944
rect 4384 12884 4388 12940
rect 4388 12884 4444 12940
rect 4444 12884 4448 12940
rect 4384 12880 4448 12884
rect 4464 12940 4528 12944
rect 4464 12884 4468 12940
rect 4468 12884 4524 12940
rect 4524 12884 4528 12940
rect 4464 12880 4528 12884
rect 4544 12940 4608 12944
rect 4544 12884 4548 12940
rect 4548 12884 4604 12940
rect 4604 12884 4608 12940
rect 4544 12880 4608 12884
rect 4624 12940 4688 12944
rect 4624 12884 4628 12940
rect 4628 12884 4684 12940
rect 4684 12884 4688 12940
rect 4624 12880 4688 12884
rect 11248 12940 11312 12944
rect 11248 12884 11252 12940
rect 11252 12884 11308 12940
rect 11308 12884 11312 12940
rect 11248 12880 11312 12884
rect 11328 12940 11392 12944
rect 11328 12884 11332 12940
rect 11332 12884 11388 12940
rect 11388 12884 11392 12940
rect 11328 12880 11392 12884
rect 11408 12940 11472 12944
rect 11408 12884 11412 12940
rect 11412 12884 11468 12940
rect 11468 12884 11472 12940
rect 11408 12880 11472 12884
rect 11488 12940 11552 12944
rect 11488 12884 11492 12940
rect 11492 12884 11548 12940
rect 11548 12884 11552 12940
rect 11488 12880 11552 12884
rect 18112 12940 18176 12944
rect 18112 12884 18116 12940
rect 18116 12884 18172 12940
rect 18172 12884 18176 12940
rect 18112 12880 18176 12884
rect 18192 12940 18256 12944
rect 18192 12884 18196 12940
rect 18196 12884 18252 12940
rect 18252 12884 18256 12940
rect 18192 12880 18256 12884
rect 18272 12940 18336 12944
rect 18272 12884 18276 12940
rect 18276 12884 18332 12940
rect 18332 12884 18336 12940
rect 18272 12880 18336 12884
rect 18352 12940 18416 12944
rect 18352 12884 18356 12940
rect 18356 12884 18412 12940
rect 18412 12884 18416 12940
rect 18352 12880 18416 12884
rect 7816 12396 7880 12400
rect 7816 12340 7820 12396
rect 7820 12340 7876 12396
rect 7876 12340 7880 12396
rect 7816 12336 7880 12340
rect 7896 12396 7960 12400
rect 7896 12340 7900 12396
rect 7900 12340 7956 12396
rect 7956 12340 7960 12396
rect 7896 12336 7960 12340
rect 7976 12396 8040 12400
rect 7976 12340 7980 12396
rect 7980 12340 8036 12396
rect 8036 12340 8040 12396
rect 7976 12336 8040 12340
rect 8056 12396 8120 12400
rect 8056 12340 8060 12396
rect 8060 12340 8116 12396
rect 8116 12340 8120 12396
rect 8056 12336 8120 12340
rect 14680 12396 14744 12400
rect 14680 12340 14684 12396
rect 14684 12340 14740 12396
rect 14740 12340 14744 12396
rect 14680 12336 14744 12340
rect 14760 12396 14824 12400
rect 14760 12340 14764 12396
rect 14764 12340 14820 12396
rect 14820 12340 14824 12396
rect 14760 12336 14824 12340
rect 14840 12396 14904 12400
rect 14840 12340 14844 12396
rect 14844 12340 14900 12396
rect 14900 12340 14904 12396
rect 14840 12336 14904 12340
rect 14920 12396 14984 12400
rect 14920 12340 14924 12396
rect 14924 12340 14980 12396
rect 14980 12340 14984 12396
rect 14920 12336 14984 12340
rect 4384 11852 4448 11856
rect 4384 11796 4388 11852
rect 4388 11796 4444 11852
rect 4444 11796 4448 11852
rect 4384 11792 4448 11796
rect 4464 11852 4528 11856
rect 4464 11796 4468 11852
rect 4468 11796 4524 11852
rect 4524 11796 4528 11852
rect 4464 11792 4528 11796
rect 4544 11852 4608 11856
rect 4544 11796 4548 11852
rect 4548 11796 4604 11852
rect 4604 11796 4608 11852
rect 4544 11792 4608 11796
rect 4624 11852 4688 11856
rect 4624 11796 4628 11852
rect 4628 11796 4684 11852
rect 4684 11796 4688 11852
rect 4624 11792 4688 11796
rect 11248 11852 11312 11856
rect 11248 11796 11252 11852
rect 11252 11796 11308 11852
rect 11308 11796 11312 11852
rect 11248 11792 11312 11796
rect 11328 11852 11392 11856
rect 11328 11796 11332 11852
rect 11332 11796 11388 11852
rect 11388 11796 11392 11852
rect 11328 11792 11392 11796
rect 11408 11852 11472 11856
rect 11408 11796 11412 11852
rect 11412 11796 11468 11852
rect 11468 11796 11472 11852
rect 11408 11792 11472 11796
rect 11488 11852 11552 11856
rect 11488 11796 11492 11852
rect 11492 11796 11548 11852
rect 11548 11796 11552 11852
rect 11488 11792 11552 11796
rect 18112 11852 18176 11856
rect 18112 11796 18116 11852
rect 18116 11796 18172 11852
rect 18172 11796 18176 11852
rect 18112 11792 18176 11796
rect 18192 11852 18256 11856
rect 18192 11796 18196 11852
rect 18196 11796 18252 11852
rect 18252 11796 18256 11852
rect 18192 11792 18256 11796
rect 18272 11852 18336 11856
rect 18272 11796 18276 11852
rect 18276 11796 18332 11852
rect 18332 11796 18336 11852
rect 18272 11792 18336 11796
rect 18352 11852 18416 11856
rect 18352 11796 18356 11852
rect 18356 11796 18412 11852
rect 18412 11796 18416 11852
rect 18352 11792 18416 11796
rect 7816 11308 7880 11312
rect 7816 11252 7820 11308
rect 7820 11252 7876 11308
rect 7876 11252 7880 11308
rect 7816 11248 7880 11252
rect 7896 11308 7960 11312
rect 7896 11252 7900 11308
rect 7900 11252 7956 11308
rect 7956 11252 7960 11308
rect 7896 11248 7960 11252
rect 7976 11308 8040 11312
rect 7976 11252 7980 11308
rect 7980 11252 8036 11308
rect 8036 11252 8040 11308
rect 7976 11248 8040 11252
rect 8056 11308 8120 11312
rect 8056 11252 8060 11308
rect 8060 11252 8116 11308
rect 8116 11252 8120 11308
rect 8056 11248 8120 11252
rect 14680 11308 14744 11312
rect 14680 11252 14684 11308
rect 14684 11252 14740 11308
rect 14740 11252 14744 11308
rect 14680 11248 14744 11252
rect 14760 11308 14824 11312
rect 14760 11252 14764 11308
rect 14764 11252 14820 11308
rect 14820 11252 14824 11308
rect 14760 11248 14824 11252
rect 14840 11308 14904 11312
rect 14840 11252 14844 11308
rect 14844 11252 14900 11308
rect 14900 11252 14904 11308
rect 14840 11248 14904 11252
rect 14920 11308 14984 11312
rect 14920 11252 14924 11308
rect 14924 11252 14980 11308
rect 14980 11252 14984 11308
rect 14920 11248 14984 11252
rect 4384 10764 4448 10768
rect 4384 10708 4388 10764
rect 4388 10708 4444 10764
rect 4444 10708 4448 10764
rect 4384 10704 4448 10708
rect 4464 10764 4528 10768
rect 4464 10708 4468 10764
rect 4468 10708 4524 10764
rect 4524 10708 4528 10764
rect 4464 10704 4528 10708
rect 4544 10764 4608 10768
rect 4544 10708 4548 10764
rect 4548 10708 4604 10764
rect 4604 10708 4608 10764
rect 4544 10704 4608 10708
rect 4624 10764 4688 10768
rect 4624 10708 4628 10764
rect 4628 10708 4684 10764
rect 4684 10708 4688 10764
rect 4624 10704 4688 10708
rect 11248 10764 11312 10768
rect 11248 10708 11252 10764
rect 11252 10708 11308 10764
rect 11308 10708 11312 10764
rect 11248 10704 11312 10708
rect 11328 10764 11392 10768
rect 11328 10708 11332 10764
rect 11332 10708 11388 10764
rect 11388 10708 11392 10764
rect 11328 10704 11392 10708
rect 11408 10764 11472 10768
rect 11408 10708 11412 10764
rect 11412 10708 11468 10764
rect 11468 10708 11472 10764
rect 11408 10704 11472 10708
rect 11488 10764 11552 10768
rect 11488 10708 11492 10764
rect 11492 10708 11548 10764
rect 11548 10708 11552 10764
rect 11488 10704 11552 10708
rect 18112 10764 18176 10768
rect 18112 10708 18116 10764
rect 18116 10708 18172 10764
rect 18172 10708 18176 10764
rect 18112 10704 18176 10708
rect 18192 10764 18256 10768
rect 18192 10708 18196 10764
rect 18196 10708 18252 10764
rect 18252 10708 18256 10764
rect 18192 10704 18256 10708
rect 18272 10764 18336 10768
rect 18272 10708 18276 10764
rect 18276 10708 18332 10764
rect 18332 10708 18336 10764
rect 18272 10704 18336 10708
rect 18352 10764 18416 10768
rect 18352 10708 18356 10764
rect 18356 10708 18412 10764
rect 18412 10708 18416 10764
rect 18352 10704 18416 10708
rect 7816 10220 7880 10224
rect 7816 10164 7820 10220
rect 7820 10164 7876 10220
rect 7876 10164 7880 10220
rect 7816 10160 7880 10164
rect 7896 10220 7960 10224
rect 7896 10164 7900 10220
rect 7900 10164 7956 10220
rect 7956 10164 7960 10220
rect 7896 10160 7960 10164
rect 7976 10220 8040 10224
rect 7976 10164 7980 10220
rect 7980 10164 8036 10220
rect 8036 10164 8040 10220
rect 7976 10160 8040 10164
rect 8056 10220 8120 10224
rect 8056 10164 8060 10220
rect 8060 10164 8116 10220
rect 8116 10164 8120 10220
rect 8056 10160 8120 10164
rect 14680 10220 14744 10224
rect 14680 10164 14684 10220
rect 14684 10164 14740 10220
rect 14740 10164 14744 10220
rect 14680 10160 14744 10164
rect 14760 10220 14824 10224
rect 14760 10164 14764 10220
rect 14764 10164 14820 10220
rect 14820 10164 14824 10220
rect 14760 10160 14824 10164
rect 14840 10220 14904 10224
rect 14840 10164 14844 10220
rect 14844 10164 14900 10220
rect 14900 10164 14904 10220
rect 14840 10160 14904 10164
rect 14920 10220 14984 10224
rect 14920 10164 14924 10220
rect 14924 10164 14980 10220
rect 14980 10164 14984 10220
rect 14920 10160 14984 10164
rect 4384 9676 4448 9680
rect 4384 9620 4388 9676
rect 4388 9620 4444 9676
rect 4444 9620 4448 9676
rect 4384 9616 4448 9620
rect 4464 9676 4528 9680
rect 4464 9620 4468 9676
rect 4468 9620 4524 9676
rect 4524 9620 4528 9676
rect 4464 9616 4528 9620
rect 4544 9676 4608 9680
rect 4544 9620 4548 9676
rect 4548 9620 4604 9676
rect 4604 9620 4608 9676
rect 4544 9616 4608 9620
rect 4624 9676 4688 9680
rect 4624 9620 4628 9676
rect 4628 9620 4684 9676
rect 4684 9620 4688 9676
rect 4624 9616 4688 9620
rect 11248 9676 11312 9680
rect 11248 9620 11252 9676
rect 11252 9620 11308 9676
rect 11308 9620 11312 9676
rect 11248 9616 11312 9620
rect 11328 9676 11392 9680
rect 11328 9620 11332 9676
rect 11332 9620 11388 9676
rect 11388 9620 11392 9676
rect 11328 9616 11392 9620
rect 11408 9676 11472 9680
rect 11408 9620 11412 9676
rect 11412 9620 11468 9676
rect 11468 9620 11472 9676
rect 11408 9616 11472 9620
rect 11488 9676 11552 9680
rect 11488 9620 11492 9676
rect 11492 9620 11548 9676
rect 11548 9620 11552 9676
rect 11488 9616 11552 9620
rect 18112 9676 18176 9680
rect 18112 9620 18116 9676
rect 18116 9620 18172 9676
rect 18172 9620 18176 9676
rect 18112 9616 18176 9620
rect 18192 9676 18256 9680
rect 18192 9620 18196 9676
rect 18196 9620 18252 9676
rect 18252 9620 18256 9676
rect 18192 9616 18256 9620
rect 18272 9676 18336 9680
rect 18272 9620 18276 9676
rect 18276 9620 18332 9676
rect 18332 9620 18336 9676
rect 18272 9616 18336 9620
rect 18352 9676 18416 9680
rect 18352 9620 18356 9676
rect 18356 9620 18412 9676
rect 18412 9620 18416 9676
rect 18352 9616 18416 9620
rect 18828 9412 18892 9476
rect 7816 9132 7880 9136
rect 7816 9076 7820 9132
rect 7820 9076 7876 9132
rect 7876 9076 7880 9132
rect 7816 9072 7880 9076
rect 7896 9132 7960 9136
rect 7896 9076 7900 9132
rect 7900 9076 7956 9132
rect 7956 9076 7960 9132
rect 7896 9072 7960 9076
rect 7976 9132 8040 9136
rect 7976 9076 7980 9132
rect 7980 9076 8036 9132
rect 8036 9076 8040 9132
rect 7976 9072 8040 9076
rect 8056 9132 8120 9136
rect 8056 9076 8060 9132
rect 8060 9076 8116 9132
rect 8116 9076 8120 9132
rect 8056 9072 8120 9076
rect 14680 9132 14744 9136
rect 14680 9076 14684 9132
rect 14684 9076 14740 9132
rect 14740 9076 14744 9132
rect 14680 9072 14744 9076
rect 14760 9132 14824 9136
rect 14760 9076 14764 9132
rect 14764 9076 14820 9132
rect 14820 9076 14824 9132
rect 14760 9072 14824 9076
rect 14840 9132 14904 9136
rect 14840 9076 14844 9132
rect 14844 9076 14900 9132
rect 14900 9076 14904 9132
rect 14840 9072 14904 9076
rect 14920 9132 14984 9136
rect 14920 9076 14924 9132
rect 14924 9076 14980 9132
rect 14980 9076 14984 9132
rect 14920 9072 14984 9076
rect 4384 8588 4448 8592
rect 4384 8532 4388 8588
rect 4388 8532 4444 8588
rect 4444 8532 4448 8588
rect 4384 8528 4448 8532
rect 4464 8588 4528 8592
rect 4464 8532 4468 8588
rect 4468 8532 4524 8588
rect 4524 8532 4528 8588
rect 4464 8528 4528 8532
rect 4544 8588 4608 8592
rect 4544 8532 4548 8588
rect 4548 8532 4604 8588
rect 4604 8532 4608 8588
rect 4544 8528 4608 8532
rect 4624 8588 4688 8592
rect 4624 8532 4628 8588
rect 4628 8532 4684 8588
rect 4684 8532 4688 8588
rect 4624 8528 4688 8532
rect 11248 8588 11312 8592
rect 11248 8532 11252 8588
rect 11252 8532 11308 8588
rect 11308 8532 11312 8588
rect 11248 8528 11312 8532
rect 11328 8588 11392 8592
rect 11328 8532 11332 8588
rect 11332 8532 11388 8588
rect 11388 8532 11392 8588
rect 11328 8528 11392 8532
rect 11408 8588 11472 8592
rect 11408 8532 11412 8588
rect 11412 8532 11468 8588
rect 11468 8532 11472 8588
rect 11408 8528 11472 8532
rect 11488 8588 11552 8592
rect 11488 8532 11492 8588
rect 11492 8532 11548 8588
rect 11548 8532 11552 8588
rect 11488 8528 11552 8532
rect 18112 8588 18176 8592
rect 18112 8532 18116 8588
rect 18116 8532 18172 8588
rect 18172 8532 18176 8588
rect 18112 8528 18176 8532
rect 18192 8588 18256 8592
rect 18192 8532 18196 8588
rect 18196 8532 18252 8588
rect 18252 8532 18256 8588
rect 18192 8528 18256 8532
rect 18272 8588 18336 8592
rect 18272 8532 18276 8588
rect 18276 8532 18332 8588
rect 18332 8532 18336 8588
rect 18272 8528 18336 8532
rect 18352 8588 18416 8592
rect 18352 8532 18356 8588
rect 18356 8532 18412 8588
rect 18412 8532 18416 8588
rect 18352 8528 18416 8532
rect 7816 8044 7880 8048
rect 7816 7988 7820 8044
rect 7820 7988 7876 8044
rect 7876 7988 7880 8044
rect 7816 7984 7880 7988
rect 7896 8044 7960 8048
rect 7896 7988 7900 8044
rect 7900 7988 7956 8044
rect 7956 7988 7960 8044
rect 7896 7984 7960 7988
rect 7976 8044 8040 8048
rect 7976 7988 7980 8044
rect 7980 7988 8036 8044
rect 8036 7988 8040 8044
rect 7976 7984 8040 7988
rect 8056 8044 8120 8048
rect 8056 7988 8060 8044
rect 8060 7988 8116 8044
rect 8116 7988 8120 8044
rect 8056 7984 8120 7988
rect 14680 8044 14744 8048
rect 14680 7988 14684 8044
rect 14684 7988 14740 8044
rect 14740 7988 14744 8044
rect 14680 7984 14744 7988
rect 14760 8044 14824 8048
rect 14760 7988 14764 8044
rect 14764 7988 14820 8044
rect 14820 7988 14824 8044
rect 14760 7984 14824 7988
rect 14840 8044 14904 8048
rect 14840 7988 14844 8044
rect 14844 7988 14900 8044
rect 14900 7988 14904 8044
rect 14840 7984 14904 7988
rect 14920 8044 14984 8048
rect 14920 7988 14924 8044
rect 14924 7988 14980 8044
rect 14980 7988 14984 8044
rect 14920 7984 14984 7988
rect 4384 7500 4448 7504
rect 4384 7444 4388 7500
rect 4388 7444 4444 7500
rect 4444 7444 4448 7500
rect 4384 7440 4448 7444
rect 4464 7500 4528 7504
rect 4464 7444 4468 7500
rect 4468 7444 4524 7500
rect 4524 7444 4528 7500
rect 4464 7440 4528 7444
rect 4544 7500 4608 7504
rect 4544 7444 4548 7500
rect 4548 7444 4604 7500
rect 4604 7444 4608 7500
rect 4544 7440 4608 7444
rect 4624 7500 4688 7504
rect 4624 7444 4628 7500
rect 4628 7444 4684 7500
rect 4684 7444 4688 7500
rect 4624 7440 4688 7444
rect 11248 7500 11312 7504
rect 11248 7444 11252 7500
rect 11252 7444 11308 7500
rect 11308 7444 11312 7500
rect 11248 7440 11312 7444
rect 11328 7500 11392 7504
rect 11328 7444 11332 7500
rect 11332 7444 11388 7500
rect 11388 7444 11392 7500
rect 11328 7440 11392 7444
rect 11408 7500 11472 7504
rect 11408 7444 11412 7500
rect 11412 7444 11468 7500
rect 11468 7444 11472 7500
rect 11408 7440 11472 7444
rect 11488 7500 11552 7504
rect 11488 7444 11492 7500
rect 11492 7444 11548 7500
rect 11548 7444 11552 7500
rect 11488 7440 11552 7444
rect 18112 7500 18176 7504
rect 18112 7444 18116 7500
rect 18116 7444 18172 7500
rect 18172 7444 18176 7500
rect 18112 7440 18176 7444
rect 18192 7500 18256 7504
rect 18192 7444 18196 7500
rect 18196 7444 18252 7500
rect 18252 7444 18256 7500
rect 18192 7440 18256 7444
rect 18272 7500 18336 7504
rect 18272 7444 18276 7500
rect 18276 7444 18332 7500
rect 18332 7444 18336 7500
rect 18272 7440 18336 7444
rect 18352 7500 18416 7504
rect 18352 7444 18356 7500
rect 18356 7444 18412 7500
rect 18412 7444 18416 7500
rect 18352 7440 18416 7444
rect 7816 6956 7880 6960
rect 7816 6900 7820 6956
rect 7820 6900 7876 6956
rect 7876 6900 7880 6956
rect 7816 6896 7880 6900
rect 7896 6956 7960 6960
rect 7896 6900 7900 6956
rect 7900 6900 7956 6956
rect 7956 6900 7960 6956
rect 7896 6896 7960 6900
rect 7976 6956 8040 6960
rect 7976 6900 7980 6956
rect 7980 6900 8036 6956
rect 8036 6900 8040 6956
rect 7976 6896 8040 6900
rect 8056 6956 8120 6960
rect 8056 6900 8060 6956
rect 8060 6900 8116 6956
rect 8116 6900 8120 6956
rect 8056 6896 8120 6900
rect 14680 6956 14744 6960
rect 14680 6900 14684 6956
rect 14684 6900 14740 6956
rect 14740 6900 14744 6956
rect 14680 6896 14744 6900
rect 14760 6956 14824 6960
rect 14760 6900 14764 6956
rect 14764 6900 14820 6956
rect 14820 6900 14824 6956
rect 14760 6896 14824 6900
rect 14840 6956 14904 6960
rect 14840 6900 14844 6956
rect 14844 6900 14900 6956
rect 14900 6900 14904 6956
rect 14840 6896 14904 6900
rect 14920 6956 14984 6960
rect 14920 6900 14924 6956
rect 14924 6900 14980 6956
rect 14980 6900 14984 6956
rect 14920 6896 14984 6900
rect 4384 6412 4448 6416
rect 4384 6356 4388 6412
rect 4388 6356 4444 6412
rect 4444 6356 4448 6412
rect 4384 6352 4448 6356
rect 4464 6412 4528 6416
rect 4464 6356 4468 6412
rect 4468 6356 4524 6412
rect 4524 6356 4528 6412
rect 4464 6352 4528 6356
rect 4544 6412 4608 6416
rect 4544 6356 4548 6412
rect 4548 6356 4604 6412
rect 4604 6356 4608 6412
rect 4544 6352 4608 6356
rect 4624 6412 4688 6416
rect 4624 6356 4628 6412
rect 4628 6356 4684 6412
rect 4684 6356 4688 6412
rect 4624 6352 4688 6356
rect 11248 6412 11312 6416
rect 11248 6356 11252 6412
rect 11252 6356 11308 6412
rect 11308 6356 11312 6412
rect 11248 6352 11312 6356
rect 11328 6412 11392 6416
rect 11328 6356 11332 6412
rect 11332 6356 11388 6412
rect 11388 6356 11392 6412
rect 11328 6352 11392 6356
rect 11408 6412 11472 6416
rect 11408 6356 11412 6412
rect 11412 6356 11468 6412
rect 11468 6356 11472 6412
rect 11408 6352 11472 6356
rect 11488 6412 11552 6416
rect 11488 6356 11492 6412
rect 11492 6356 11548 6412
rect 11548 6356 11552 6412
rect 11488 6352 11552 6356
rect 18112 6412 18176 6416
rect 18112 6356 18116 6412
rect 18116 6356 18172 6412
rect 18172 6356 18176 6412
rect 18112 6352 18176 6356
rect 18192 6412 18256 6416
rect 18192 6356 18196 6412
rect 18196 6356 18252 6412
rect 18252 6356 18256 6412
rect 18192 6352 18256 6356
rect 18272 6412 18336 6416
rect 18272 6356 18276 6412
rect 18276 6356 18332 6412
rect 18332 6356 18336 6412
rect 18272 6352 18336 6356
rect 18352 6412 18416 6416
rect 18352 6356 18356 6412
rect 18356 6356 18412 6412
rect 18412 6356 18416 6412
rect 18352 6352 18416 6356
rect 7816 5868 7880 5872
rect 7816 5812 7820 5868
rect 7820 5812 7876 5868
rect 7876 5812 7880 5868
rect 7816 5808 7880 5812
rect 7896 5868 7960 5872
rect 7896 5812 7900 5868
rect 7900 5812 7956 5868
rect 7956 5812 7960 5868
rect 7896 5808 7960 5812
rect 7976 5868 8040 5872
rect 7976 5812 7980 5868
rect 7980 5812 8036 5868
rect 8036 5812 8040 5868
rect 7976 5808 8040 5812
rect 8056 5868 8120 5872
rect 8056 5812 8060 5868
rect 8060 5812 8116 5868
rect 8116 5812 8120 5868
rect 8056 5808 8120 5812
rect 14680 5868 14744 5872
rect 14680 5812 14684 5868
rect 14684 5812 14740 5868
rect 14740 5812 14744 5868
rect 14680 5808 14744 5812
rect 14760 5868 14824 5872
rect 14760 5812 14764 5868
rect 14764 5812 14820 5868
rect 14820 5812 14824 5868
rect 14760 5808 14824 5812
rect 14840 5868 14904 5872
rect 14840 5812 14844 5868
rect 14844 5812 14900 5868
rect 14900 5812 14904 5868
rect 14840 5808 14904 5812
rect 14920 5868 14984 5872
rect 14920 5812 14924 5868
rect 14924 5812 14980 5868
rect 14980 5812 14984 5868
rect 14920 5808 14984 5812
rect 4384 5324 4448 5328
rect 4384 5268 4388 5324
rect 4388 5268 4444 5324
rect 4444 5268 4448 5324
rect 4384 5264 4448 5268
rect 4464 5324 4528 5328
rect 4464 5268 4468 5324
rect 4468 5268 4524 5324
rect 4524 5268 4528 5324
rect 4464 5264 4528 5268
rect 4544 5324 4608 5328
rect 4544 5268 4548 5324
rect 4548 5268 4604 5324
rect 4604 5268 4608 5324
rect 4544 5264 4608 5268
rect 4624 5324 4688 5328
rect 4624 5268 4628 5324
rect 4628 5268 4684 5324
rect 4684 5268 4688 5324
rect 4624 5264 4688 5268
rect 11248 5324 11312 5328
rect 11248 5268 11252 5324
rect 11252 5268 11308 5324
rect 11308 5268 11312 5324
rect 11248 5264 11312 5268
rect 11328 5324 11392 5328
rect 11328 5268 11332 5324
rect 11332 5268 11388 5324
rect 11388 5268 11392 5324
rect 11328 5264 11392 5268
rect 11408 5324 11472 5328
rect 11408 5268 11412 5324
rect 11412 5268 11468 5324
rect 11468 5268 11472 5324
rect 11408 5264 11472 5268
rect 11488 5324 11552 5328
rect 11488 5268 11492 5324
rect 11492 5268 11548 5324
rect 11548 5268 11552 5324
rect 11488 5264 11552 5268
rect 18112 5324 18176 5328
rect 18112 5268 18116 5324
rect 18116 5268 18172 5324
rect 18172 5268 18176 5324
rect 18112 5264 18176 5268
rect 18192 5324 18256 5328
rect 18192 5268 18196 5324
rect 18196 5268 18252 5324
rect 18252 5268 18256 5324
rect 18192 5264 18256 5268
rect 18272 5324 18336 5328
rect 18272 5268 18276 5324
rect 18276 5268 18332 5324
rect 18332 5268 18336 5324
rect 18272 5264 18336 5268
rect 18352 5324 18416 5328
rect 18352 5268 18356 5324
rect 18356 5268 18412 5324
rect 18412 5268 18416 5324
rect 18352 5264 18416 5268
rect 7816 4780 7880 4784
rect 7816 4724 7820 4780
rect 7820 4724 7876 4780
rect 7876 4724 7880 4780
rect 7816 4720 7880 4724
rect 7896 4780 7960 4784
rect 7896 4724 7900 4780
rect 7900 4724 7956 4780
rect 7956 4724 7960 4780
rect 7896 4720 7960 4724
rect 7976 4780 8040 4784
rect 7976 4724 7980 4780
rect 7980 4724 8036 4780
rect 8036 4724 8040 4780
rect 7976 4720 8040 4724
rect 8056 4780 8120 4784
rect 8056 4724 8060 4780
rect 8060 4724 8116 4780
rect 8116 4724 8120 4780
rect 8056 4720 8120 4724
rect 14680 4780 14744 4784
rect 14680 4724 14684 4780
rect 14684 4724 14740 4780
rect 14740 4724 14744 4780
rect 14680 4720 14744 4724
rect 14760 4780 14824 4784
rect 14760 4724 14764 4780
rect 14764 4724 14820 4780
rect 14820 4724 14824 4780
rect 14760 4720 14824 4724
rect 14840 4780 14904 4784
rect 14840 4724 14844 4780
rect 14844 4724 14900 4780
rect 14900 4724 14904 4780
rect 14840 4720 14904 4724
rect 14920 4780 14984 4784
rect 14920 4724 14924 4780
rect 14924 4724 14980 4780
rect 14980 4724 14984 4780
rect 14920 4720 14984 4724
rect 4384 4236 4448 4240
rect 4384 4180 4388 4236
rect 4388 4180 4444 4236
rect 4444 4180 4448 4236
rect 4384 4176 4448 4180
rect 4464 4236 4528 4240
rect 4464 4180 4468 4236
rect 4468 4180 4524 4236
rect 4524 4180 4528 4236
rect 4464 4176 4528 4180
rect 4544 4236 4608 4240
rect 4544 4180 4548 4236
rect 4548 4180 4604 4236
rect 4604 4180 4608 4236
rect 4544 4176 4608 4180
rect 4624 4236 4688 4240
rect 4624 4180 4628 4236
rect 4628 4180 4684 4236
rect 4684 4180 4688 4236
rect 4624 4176 4688 4180
rect 11248 4236 11312 4240
rect 11248 4180 11252 4236
rect 11252 4180 11308 4236
rect 11308 4180 11312 4236
rect 11248 4176 11312 4180
rect 11328 4236 11392 4240
rect 11328 4180 11332 4236
rect 11332 4180 11388 4236
rect 11388 4180 11392 4236
rect 11328 4176 11392 4180
rect 11408 4236 11472 4240
rect 11408 4180 11412 4236
rect 11412 4180 11468 4236
rect 11468 4180 11472 4236
rect 11408 4176 11472 4180
rect 11488 4236 11552 4240
rect 11488 4180 11492 4236
rect 11492 4180 11548 4236
rect 11548 4180 11552 4236
rect 11488 4176 11552 4180
rect 18112 4236 18176 4240
rect 18112 4180 18116 4236
rect 18116 4180 18172 4236
rect 18172 4180 18176 4236
rect 18112 4176 18176 4180
rect 18192 4236 18256 4240
rect 18192 4180 18196 4236
rect 18196 4180 18252 4236
rect 18252 4180 18256 4236
rect 18192 4176 18256 4180
rect 18272 4236 18336 4240
rect 18272 4180 18276 4236
rect 18276 4180 18332 4236
rect 18332 4180 18336 4236
rect 18272 4176 18336 4180
rect 18352 4236 18416 4240
rect 18352 4180 18356 4236
rect 18356 4180 18412 4236
rect 18412 4180 18416 4236
rect 18352 4176 18416 4180
rect 7816 3692 7880 3696
rect 7816 3636 7820 3692
rect 7820 3636 7876 3692
rect 7876 3636 7880 3692
rect 7816 3632 7880 3636
rect 7896 3692 7960 3696
rect 7896 3636 7900 3692
rect 7900 3636 7956 3692
rect 7956 3636 7960 3692
rect 7896 3632 7960 3636
rect 7976 3692 8040 3696
rect 7976 3636 7980 3692
rect 7980 3636 8036 3692
rect 8036 3636 8040 3692
rect 7976 3632 8040 3636
rect 8056 3692 8120 3696
rect 8056 3636 8060 3692
rect 8060 3636 8116 3692
rect 8116 3636 8120 3692
rect 8056 3632 8120 3636
rect 14680 3692 14744 3696
rect 14680 3636 14684 3692
rect 14684 3636 14740 3692
rect 14740 3636 14744 3692
rect 14680 3632 14744 3636
rect 14760 3692 14824 3696
rect 14760 3636 14764 3692
rect 14764 3636 14820 3692
rect 14820 3636 14824 3692
rect 14760 3632 14824 3636
rect 14840 3692 14904 3696
rect 14840 3636 14844 3692
rect 14844 3636 14900 3692
rect 14900 3636 14904 3692
rect 14840 3632 14904 3636
rect 14920 3692 14984 3696
rect 14920 3636 14924 3692
rect 14924 3636 14980 3692
rect 14980 3636 14984 3692
rect 14920 3632 14984 3636
rect 4384 3148 4448 3152
rect 4384 3092 4388 3148
rect 4388 3092 4444 3148
rect 4444 3092 4448 3148
rect 4384 3088 4448 3092
rect 4464 3148 4528 3152
rect 4464 3092 4468 3148
rect 4468 3092 4524 3148
rect 4524 3092 4528 3148
rect 4464 3088 4528 3092
rect 4544 3148 4608 3152
rect 4544 3092 4548 3148
rect 4548 3092 4604 3148
rect 4604 3092 4608 3148
rect 4544 3088 4608 3092
rect 4624 3148 4688 3152
rect 4624 3092 4628 3148
rect 4628 3092 4684 3148
rect 4684 3092 4688 3148
rect 4624 3088 4688 3092
rect 11248 3148 11312 3152
rect 11248 3092 11252 3148
rect 11252 3092 11308 3148
rect 11308 3092 11312 3148
rect 11248 3088 11312 3092
rect 11328 3148 11392 3152
rect 11328 3092 11332 3148
rect 11332 3092 11388 3148
rect 11388 3092 11392 3148
rect 11328 3088 11392 3092
rect 11408 3148 11472 3152
rect 11408 3092 11412 3148
rect 11412 3092 11468 3148
rect 11468 3092 11472 3148
rect 11408 3088 11472 3092
rect 11488 3148 11552 3152
rect 11488 3092 11492 3148
rect 11492 3092 11548 3148
rect 11548 3092 11552 3148
rect 11488 3088 11552 3092
rect 18112 3148 18176 3152
rect 18112 3092 18116 3148
rect 18116 3092 18172 3148
rect 18172 3092 18176 3148
rect 18112 3088 18176 3092
rect 18192 3148 18256 3152
rect 18192 3092 18196 3148
rect 18196 3092 18252 3148
rect 18252 3092 18256 3148
rect 18192 3088 18256 3092
rect 18272 3148 18336 3152
rect 18272 3092 18276 3148
rect 18276 3092 18332 3148
rect 18332 3092 18336 3148
rect 18272 3088 18336 3092
rect 18352 3148 18416 3152
rect 18352 3092 18356 3148
rect 18356 3092 18412 3148
rect 18412 3092 18416 3148
rect 18352 3088 18416 3092
rect 7816 2604 7880 2608
rect 7816 2548 7820 2604
rect 7820 2548 7876 2604
rect 7876 2548 7880 2604
rect 7816 2544 7880 2548
rect 7896 2604 7960 2608
rect 7896 2548 7900 2604
rect 7900 2548 7956 2604
rect 7956 2548 7960 2604
rect 7896 2544 7960 2548
rect 7976 2604 8040 2608
rect 7976 2548 7980 2604
rect 7980 2548 8036 2604
rect 8036 2548 8040 2604
rect 7976 2544 8040 2548
rect 8056 2604 8120 2608
rect 8056 2548 8060 2604
rect 8060 2548 8116 2604
rect 8116 2548 8120 2604
rect 8056 2544 8120 2548
rect 14680 2604 14744 2608
rect 14680 2548 14684 2604
rect 14684 2548 14740 2604
rect 14740 2548 14744 2604
rect 14680 2544 14744 2548
rect 14760 2604 14824 2608
rect 14760 2548 14764 2604
rect 14764 2548 14820 2604
rect 14820 2548 14824 2604
rect 14760 2544 14824 2548
rect 14840 2604 14904 2608
rect 14840 2548 14844 2604
rect 14844 2548 14900 2604
rect 14900 2548 14904 2604
rect 14840 2544 14904 2548
rect 14920 2604 14984 2608
rect 14920 2548 14924 2604
rect 14924 2548 14980 2604
rect 14980 2548 14984 2604
rect 14920 2544 14984 2548
rect 4384 2060 4448 2064
rect 4384 2004 4388 2060
rect 4388 2004 4444 2060
rect 4444 2004 4448 2060
rect 4384 2000 4448 2004
rect 4464 2060 4528 2064
rect 4464 2004 4468 2060
rect 4468 2004 4524 2060
rect 4524 2004 4528 2060
rect 4464 2000 4528 2004
rect 4544 2060 4608 2064
rect 4544 2004 4548 2060
rect 4548 2004 4604 2060
rect 4604 2004 4608 2060
rect 4544 2000 4608 2004
rect 4624 2060 4688 2064
rect 4624 2004 4628 2060
rect 4628 2004 4684 2060
rect 4684 2004 4688 2060
rect 4624 2000 4688 2004
rect 11248 2060 11312 2064
rect 11248 2004 11252 2060
rect 11252 2004 11308 2060
rect 11308 2004 11312 2060
rect 11248 2000 11312 2004
rect 11328 2060 11392 2064
rect 11328 2004 11332 2060
rect 11332 2004 11388 2060
rect 11388 2004 11392 2060
rect 11328 2000 11392 2004
rect 11408 2060 11472 2064
rect 11408 2004 11412 2060
rect 11412 2004 11468 2060
rect 11468 2004 11472 2060
rect 11408 2000 11472 2004
rect 11488 2060 11552 2064
rect 11488 2004 11492 2060
rect 11492 2004 11548 2060
rect 11548 2004 11552 2060
rect 11488 2000 11552 2004
rect 18112 2060 18176 2064
rect 18112 2004 18116 2060
rect 18116 2004 18172 2060
rect 18172 2004 18176 2060
rect 18112 2000 18176 2004
rect 18192 2060 18256 2064
rect 18192 2004 18196 2060
rect 18196 2004 18252 2060
rect 18252 2004 18256 2060
rect 18192 2000 18256 2004
rect 18272 2060 18336 2064
rect 18272 2004 18276 2060
rect 18276 2004 18332 2060
rect 18332 2004 18336 2060
rect 18272 2000 18336 2004
rect 18352 2060 18416 2064
rect 18352 2004 18356 2060
rect 18356 2004 18412 2060
rect 18412 2004 18416 2060
rect 18352 2000 18416 2004
rect 18828 1796 18892 1860
<< metal4 >>
rect 4376 19472 4696 20032
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 18384 4696 19408
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 17296 4696 18320
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 16208 4696 17232
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 15120 4696 16144
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 14032 4696 15056
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 12944 4696 13968
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 11856 4696 12880
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 10768 4696 11792
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 9680 4696 10704
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 8592 4696 9616
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 7504 4696 8528
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 6416 4696 7440
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 5328 4696 6352
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 4240 4696 5264
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 3152 4696 4176
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 2064 4696 3088
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1984 4696 2000
rect 7808 20016 8128 20032
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 18928 8128 19952
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 17840 8128 18864
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 16752 8128 17776
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 15664 8128 16688
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 14576 8128 15600
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 13488 8128 14512
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 12400 8128 13424
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 11312 8128 12336
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 10224 8128 11248
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 9136 8128 10160
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 8048 8128 9072
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 6960 8128 7984
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 5872 8128 6896
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 4784 8128 5808
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 3696 8128 4720
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 2608 8128 3632
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 1984 8128 2544
rect 11240 19472 11560 20032
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 18384 11560 19408
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 17296 11560 18320
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 16208 11560 17232
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 15120 11560 16144
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 14032 11560 15056
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 12944 11560 13968
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 11856 11560 12880
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 10768 11560 11792
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 9680 11560 10704
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 8592 11560 9616
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 7504 11560 8528
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 6416 11560 7440
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 5328 11560 6352
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 4240 11560 5264
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 3152 11560 4176
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 2064 11560 3088
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1984 11560 2000
rect 14672 20016 14992 20032
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 14672 18928 14992 19952
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 17840 14992 18864
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 14672 16752 14992 17776
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 15664 14992 16688
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 14576 14992 15600
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 14672 13488 14992 14512
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 12400 14992 13424
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 11312 14992 12336
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 10224 14992 11248
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 9136 14992 10160
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 14672 8048 14992 9072
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 6960 14992 7984
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 5872 14992 6896
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 14672 4784 14992 5808
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 3696 14992 4720
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 2608 14992 3632
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 1984 14992 2544
rect 18104 19472 18424 20032
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 18384 18424 19408
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 17296 18424 18320
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 18104 16208 18424 17232
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 15120 18424 16144
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 14032 18424 15056
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 12944 18424 13968
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 11856 18424 12880
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 18104 10768 18424 11792
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 9680 18424 10704
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 8592 18424 9616
rect 18827 9476 18893 9477
rect 18827 9412 18828 9476
rect 18892 9412 18893 9476
rect 18827 9411 18893 9412
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 18104 7504 18424 8528
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 6416 18424 7440
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 18104 5328 18424 6352
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 4240 18424 5264
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 3152 18424 4176
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 18104 2064 18424 3088
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1984 18424 2000
rect 18830 1861 18890 9411
rect 18827 1860 18893 1861
rect 18827 1796 18828 1860
rect 18892 1796 18893 1860
rect 18827 1795 18893 1796
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1606821651
transform 1 0 3588 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1606821651
transform 1 0 4048 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1606821651
transform 1 0 5152 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1606821651
transform 1 0 6256 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606821651
transform 1 0 8004 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1606821651
transform 1 0 7360 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1606821651
transform 1 0 8464 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606821651
transform 1 0 9108 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1606821651
transform 1 0 9660 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606821651
transform 1 0 11960 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1606821651
transform 1 0 10764 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1606821651
transform 1 0 11868 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606821651
transform 1 0 13708 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1606821651
transform 1 0 12972 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1606821651
transform 1 0 14076 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606821651
transform 1 0 14812 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1606821651
transform 1 0 15272 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1606821651
transform 1 0 16376 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606821651
transform 1 0 16560 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606821651
transform 1 0 17664 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1606821651
transform 1 0 17480 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606821651
transform 1 0 19412 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1606821651
transform 1 0 18584 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1606821651
transform 1 0 19688 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 20792 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606821651
transform 1 0 20516 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 21160 0 -1 2576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606821651
transform 1 0 20884 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 21252 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1606821651
transform 1 0 4692 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 6716 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5796 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1606821651
transform 1 0 6532 0 -1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1606821651
transform 1 0 6808 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1606821651
transform 1 0 7912 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1606821651
transform 1 0 9016 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1606821651
transform 1 0 10120 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 12328 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1606821651
transform 1 0 11224 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1606821651
transform 1 0 12420 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1606821651
transform 1 0 13524 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1606821651
transform 1 0 14628 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1606821651
transform 1 0 15732 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 17940 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1606821651
transform 1 0 16836 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1606821651
transform 1 0 18032 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1606821651
transform 1 0 19136 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1606821651
transform 1 0 20240 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 3956 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1606821651
transform 1 0 4048 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1606821651
transform 1 0 5152 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1606821651
transform 1 0 6256 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1606821651
transform 1 0 7360 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1606821651
transform 1 0 8464 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 9568 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1606821651
transform 1 0 9660 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1606821651
transform 1 0 10764 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1606821651
transform 1 0 11868 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1606821651
transform 1 0 12972 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1606821651
transform 1 0 14076 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 15180 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1606821651
transform 1 0 15272 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1606821651
transform 1 0 16376 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1606821651
transform 1 0 17480 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1606821651
transform 1 0 18584 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1606821651
transform 1 0 19688 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 20792 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1606821651
transform 1 0 20884 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1606821651
transform 1 0 21252 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1606821651
transform 1 0 4692 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 6716 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1606821651
transform 1 0 5796 0 -1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1606821651
transform 1 0 6532 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1606821651
transform 1 0 6808 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1606821651
transform 1 0 7912 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1606821651
transform 1 0 9016 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1606821651
transform 1 0 10120 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 12328 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1606821651
transform 1 0 11224 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1606821651
transform 1 0 12420 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1606821651
transform 1 0 13524 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1606821651
transform 1 0 14628 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1606821651
transform 1 0 15732 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 17940 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1606821651
transform 1 0 16836 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1606821651
transform 1 0 18032 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1606821651
transform 1 0 19136 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_208
timestamp 1606821651
transform 1 0 20240 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 20516 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 3956 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1606821651
transform 1 0 4048 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1606821651
transform 1 0 5152 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1606821651
transform 1 0 6256 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1606821651
transform 1 0 7360 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1606821651
transform 1 0 8464 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 9568 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1606821651
transform 1 0 9660 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1606821651
transform 1 0 10764 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1606821651
transform 1 0 11868 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1606821651
transform 1 0 12972 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1606821651
transform 1 0 14076 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 15180 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1606821651
transform 1 0 15272 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1606821651
transform 1 0 16376 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1606821651
transform 1 0 17480 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1606821651
transform 1 0 18584 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1606821651
transform 1 0 19688 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 20792 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1606821651
transform 1 0 20884 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606821651
transform 1 0 21252 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 3956 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1606821651
transform 1 0 4692 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1606821651
transform 1 0 4048 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 6716 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1606821651
transform 1 0 5796 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1606821651
transform 1 0 6532 0 -1 5840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1606821651
transform 1 0 6808 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1606821651
transform 1 0 5152 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1606821651
transform 1 0 6256 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1606821651
transform 1 0 7912 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1606821651
transform 1 0 7360 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1606821651
transform 1 0 8464 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 9568 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1606821651
transform 1 0 9016 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1606821651
transform 1 0 10120 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1606821651
transform 1 0 9660 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 12328 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1606821651
transform 1 0 11224 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1606821651
transform 1 0 12420 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1606821651
transform 1 0 10764 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1606821651
transform 1 0 11868 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1606821651
transform 1 0 13524 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1606821651
transform 1 0 12972 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1606821651
transform 1 0 14076 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 15180 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1606821651
transform 1 0 14628 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1606821651
transform 1 0 15732 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1606821651
transform 1 0 15272 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1606821651
transform 1 0 16376 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 17940 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1606821651
transform 1 0 16836 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1606821651
transform 1 0 18032 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1606821651
transform 1 0 17480 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1606821651
transform 1 0 19136 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_208
timestamp 1606821651
transform 1 0 20240 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1606821651
transform 1 0 18584 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1606821651
transform 1 0 19688 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606821651
transform 1 0 20516 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 20792 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1606821651
transform 1 0 20884 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1606821651
transform 1 0 21252 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606821651
transform 1 0 2484 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1606821651
transform 1 0 4692 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 6716 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1606821651
transform 1 0 5796 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1606821651
transform 1 0 6532 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_62
timestamp 1606821651
transform 1 0 6808 0 -1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7360 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10580 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_84
timestamp 1606821651
transform 1 0 8832 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_96
timestamp 1606821651
transform 1 0 9936 0 -1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_102
timestamp 1606821651
transform 1 0 10488 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 12328 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_112
timestamp 1606821651
transform 1 0 11408 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1606821651
transform 1 0 12144 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1606821651
transform 1 0 12420 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14076 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_135
timestamp 1606821651
transform 1 0 13524 0 -1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_150
timestamp 1606821651
transform 1 0 14904 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_162
timestamp 1606821651
transform 1 0 16008 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 17940 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_174
timestamp 1606821651
transform 1 0 17112 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1606821651
transform 1 0 17848 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1606821651
transform 1 0 18032 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1606821651
transform 1 0 19136 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_208
timestamp 1606821651
transform 1 0 20240 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606821651
transform 1 0 20516 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 3956 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1606821651
transform 1 0 3588 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1606821651
transform 1 0 4048 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1606821651
transform 1 0 5152 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1606821651
transform 1 0 6256 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1606821651
transform 1 0 7360 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1606821651
transform 1 0 8464 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 9568 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11316 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1606821651
transform 1 0 11132 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12972 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1606821651
transform 1 0 12788 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1606821651
transform 1 0 14444 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14628 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 15180 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_150
timestamp 1606821651
transform 1 0 14904 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1606821651
transform 1 0 16744 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1606821651
transform 1 0 17756 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1606821651
transform 1 0 18860 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_205
timestamp 1606821651
transform 1 0 19964 0 1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 20792 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_213
timestamp 1606821651
transform 1 0 20700 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1606821651
transform 1 0 20884 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606821651
transform 1 0 21252 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606821651
transform 1 0 2484 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1606821651
transform 1 0 3588 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1606821651
transform 1 0 4692 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 6716 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1606821651
transform 1 0 5796 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1606821651
transform 1 0 6532 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1606821651
transform 1 0 6808 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1606821651
transform 1 0 7912 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10396 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_86
timestamp 1606821651
transform 1 0 9016 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_98
timestamp 1606821651
transform 1 0 10120 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11408 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 12328 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp 1606821651
transform 1 0 11224 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1606821651
transform 1 0 11960 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1606821651
transform 1 0 12420 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13708 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_135
timestamp 1606821651
transform 1 0 13524 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16284 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_146
timestamp 1606821651
transform 1 0 14536 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_158
timestamp 1606821651
transform 1 0 15640 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_164
timestamp 1606821651
transform 1 0 16192 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 17940 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1606821651
transform 1 0 17756 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606821651
transform 1 0 19964 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1606821651
transform 1 0 19504 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1606821651
transform 1 0 19872 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606821651
transform 1 0 20516 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1606821651
transform 1 0 20332 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606821651
transform 1 0 21252 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606821651
transform 1 0 2484 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 3956 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1606821651
transform 1 0 3588 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1606821651
transform 1 0 4048 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1606821651
transform 1 0 5152 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1606821651
transform 1 0 6256 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1606821651
transform 1 0 7360 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1606821651
transform 1 0 8464 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606821651
transform 1 0 10672 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 9568 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1606821651
transform 1 0 9660 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_101
timestamp 1606821651
transform 1 0 10396 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1606821651
transform 1 0 11316 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1606821651
transform 1 0 10948 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1606821651
transform 1 0 11684 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13340 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_127
timestamp 1606821651
transform 1 0 12788 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1606821651
transform 1 0 13892 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16284 0 1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 15180 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1606821651
transform 1 0 14996 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_154
timestamp 1606821651
transform 1 0 15272 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_162
timestamp 1606821651
transform 1 0 16008 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1606821651
transform 1 0 17296 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_174
timestamp 1606821651
transform 1 0 17112 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_179
timestamp 1606821651
transform 1 0 17572 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606821651
transform 1 0 20240 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_191
timestamp 1606821651
transform 1 0 18676 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_203
timestamp 1606821651
transform 1 0 19780 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_207
timestamp 1606821651
transform 1 0 20148 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 20792 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1606821651
transform 1 0 20608 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1606821651
transform 1 0 20884 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1606821651
transform 1 0 21252 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606821651
transform 1 0 2484 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1606821651
transform 1 0 3588 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1606821651
transform 1 0 4692 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 6716 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1606821651
transform 1 0 5796 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1606821651
transform 1 0 6532 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1606821651
transform 1 0 6808 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8188 0 -1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_74
timestamp 1606821651
transform 1 0 7912 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1606821651
transform 1 0 9660 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10948 0 -1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 12328 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1606821651
transform 1 0 10764 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_116
timestamp 1606821651
transform 1 0 11776 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_123
timestamp 1606821651
transform 1 0 12420 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606821651
transform 1 0 13248 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_131
timestamp 1606821651
transform 1 0 13156 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_136
timestamp 1606821651
transform 1 0 13616 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15456 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_148
timestamp 1606821651
transform 1 0 14720 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_162
timestamp 1606821651
transform 1 0 16008 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18308 0 -1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 17940 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_174
timestamp 1606821651
transform 1 0 17112 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_182
timestamp 1606821651
transform 1 0 17848 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_184
timestamp 1606821651
transform 1 0 18032 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606821651
transform 1 0 19964 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1606821651
transform 1 0 19780 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606821651
transform 1 0 20516 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1606821651
transform 1 0 20332 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606821651
transform 1 0 2484 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606821651
transform 1 0 2484 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 3956 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1606821651
transform 1 0 3588 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1606821651
transform 1 0 4048 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1606821651
transform 1 0 3588 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1606821651
transform 1 0 4692 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 6716 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1606821651
transform 1 0 5152 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1606821651
transform 1 0 6256 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1606821651
transform 1 0 5796 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1606821651
transform 1 0 6532 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1606821651
transform 1 0 6808 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7912 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_68
timestamp 1606821651
transform 1 0 7360 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_74
timestamp 1606821651
transform 1 0 7912 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10028 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 9568 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1606821651
transform 1 0 9384 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1606821651
transform 1 0 9660 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_101
timestamp 1606821651
transform 1 0 10396 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_86
timestamp 1606821651
transform 1 0 9016 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_94
timestamp 1606821651
transform 1 0 9752 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1606821651
transform 1 0 10856 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_111
timestamp 1606821651
transform 1 0 11316 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 11040 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606821651
transform 1 0 11500 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1606821651
transform 1 0 12236 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1606821651
transform 1 0 11868 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_116
timestamp 1606821651
transform 1 0 11776 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 12328 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12328 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1606821651
transform 1 0 12420 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13524 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1606821651
transform 1 0 13156 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_135
timestamp 1606821651
transform 1 0 13524 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606821651
transform 1 0 15272 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15916 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 15180 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1606821651
transform 1 0 14996 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1606821651
transform 1 0 15640 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_147
timestamp 1606821651
transform 1 0 14628 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_159
timestamp 1606821651
transform 1 0 15732 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 17940 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_170
timestamp 1606821651
transform 1 0 16744 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_182
timestamp 1606821651
transform 1 0 17848 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_177
timestamp 1606821651
transform 1 0 17388 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1606821651
transform 1 0 18032 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606821651
transform 1 0 19688 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18492 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18676 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1606821651
transform 1 0 18584 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1606821651
transform 1 0 19504 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_205
timestamp 1606821651
transform 1 0 19964 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_188
timestamp 1606821651
transform 1 0 18400 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1606821651
transform 1 0 19964 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606821651
transform 1 0 20516 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 20792 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_213
timestamp 1606821651
transform 1 0 20700 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606821651
transform 1 0 20884 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606821651
transform 1 0 21252 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606821651
transform 1 0 2484 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 3956 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1606821651
transform 1 0 3588 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1606821651
transform 1 0 4048 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1606821651
transform 1 0 5152 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_56
timestamp 1606821651
transform 1 0 6256 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7176 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_64
timestamp 1606821651
transform 1 0 6992 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_82
timestamp 1606821651
transform 1 0 8648 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 9568 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1606821651
transform 1 0 9384 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1606821651
transform 1 0 9660 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11040 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_105
timestamp 1606821651
transform 1 0 10764 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_117
timestamp 1606821651
transform 1 0 11868 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_125
timestamp 1606821651
transform 1 0 12604 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12696 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_142
timestamp 1606821651
transform 1 0 14168 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 15180 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_150
timestamp 1606821651
transform 1 0 14904 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_154
timestamp 1606821651
transform 1 0 15272 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1606821651
transform 1 0 16376 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16560 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1606821651
transform 1 0 17388 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_185
timestamp 1606821651
transform 1 0 18124 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 20240 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18400 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_197
timestamp 1606821651
transform 1 0 19228 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_205
timestamp 1606821651
transform 1 0 19964 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 20792 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1606821651
transform 1 0 20608 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1606821651
transform 1 0 20884 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1606821651
transform 1 0 21252 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606821651
transform 1 0 2484 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1606821651
transform 1 0 4692 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 6716 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1606821651
transform 1 0 5796 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1606821651
transform 1 0 6532 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1606821651
transform 1 0 6808 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8280 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_74
timestamp 1606821651
transform 1 0 7912 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10672 0 -1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1606821651
transform 1 0 9108 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1606821651
transform 1 0 10212 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_103
timestamp 1606821651
transform 1 0 10580 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 12328 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_110
timestamp 1606821651
transform 1 0 11224 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1606821651
transform 1 0 12420 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13708 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1606821651
transform 1 0 13524 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1606821651
transform 1 0 14720 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15916 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1606821651
transform 1 0 14536 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_151
timestamp 1606821651
transform 1 0 14996 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1606821651
transform 1 0 15732 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 17940 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606821651
transform 1 0 16744 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1606821651
transform 1 0 17756 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1606821651
transform 1 0 18032 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 19964 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 18768 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_201
timestamp 1606821651
transform 1 0 19596 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 20516 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_209
timestamp 1606821651
transform 1 0 20332 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606821651
transform 1 0 2484 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 3956 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1606821651
transform 1 0 3588 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1606821651
transform 1 0 4048 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6716 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1606821651
transform 1 0 5152 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1606821651
transform 1 0 6256 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1606821651
transform 1 0 6624 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8004 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_70
timestamp 1606821651
transform 1 0 7544 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1606821651
transform 1 0 7912 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10396 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 9568 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1606821651
transform 1 0 8832 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1606821651
transform 1 0 9660 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606821651
transform 1 0 11408 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1606821651
transform 1 0 11224 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1606821651
transform 1 0 11684 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13524 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_track_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13248 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1606821651
transform 1 0 12788 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 1606821651
transform 1 0 13156 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_144
timestamp 1606821651
transform 1 0 14352 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 15180 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1606821651
transform 1 0 15088 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1606821651
transform 1 0 15272 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1606821651
transform 1 0 16376 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_178
timestamp 1606821651
transform 1 0 17480 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1606821651
transform 1 0 19044 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 20240 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606821651
transform 1 0 18860 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_198
timestamp 1606821651
transform 1 0 19320 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1606821651
transform 1 0 20056 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 20792 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1606821651
transform 1 0 20608 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1606821651
transform 1 0 20884 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1606821651
transform 1 0 21252 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606821651
transform 1 0 2484 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1606821651
transform 1 0 4692 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 6716 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1606821651
transform 1 0 5796 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1606821651
transform 1 0 6532 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_62
timestamp 1606821651
transform 1 0 6808 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6992 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8740 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_80
timestamp 1606821651
transform 1 0 8464 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10396 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_99
timestamp 1606821651
transform 1 0 10212 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 12328 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_110
timestamp 1606821651
transform 1 0 11224 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14076 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_139
timestamp 1606821651
transform 1 0 13892 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15180 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606821651
transform 1 0 14904 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18032 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 17940 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_169
timestamp 1606821651
transform 1 0 16652 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1606821651
transform 1 0 17756 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 19964 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_193
timestamp 1606821651
transform 1 0 18860 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 20516 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1606821651
transform 1 0 20332 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606821651
transform 1 0 20884 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606821651
transform 1 0 21252 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606821651
transform 1 0 2484 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606821651
transform 1 0 2484 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 3956 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1606821651
transform 1 0 3588 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1606821651
transform 1 0 4048 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1606821651
transform 1 0 3588 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_39
timestamp 1606821651
transform 1 0 4692 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5612 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 6716 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1606821651
transform 1 0 5152 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1606821651
transform 1 0 6256 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_47
timestamp 1606821651
transform 1 0 5428 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_58
timestamp 1606821651
transform 1 0 6440 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1606821651
transform 1 0 6808 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_track_0.prog_clk
timestamp 1606821651
transform 1 0 7544 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_68
timestamp 1606821651
transform 1 0 7360 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_73
timestamp 1606821651
transform 1 0 7820 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1606821651
transform 1 0 7912 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9936 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 9568 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_track_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10028 0 -1 13456
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_19_85
timestamp 1606821651
transform 1 0 8924 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_91
timestamp 1606821651
transform 1 0 9476 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_93
timestamp 1606821651
transform 1 0 9660 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_86
timestamp 1606821651
transform 1 0 9016 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_94
timestamp 1606821651
transform 1 0 9752 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11408 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 12328 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_track_0.prog_clk
timestamp 1606821651
transform 1 0 12420 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1606821651
transform 1 0 11960 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_122
timestamp 1606821651
transform 1 0 12328 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1606821651
transform 1 0 11868 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_121
timestamp 1606821651
transform 1 0 12236 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1606821651
transform 1 0 12420 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12972 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13984 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_126
timestamp 1606821651
transform 1 0 12696 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1606821651
transform 1 0 13800 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_135
timestamp 1606821651
transform 1 0 13524 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 15180 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1606821651
transform 1 0 14812 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1606821651
transform 1 0 15824 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_147
timestamp 1606821651
transform 1 0 14628 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_159
timestamp 1606821651
transform 1 0 15732 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16560 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 17940 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_171
timestamp 1606821651
transform 1 0 16836 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1606821651
transform 1 0 18032 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 19964 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 19964 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 19412 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19136 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18676 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_202
timestamp 1606821651
transform 1 0 19688 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_190
timestamp 1606821651
transform 1 0 18584 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1606821651
transform 1 0 19228 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_203
timestamp 1606821651
transform 1 0 19780 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1606821651
transform 1 0 20332 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1606821651
transform 1 0 20700 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1606821651
transform 1 0 20332 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 20516 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1606821651
transform 1 0 20884 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 20792 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1606821651
transform 1 0 21252 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2208 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1606821651
transform 1 0 2116 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4876 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 3956 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_28
timestamp 1606821651
transform 1 0 3680 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1606821651
transform 1 0 4048 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_40
timestamp 1606821651
transform 1 0 4784 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1606821651
transform 1 0 6532 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1606821651
transform 1 0 6348 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7268 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1606821651
transform 1 0 7176 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1606821651
transform 1 0 8740 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 9568 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_track_0.prog_clk
timestamp 1606821651
transform 1 0 8924 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_88
timestamp 1606821651
transform 1 0 9200 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1606821651
transform 1 0 9660 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10948 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12604 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1606821651
transform 1 0 10764 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606821651
transform 1 0 13616 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1606821651
transform 1 0 13432 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1606821651
transform 1 0 13892 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16376 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 15180 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_151
timestamp 1606821651
transform 1 0 14996 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1606821651
transform 1 0 15272 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 17388 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1606821651
transform 1 0 17204 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_186
timestamp 1606821651
transform 1 0 18216 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 20240 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 18400 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_192
timestamp 1606821651
transform 1 0 18768 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_204
timestamp 1606821651
transform 1 0 19872 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 20792 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1606821651
transform 1 0 20608 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1606821651
transform 1 0 20884 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_219
timestamp 1606821651
transform 1 0 21252 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606821651
transform 1 0 2484 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3864 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 6716 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1606821651
transform 1 0 5336 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1606821651
transform 1 0 6532 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1606821651
transform 1 0 6808 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8372 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1606821651
transform 1 0 7912 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1606821651
transform 1 0 8280 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_95
timestamp 1606821651
transform 1 0 9844 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 12328 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_107
timestamp 1606821651
transform 1 0 10948 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_119
timestamp 1606821651
transform 1 0 12052 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13800 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_132
timestamp 1606821651
transform 1 0 13248 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15456 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1606821651
transform 1 0 17296 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 17940 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1606821651
transform 1 0 16928 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1606821651
transform 1 0 17572 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1606821651
transform 1 0 18032 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19228 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19964 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_196
timestamp 1606821651
transform 1 0 19136 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1606821651
transform 1 0 19780 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 20700 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_211
timestamp 1606821651
transform 1 0 20516 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_217
timestamp 1606821651
transform 1 0 21068 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606821651
transform 1 0 2484 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 3956 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1606821651
transform 1 0 3588 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_41
timestamp 1606821651
transform 1 0 4876 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_53
timestamp 1606821651
transform 1 0 5980 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8004 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1606821651
transform 1 0 7084 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1606821651
transform 1 0 7820 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1606821651
transform 1 0 10672 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 9568 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_84
timestamp 1606821651
transform 1 0 8832 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_102
timestamp 1606821651
transform 1 0 10488 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11960 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_107
timestamp 1606821651
transform 1 0 10948 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_115
timestamp 1606821651
transform 1 0 11684 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13524 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_track_0.prog_clk
timestamp 1606821651
transform 1 0 13156 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1606821651
transform 1 0 12788 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_134
timestamp 1606821651
transform 1 0 13432 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 15180 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1606821651
transform 1 0 14996 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1606821651
transform 1 0 15272 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_166
timestamp 1606821651
transform 1 0 16376 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16468 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_176
timestamp 1606821651
transform 1 0 17296 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 20240 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 19688 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18768 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1606821651
transform 1 0 18400 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1606821651
transform 1 0 19320 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_206
timestamp 1606821651
transform 1 0 20056 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 20792 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_212
timestamp 1606821651
transform 1 0 20608 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606821651
transform 1 0 20884 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606821651
transform 1 0 21252 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1564 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1606821651
transform 1 0 4232 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4784 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3220 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_21
timestamp 1606821651
transform 1 0 3036 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_37
timestamp 1606821651
transform 1 0 4508 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 6716 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1606821651
transform 1 0 6256 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_60
timestamp 1606821651
transform 1 0 6624 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1606821651
transform 1 0 6808 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_track_0.prog_clk
timestamp 1606821651
transform 1 0 7176 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_69
timestamp 1606821651
transform 1 0 7452 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_81
timestamp 1606821651
transform 1 0 8556 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606821651
transform 1 0 9660 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 12328 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606821651
transform 1 0 10764 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1606821651
transform 1 0 11868 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1606821651
transform 1 0 12236 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1606821651
transform 1 0 12420 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_135
timestamp 1606821651
transform 1 0 13524 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1606821651
transform 1 0 14628 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_159
timestamp 1606821651
transform 1 0 15732 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 17940 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_171
timestamp 1606821651
transform 1 0 16836 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1606821651
transform 1 0 18032 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 19964 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18952 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1606821651
transform 1 0 18768 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_200
timestamp 1606821651
transform 1 0 19504 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_204
timestamp 1606821651
transform 1 0 19872 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 20516 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1606821651
transform 1 0 20332 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1748 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 3956 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_23
timestamp 1606821651
transform 1 0 3220 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1606821651
transform 1 0 4048 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5704 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_44
timestamp 1606821651
transform 1 0 5152 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7360 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1606821651
transform 1 0 7176 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_77
timestamp 1606821651
transform 1 0 8188 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1606821651
transform 1 0 10120 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 9568 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_89
timestamp 1606821651
transform 1 0 9292 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1606821651
transform 1 0 9660 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1606821651
transform 1 0 10028 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_101
timestamp 1606821651
transform 1 0 10396 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11500 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1606821651
transform 1 0 13156 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14076 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1606821651
transform 1 0 12972 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_134
timestamp 1606821651
transform 1 0 13432 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_140
timestamp 1606821651
transform 1 0 13984 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15272 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 15180 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_150
timestamp 1606821651
transform 1 0 14904 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1606821651
transform 1 0 16100 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16560 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1606821651
transform 1 0 16468 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_177
timestamp 1606821651
transform 1 0 17388 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 20240 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18860 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_189
timestamp 1606821651
transform 1 0 18492 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_199
timestamp 1606821651
transform 1 0 19412 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1606821651
transform 1 0 20148 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 20792 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1606821651
transform 1 0 20608 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606821651
transform 1 0 20884 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606821651
transform 1 0 21252 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606821651
transform 1 0 2484 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1606821651
transform 1 0 2484 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1606821651
transform 1 0 2852 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3864 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 3956 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_27
timestamp 1606821651
transform 1 0 3588 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_36
timestamp 1606821651
transform 1 0 4416 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1606821651
transform 1 0 3772 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_41
timestamp 1606821651
transform 1 0 4876 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6532 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 6716 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_48
timestamp 1606821651
transform 1 0 5520 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1606821651
transform 1 0 6624 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_62
timestamp 1606821651
transform 1 0 6808 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_53
timestamp 1606821651
transform 1 0 5980 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1606821651
transform 1 0 7912 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8740 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1606821651
transform 1 0 7728 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1606821651
transform 1 0 8188 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_75
timestamp 1606821651
transform 1 0 8004 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10396 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9752 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 9568 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_99
timestamp 1606821651
transform 1 0 10212 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1606821651
transform 1 0 9384 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1606821651
transform 1 0 9660 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_103
timestamp 1606821651
transform 1 0 10580 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11776 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 12328 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1606821651
transform 1 0 11868 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1606821651
transform 1 0 12236 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_123
timestamp 1606821651
transform 1 0 12420 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_115
timestamp 1606821651
transform 1 0 11684 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1606821651
transform 1 0 12604 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12972 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12788 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_26_145
timestamp 1606821651
transform 1 0 14444 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_136
timestamp 1606821651
transform 1 0 13616 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1606821651
transform 1 0 14996 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15548 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 15180 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1606821651
transform 1 0 14720 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_152
timestamp 1606821651
transform 1 0 15088 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1606821651
transform 1 0 15272 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_166
timestamp 1606821651
transform 1 0 16376 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606821651
transform 1 0 18032 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16468 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18124 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 17940 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_173
timestamp 1606821651
transform 1 0 17020 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1606821651
transform 1 0 17756 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1606821651
transform 1 0 18308 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_183
timestamp 1606821651
transform 1 0 17940 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19228 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19412 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19964 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18676 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1606821651
transform 1 0 19228 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_205
timestamp 1606821651
transform 1 0 19964 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_194
timestamp 1606821651
transform 1 0 18952 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1606821651
transform 1 0 19780 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 20516 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 20792 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_211
timestamp 1606821651
transform 1 0 20516 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606821651
transform 1 0 20884 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606821651
transform 1 0 21252 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1472 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_20
timestamp 1606821651
transform 1 0 2944 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1606821651
transform 1 0 3312 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1606821651
transform 1 0 3588 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_39
timestamp 1606821651
transform 1 0 4692 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4968 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 6716 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1606821651
transform 1 0 6440 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1606821651
transform 1 0 6808 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1606821651
transform 1 0 7912 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1606821651
transform 1 0 9016 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1606821651
transform 1 0 10120 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 12328 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1606821651
transform 1 0 11224 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1606821651
transform 1 0 12420 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_135
timestamp 1606821651
transform 1 0 13524 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_147
timestamp 1606821651
transform 1 0 14628 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_159
timestamp 1606821651
transform 1 0 15732 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 17940 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1606821651
transform 1 0 16836 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1606821651
transform 1 0 18032 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 20240 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 19688 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_196
timestamp 1606821651
transform 1 0 19136 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1606821651
transform 1 0 20056 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 20792 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606821651
transform 1 0 20608 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_218
timestamp 1606821651
transform 1 0 21160 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606821651
transform 1 0 2484 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 3956 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1606821651
transform 1 0 3588 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1606821651
transform 1 0 4048 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5244 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_44
timestamp 1606821651
transform 1 0 5152 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_51
timestamp 1606821651
transform 1 0 5796 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8372 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7360 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_63
timestamp 1606821651
transform 1 0 6900 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_67
timestamp 1606821651
transform 1 0 7268 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_77
timestamp 1606821651
transform 1 0 8188 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 9568 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1606821651
transform 1 0 9200 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1606821651
transform 1 0 9660 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606821651
transform 1 0 10764 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_108
timestamp 1606821651
transform 1 0 11040 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_120
timestamp 1606821651
transform 1 0 12144 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13340 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_132
timestamp 1606821651
transform 1 0 13248 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_142
timestamp 1606821651
transform 1 0 14168 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 15180 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_150
timestamp 1606821651
transform 1 0 14904 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1606821651
transform 1 0 15272 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1606821651
transform 1 0 16376 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606821651
transform 1 0 16560 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606821651
transform 1 0 16836 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_183
timestamp 1606821651
transform 1 0 17940 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606821651
transform 1 0 19504 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1606821651
transform 1 0 19044 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1606821651
transform 1 0 19412 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_204
timestamp 1606821651
transform 1 0 19872 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 20792 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1606821651
transform 1 0 20608 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606821651
transform 1 0 20884 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606821651
transform 1 0 21252 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2392 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_11
timestamp 1606821651
transform 1 0 2116 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4784 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_30
timestamp 1606821651
transform 1 0 3864 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_38
timestamp 1606821651
transform 1 0 4600 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1606821651
transform 1 0 5796 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 6716 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 1606821651
transform 1 0 5612 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_54
timestamp 1606821651
transform 1 0 6072 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_60
timestamp 1606821651
transform 1 0 6624 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606821651
transform 1 0 8464 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1606821651
transform 1 0 8280 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_83
timestamp 1606821651
transform 1 0 8740 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10672 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9200 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_87
timestamp 1606821651
transform 1 0 9108 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1606821651
transform 1 0 10028 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1606821651
transform 1 0 10580 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 12328 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1606821651
transform 1 0 12144 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13432 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_132
timestamp 1606821651
transform 1 0 13248 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15088 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_150
timestamp 1606821651
transform 1 0 14904 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16744 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 17940 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1606821651
transform 1 0 16560 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1606821651
transform 1 0 17572 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19504 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_190
timestamp 1606821651
transform 1 0 18584 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1606821651
transform 1 0 19320 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_206
timestamp 1606821651
transform 1 0 20056 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 20516 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1606821651
transform 1 0 20424 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606821651
transform 1 0 2484 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 3956 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1606821651
transform 1 0 3588 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_48
timestamp 1606821651
transform 1 0 5520 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_60
timestamp 1606821651
transform 1 0 6624 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7728 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 9568 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1606821651
transform 1 0 9200 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12328 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1606821651
transform 1 0 11132 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606821651
transform 1 0 12144 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606821651
transform 1 0 13984 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1606821651
transform 1 0 13800 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_143
timestamp 1606821651
transform 1 0 14260 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 15180 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1606821651
transform 1 0 14996 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1606821651
transform 1 0 16100 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16928 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 17940 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_171
timestamp 1606821651
transform 1 0 16836 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1606821651
transform 1 0 17480 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1606821651
transform 1 0 17848 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 20240 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19504 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1606821651
transform 1 0 19044 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1606821651
transform 1 0 19412 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1606821651
transform 1 0 20056 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 20792 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1606821651
transform 1 0 20608 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606821651
transform 1 0 20884 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606821651
transform 1 0 21252 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606821651
transform 1 0 2484 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4600 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 3956 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606821651
transform 1 0 3588 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 6808 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_47
timestamp 1606821651
transform 1 0 5428 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1606821651
transform 1 0 6532 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 9660 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606821651
transform 1 0 9108 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606821651
transform 1 0 9752 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 12512 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606821651
transform 1 0 10856 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606821651
transform 1 0 11960 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606821651
transform 1 0 12604 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606821651
transform 1 0 13708 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 15364 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606821651
transform 1 0 14812 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606821651
transform 1 0 17664 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 18216 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606821651
transform 1 0 16560 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1606821651
transform 1 0 18032 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_187
timestamp 1606821651
transform 1 0 18308 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 18400 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19504 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1606821651
transform 1 0 18768 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1606821651
transform 1 0 20056 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 20516 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1606821651
transform 1 0 21068 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 1606821651
transform 1 0 20424 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 19984
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 5576 480 5696 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 17000 480 17120 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 22320 4080 22800 4200 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 22320 8568 22800 8688 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 22320 9112 22800 9232 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 22320 9520 22800 9640 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 22320 9928 22800 10048 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 22320 10472 22800 10592 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 22320 10880 22800 11000 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 22320 11424 22800 11544 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 22320 11832 22800 11952 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 22320 12240 22800 12360 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 22320 12784 22800 12904 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 22320 4488 22800 4608 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 22320 4896 22800 5016 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 22320 5440 22800 5560 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 22320 5848 22800 5968 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 22320 6392 22800 6512 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 22320 6800 22800 6920 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 22320 7208 22800 7328 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 22320 7752 22800 7872 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 22320 8160 22800 8280 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 22320 13192 22800 13312 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 22320 17816 22800 17936 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 22320 18224 22800 18344 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 22320 18632 22800 18752 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 22320 19176 22800 19296 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 22320 19584 22800 19704 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 22320 19992 22800 20112 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 22320 20536 22800 20656 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 22320 20944 22800 21064 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 22320 21352 22800 21472 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 22320 21896 22800 22016 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 22320 13600 22800 13720 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 22320 14144 22800 14264 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 22320 14552 22800 14672 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 22320 14960 22800 15080 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 22320 15504 22800 15624 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 22320 15912 22800 16032 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 22320 16320 22800 16440 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 22320 16864 22800 16984 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 22320 17272 22800 17392 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 846 22176 902 22656 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 6366 22176 6422 22656 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 6918 22176 6974 22656 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 7470 22176 7526 22656 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 8022 22176 8078 22656 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 8574 22176 8630 22656 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 9126 22176 9182 22656 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 9678 22176 9734 22656 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 10230 22176 10286 22656 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 10782 22176 10838 22656 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 11334 22176 11390 22656 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1398 22176 1454 22656 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 1950 22176 2006 22656 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2502 22176 2558 22656 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3054 22176 3110 22656 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 3606 22176 3662 22656 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4158 22176 4214 22656 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 4710 22176 4766 22656 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 5262 22176 5318 22656 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 5814 22176 5870 22656 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 11978 22176 12034 22656 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17498 22176 17554 22656 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 18050 22176 18106 22656 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18602 22176 18658 22656 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 19154 22176 19210 22656 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19706 22176 19762 22656 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 20258 22176 20314 22656 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20810 22176 20866 22656 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 21362 22176 21418 22656 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21914 22176 21970 22656 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 22466 22176 22522 22656 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 12530 22176 12586 22656 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 13082 22176 13138 22656 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 13634 22176 13690 22656 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 14186 22176 14242 22656 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 14738 22176 14794 22656 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 15290 22176 15346 22656 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 15842 22176 15898 22656 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16394 22176 16450 22656 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 16946 22176 17002 22656 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 22320 22304 22800 22424 6 prog_clk_0_E_in
port 82 nsew default input
rlabel metal3 s 22320 2176 22800 2296 6 right_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 22320 2720 22800 2840 6 right_bottom_grid_pin_13_
port 84 nsew default input
rlabel metal3 s 22320 3128 22800 3248 6 right_bottom_grid_pin_15_
port 85 nsew default input
rlabel metal3 s 22320 3536 22800 3656 6 right_bottom_grid_pin_17_
port 86 nsew default input
rlabel metal3 s 22320 0 22800 120 6 right_bottom_grid_pin_1_
port 87 nsew default input
rlabel metal3 s 22320 408 22800 528 6 right_bottom_grid_pin_3_
port 88 nsew default input
rlabel metal3 s 22320 816 22800 936 6 right_bottom_grid_pin_5_
port 89 nsew default input
rlabel metal3 s 22320 1360 22800 1480 6 right_bottom_grid_pin_7_
port 90 nsew default input
rlabel metal3 s 22320 1768 22800 1888 6 right_bottom_grid_pin_9_
port 91 nsew default input
rlabel metal2 s 294 22176 350 22656 6 top_left_grid_pin_1_
port 92 nsew default input
rlabel metal4 s 4376 1984 4696 20032 6 VPWR
port 93 nsew default input
rlabel metal4 s 7808 1984 8128 20032 6 VGND
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22656
<< end >>
