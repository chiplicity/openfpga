magic
tech EFS8A
magscale 1 2
timestamp 1602873728
<< locali >>
rect 4537 25347 4571 25449
rect 12357 25279 12391 25449
rect 15485 25347 15519 25449
rect 12943 25313 12978 25347
rect 13955 25313 13990 25347
rect 15485 25313 15646 25347
rect 16623 25313 16658 25347
rect 18279 25313 18406 25347
rect 19383 25313 19418 25347
rect 15887 24701 16014 24735
rect 16497 24225 16658 24259
rect 16497 24055 16531 24225
rect 17267 23137 17302 23171
rect 6469 22491 6503 22593
rect 13271 22423 13305 22491
rect 13271 22389 13277 22423
rect 2973 20247 3007 20417
rect 14933 19227 14967 19465
rect 17693 19295 17727 19465
rect 13363 19159 13397 19227
rect 13363 19125 13369 19159
rect 5267 18071 5301 18139
rect 13369 18071 13403 18173
rect 5267 18037 5273 18071
rect 13369 18037 13495 18071
rect 16767 17833 16773 17867
rect 16767 17765 16801 17833
rect 13277 17527 13311 17697
rect 12725 17119 12759 17289
rect 16991 17085 17026 17119
rect 6187 16745 6193 16779
rect 6187 16677 6221 16745
rect 8401 15895 8435 16065
rect 16991 14433 17026 14467
rect 5359 12631 5393 12699
rect 5359 12597 5365 12631
rect 4169 10557 4261 10591
rect 4169 10455 4203 10557
rect 3571 9673 3617 9707
rect 3157 9503 3191 9605
rect 2559 8585 2697 8619
rect 1547 8517 1685 8551
rect 1443 7905 1478 7939
rect 1443 6817 1478 6851
rect 1547 3689 1593 3723
<< viali >>
rect 4261 25449 4295 25483
rect 4537 25449 4571 25483
rect 4721 25449 4755 25483
rect 12357 25449 12391 25483
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 4537 25313 4571 25347
rect 5825 25313 5859 25347
rect 8309 25313 8343 25347
rect 9873 25313 9907 25347
rect 11412 25313 11446 25347
rect 15485 25449 15519 25483
rect 18475 25381 18509 25415
rect 12909 25313 12943 25347
rect 13921 25313 13955 25347
rect 16589 25313 16623 25347
rect 18245 25313 18279 25347
rect 19349 25313 19383 25347
rect 1409 25245 1443 25279
rect 2421 25245 2455 25279
rect 5181 25245 5215 25279
rect 7757 25245 7791 25279
rect 12357 25245 12391 25279
rect 16727 25177 16761 25211
rect 10057 25109 10091 25143
rect 11483 25109 11517 25143
rect 13047 25109 13081 25143
rect 14059 25109 14093 25143
rect 15715 25109 15749 25143
rect 19487 25109 19521 25143
rect 5089 24905 5123 24939
rect 9873 24905 9907 24939
rect 11805 24905 11839 24939
rect 13461 24905 13495 24939
rect 14473 24905 14507 24939
rect 14841 24905 14875 24939
rect 15669 24905 15703 24939
rect 16589 24905 16623 24939
rect 18521 24905 18555 24939
rect 1961 24769 1995 24803
rect 4721 24769 4755 24803
rect 19211 24769 19245 24803
rect 3525 24701 3559 24735
rect 4261 24701 4295 24735
rect 6653 24701 6687 24735
rect 6929 24701 6963 24735
rect 8493 24701 8527 24735
rect 8677 24701 8711 24735
rect 10701 24701 10735 24735
rect 10885 24701 10919 24735
rect 12265 24701 12299 24735
rect 12541 24701 12575 24735
rect 14064 24701 14098 24735
rect 15853 24701 15887 24735
rect 18096 24701 18130 24735
rect 18889 24701 18923 24735
rect 19108 24701 19142 24735
rect 19901 24701 19935 24735
rect 1777 24633 1811 24667
rect 2053 24633 2087 24667
rect 2605 24633 2639 24667
rect 5273 24633 5307 24667
rect 5365 24633 5399 24667
rect 5917 24633 5951 24667
rect 6837 24633 6871 24667
rect 10793 24633 10827 24667
rect 12449 24633 12483 24667
rect 14151 24633 14185 24667
rect 19533 24633 19567 24667
rect 2881 24565 2915 24599
rect 3893 24565 3927 24599
rect 7941 24565 7975 24599
rect 8861 24565 8895 24599
rect 16083 24565 16117 24599
rect 16957 24565 16991 24599
rect 18199 24565 18233 24599
rect 1961 24361 1995 24395
rect 11897 24361 11931 24395
rect 18521 24361 18555 24395
rect 2329 24293 2363 24327
rect 4261 24293 4295 24327
rect 5825 24293 5859 24327
rect 6377 24293 6411 24327
rect 8217 24293 8251 24327
rect 10149 24293 10183 24327
rect 12173 24293 12207 24327
rect 12265 24293 12299 24327
rect 14105 24225 14139 24259
rect 15460 24225 15494 24259
rect 16727 24225 16761 24259
rect 18337 24225 18371 24259
rect 19508 24225 19542 24259
rect 2237 24157 2271 24191
rect 2605 24157 2639 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 5733 24157 5767 24191
rect 8125 24157 8159 24191
rect 8401 24157 8435 24191
rect 10057 24157 10091 24191
rect 10701 24157 10735 24191
rect 12817 24157 12851 24191
rect 13093 24157 13127 24191
rect 14381 24157 14415 24191
rect 3157 24089 3191 24123
rect 7941 24089 7975 24123
rect 19579 24089 19613 24123
rect 5273 24021 5307 24055
rect 15531 24021 15565 24055
rect 15945 24021 15979 24055
rect 16497 24021 16531 24055
rect 19257 24021 19291 24055
rect 2605 23817 2639 23851
rect 3801 23817 3835 23851
rect 5641 23817 5675 23851
rect 6377 23817 6411 23851
rect 8769 23817 8803 23851
rect 9873 23817 9907 23851
rect 10701 23817 10735 23851
rect 12173 23817 12207 23851
rect 14105 23817 14139 23851
rect 14473 23817 14507 23851
rect 15761 23817 15795 23851
rect 17049 23817 17083 23851
rect 19073 23817 19107 23851
rect 19441 23817 19475 23851
rect 24961 23817 24995 23851
rect 18337 23749 18371 23783
rect 23857 23749 23891 23783
rect 1685 23681 1719 23715
rect 2145 23681 2179 23715
rect 3433 23681 3467 23715
rect 4629 23681 4663 23715
rect 8033 23681 8067 23715
rect 9229 23681 9263 23715
rect 13185 23681 13219 23715
rect 13829 23681 13863 23715
rect 14749 23681 14783 23715
rect 15025 23681 15059 23715
rect 16589 23681 16623 23715
rect 19809 23681 19843 23715
rect 5445 23613 5479 23647
rect 16865 23613 16899 23647
rect 17417 23613 17451 23647
rect 18153 23613 18187 23647
rect 18705 23613 18739 23647
rect 19257 23613 19291 23647
rect 20396 23613 20430 23647
rect 20821 23613 20855 23647
rect 21424 23613 21458 23647
rect 21833 23613 21867 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 24777 23613 24811 23647
rect 1777 23545 1811 23579
rect 2973 23545 3007 23579
rect 3985 23545 4019 23579
rect 4077 23545 4111 23579
rect 7389 23545 7423 23579
rect 7481 23545 7515 23579
rect 8401 23545 8435 23579
rect 8953 23545 8987 23579
rect 9045 23545 9079 23579
rect 10333 23545 10367 23579
rect 10885 23545 10919 23579
rect 10977 23545 11011 23579
rect 11529 23545 11563 23579
rect 13277 23545 13311 23579
rect 14841 23545 14875 23579
rect 21511 23545 21545 23579
rect 25329 23545 25363 23579
rect 4997 23477 5031 23511
rect 5365 23477 5399 23511
rect 6101 23477 6135 23511
rect 7205 23477 7239 23511
rect 13001 23477 13035 23511
rect 20499 23477 20533 23511
rect 2237 23273 2271 23307
rect 4261 23273 4295 23307
rect 14749 23273 14783 23307
rect 17371 23273 17405 23307
rect 18383 23273 18417 23307
rect 5911 23205 5945 23239
rect 8217 23205 8251 23239
rect 8769 23205 8803 23239
rect 10609 23205 10643 23239
rect 11161 23205 11195 23239
rect 12173 23205 12207 23239
rect 12725 23205 12759 23239
rect 13829 23205 13863 23239
rect 2605 23137 2639 23171
rect 4077 23137 4111 23171
rect 15669 23137 15703 23171
rect 17233 23137 17267 23171
rect 18280 23137 18314 23171
rect 19324 23137 19358 23171
rect 5549 23069 5583 23103
rect 8125 23069 8159 23103
rect 10517 23069 10551 23103
rect 11437 23069 11471 23103
rect 12081 23069 12115 23103
rect 13737 23069 13771 23103
rect 15301 23069 15335 23103
rect 6837 23001 6871 23035
rect 14289 23001 14323 23035
rect 1685 22933 1719 22967
rect 3065 22933 3099 22967
rect 5089 22933 5123 22967
rect 6469 22933 6503 22967
rect 7389 22933 7423 22967
rect 7941 22933 7975 22967
rect 9965 22933 9999 22967
rect 13001 22933 13035 22967
rect 16405 22933 16439 22967
rect 19395 22933 19429 22967
rect 2973 22729 3007 22763
rect 5917 22729 5951 22763
rect 7941 22729 7975 22763
rect 9321 22729 9355 22763
rect 9597 22729 9631 22763
rect 10057 22729 10091 22763
rect 12081 22729 12115 22763
rect 13829 22729 13863 22763
rect 14197 22729 14231 22763
rect 15669 22729 15703 22763
rect 17325 22729 17359 22763
rect 18889 22729 18923 22763
rect 19211 22729 19245 22763
rect 19901 22729 19935 22763
rect 11529 22661 11563 22695
rect 1961 22593 1995 22627
rect 2329 22593 2363 22627
rect 6469 22593 6503 22627
rect 10241 22593 10275 22627
rect 10701 22593 10735 22627
rect 15025 22593 15059 22627
rect 16681 22593 16715 22627
rect 20085 22593 20119 22627
rect 3341 22525 3375 22559
rect 3709 22525 3743 22559
rect 3893 22525 3927 22559
rect 4169 22525 4203 22559
rect 4997 22525 5031 22559
rect 6837 22525 6871 22559
rect 7297 22525 7331 22559
rect 8401 22525 8435 22559
rect 12909 22525 12943 22559
rect 18128 22525 18162 22559
rect 18521 22525 18555 22559
rect 19140 22525 19174 22559
rect 1777 22457 1811 22491
rect 2053 22457 2087 22491
rect 5359 22457 5393 22491
rect 6469 22457 6503 22491
rect 6561 22457 6595 22491
rect 8309 22457 8343 22491
rect 8763 22457 8797 22491
rect 10333 22457 10367 22491
rect 14749 22457 14783 22491
rect 14841 22457 14875 22491
rect 16405 22457 16439 22491
rect 16497 22457 16531 22491
rect 4537 22389 4571 22423
rect 4905 22389 4939 22423
rect 6285 22389 6319 22423
rect 6929 22389 6963 22423
rect 11253 22389 11287 22423
rect 12817 22389 12851 22423
rect 13277 22389 13311 22423
rect 14565 22389 14599 22423
rect 16221 22389 16255 22423
rect 18199 22389 18233 22423
rect 19533 22389 19567 22423
rect 2789 22185 2823 22219
rect 5733 22185 5767 22219
rect 6837 22185 6871 22219
rect 8769 22185 8803 22219
rect 11253 22185 11287 22219
rect 13001 22185 13035 22219
rect 13737 22185 13771 22219
rect 14749 22185 14783 22219
rect 15485 22185 15519 22219
rect 22661 22185 22695 22219
rect 1685 22117 1719 22151
rect 5175 22117 5209 22151
rect 8211 22117 8245 22151
rect 10695 22117 10729 22151
rect 12443 22117 12477 22151
rect 15761 22117 15795 22151
rect 15853 22117 15887 22151
rect 16405 22117 16439 22151
rect 2329 22049 2363 22083
rect 11897 22049 11931 22083
rect 14264 22049 14298 22083
rect 17268 22049 17302 22083
rect 18312 22049 18346 22083
rect 19324 22049 19358 22083
rect 21373 22049 21407 22083
rect 22477 22049 22511 22083
rect 4813 21981 4847 22015
rect 7849 21981 7883 22015
rect 10333 21981 10367 22015
rect 12081 21981 12115 22015
rect 13277 21913 13311 21947
rect 21557 21913 21591 21947
rect 3525 21845 3559 21879
rect 6009 21845 6043 21879
rect 9045 21845 9079 21879
rect 10149 21845 10183 21879
rect 14335 21845 14369 21879
rect 17371 21845 17405 21879
rect 18383 21845 18417 21879
rect 19395 21845 19429 21879
rect 3893 21641 3927 21675
rect 6193 21641 6227 21675
rect 7941 21641 7975 21675
rect 9919 21641 9953 21675
rect 10425 21641 10459 21675
rect 12173 21641 12207 21675
rect 12817 21641 12851 21675
rect 13829 21641 13863 21675
rect 16681 21641 16715 21675
rect 17417 21641 17451 21675
rect 5917 21573 5951 21607
rect 9689 21573 9723 21607
rect 14105 21573 14139 21607
rect 19211 21573 19245 21607
rect 22477 21573 22511 21607
rect 6837 21505 6871 21539
rect 18199 21505 18233 21539
rect 21373 21505 21407 21539
rect 3617 21437 3651 21471
rect 3709 21437 3743 21471
rect 4997 21437 5031 21471
rect 6561 21437 6595 21471
rect 8401 21437 8435 21471
rect 8677 21437 8711 21471
rect 9848 21437 9882 21471
rect 10885 21437 10919 21471
rect 11253 21437 11287 21471
rect 12909 21437 12943 21471
rect 14657 21437 14691 21471
rect 15577 21437 15611 21471
rect 15945 21437 15979 21471
rect 16313 21437 16347 21471
rect 16497 21437 16531 21471
rect 18112 21437 18146 21471
rect 19108 21437 19142 21471
rect 19901 21437 19935 21471
rect 1685 21369 1719 21403
rect 2237 21369 2271 21403
rect 2329 21369 2363 21403
rect 2881 21369 2915 21403
rect 4537 21369 4571 21403
rect 4905 21369 4939 21403
rect 5318 21369 5352 21403
rect 7573 21369 7607 21403
rect 9321 21369 9355 21403
rect 11529 21369 11563 21403
rect 13230 21369 13264 21403
rect 14473 21369 14507 21403
rect 14978 21369 15012 21403
rect 18889 21369 18923 21403
rect 2053 21301 2087 21335
rect 8309 21301 8343 21335
rect 18521 21301 18555 21335
rect 19533 21301 19567 21335
rect 1777 21097 1811 21131
rect 2513 21097 2547 21131
rect 4261 21097 4295 21131
rect 5641 21097 5675 21131
rect 7941 21097 7975 21131
rect 10609 21097 10643 21131
rect 10977 21097 11011 21131
rect 13185 21097 13219 21131
rect 8769 21029 8803 21063
rect 10051 21029 10085 21063
rect 12265 21029 12299 21063
rect 17325 21029 17359 21063
rect 2881 20961 2915 20995
rect 4077 20961 4111 20995
rect 5825 20961 5859 20995
rect 6101 20961 6135 20995
rect 6377 20961 6411 20995
rect 8309 20961 8343 20995
rect 8493 20961 8527 20995
rect 11805 20961 11839 20995
rect 11989 20961 12023 20995
rect 12909 20961 12943 20995
rect 13369 20961 13403 20995
rect 13553 20961 13587 20995
rect 15485 20961 15519 20995
rect 19073 20961 19107 20995
rect 5457 20893 5491 20927
rect 9689 20893 9723 20927
rect 15301 20893 15335 20927
rect 17233 20893 17267 20927
rect 18705 20893 18739 20927
rect 17785 20825 17819 20859
rect 4905 20757 4939 20791
rect 6929 20757 6963 20791
rect 9505 20757 9539 20791
rect 11253 20757 11287 20791
rect 12633 20757 12667 20791
rect 14657 20757 14691 20791
rect 16497 20757 16531 20791
rect 18153 20757 18187 20791
rect 3893 20553 3927 20587
rect 5917 20553 5951 20587
rect 6285 20553 6319 20587
rect 10425 20553 10459 20587
rect 14381 20553 14415 20587
rect 15485 20553 15519 20587
rect 17509 20553 17543 20587
rect 19073 20553 19107 20587
rect 7757 20485 7791 20519
rect 9321 20485 9355 20519
rect 2237 20417 2271 20451
rect 2881 20417 2915 20451
rect 2973 20417 3007 20451
rect 6561 20417 6595 20451
rect 10149 20417 10183 20451
rect 11345 20417 11379 20451
rect 13185 20417 13219 20451
rect 14565 20417 14599 20451
rect 14841 20417 14875 20451
rect 16486 20417 16520 20451
rect 18153 20417 18187 20451
rect 19625 20417 19659 20451
rect 20637 20417 20671 20451
rect 1685 20281 1719 20315
rect 2053 20281 2087 20315
rect 2329 20281 2363 20315
rect 3709 20349 3743 20383
rect 4721 20349 4755 20383
rect 5089 20349 5123 20383
rect 5641 20349 5675 20383
rect 5825 20349 5859 20383
rect 6837 20349 6871 20383
rect 8125 20349 8159 20383
rect 9413 20349 9447 20383
rect 9873 20349 9907 20383
rect 12449 20349 12483 20383
rect 12909 20349 12943 20383
rect 13829 20349 13863 20383
rect 3525 20281 3559 20315
rect 4353 20281 4387 20315
rect 7158 20281 7192 20315
rect 8953 20281 8987 20315
rect 14657 20281 14691 20315
rect 16313 20281 16347 20315
rect 16589 20281 16623 20315
rect 17141 20281 17175 20315
rect 18245 20281 18279 20315
rect 18797 20281 18831 20315
rect 2973 20213 3007 20247
rect 3157 20213 3191 20247
rect 8493 20213 8527 20247
rect 11161 20213 11195 20247
rect 11805 20213 11839 20247
rect 12173 20213 12207 20247
rect 13553 20213 13587 20247
rect 17877 20213 17911 20247
rect 2973 20009 3007 20043
rect 5917 20009 5951 20043
rect 9781 20009 9815 20043
rect 14657 20009 14691 20043
rect 16957 20009 16991 20043
rect 24593 20009 24627 20043
rect 2513 19941 2547 19975
rect 4261 19941 4295 19975
rect 4813 19941 4847 19975
rect 5641 19941 5675 19975
rect 7941 19941 7975 19975
rect 13829 19941 13863 19975
rect 16358 19941 16392 19975
rect 17969 19941 18003 19975
rect 18797 19941 18831 19975
rect 2053 19873 2087 19907
rect 6101 19873 6135 19907
rect 6653 19873 6687 19907
rect 8309 19873 8343 19907
rect 8585 19873 8619 19907
rect 9781 19873 9815 19907
rect 10149 19873 10183 19907
rect 11805 19873 11839 19907
rect 12173 19873 12207 19907
rect 19349 19873 19383 19907
rect 24409 19873 24443 19907
rect 2145 19805 2179 19839
rect 4169 19805 4203 19839
rect 6745 19805 6779 19839
rect 8677 19805 8711 19839
rect 12449 19805 12483 19839
rect 13553 19805 13587 19839
rect 13737 19805 13771 19839
rect 14381 19805 14415 19839
rect 16037 19805 16071 19839
rect 17877 19805 17911 19839
rect 18337 19805 18371 19839
rect 3801 19737 3835 19771
rect 17601 19737 17635 19771
rect 3433 19669 3467 19703
rect 5181 19669 5215 19703
rect 7297 19669 7331 19703
rect 9413 19669 9447 19703
rect 13001 19669 13035 19703
rect 17233 19669 17267 19703
rect 19533 19669 19567 19703
rect 4169 19465 4203 19499
rect 8309 19465 8343 19499
rect 9459 19465 9493 19499
rect 9965 19465 9999 19499
rect 10701 19465 10735 19499
rect 12173 19465 12207 19499
rect 12817 19465 12851 19499
rect 13921 19465 13955 19499
rect 14933 19465 14967 19499
rect 15117 19465 15151 19499
rect 16129 19465 16163 19499
rect 17693 19465 17727 19499
rect 17785 19465 17819 19499
rect 19349 19465 19383 19499
rect 2605 19397 2639 19431
rect 3709 19397 3743 19431
rect 9597 19397 9631 19431
rect 10425 19397 10459 19431
rect 11805 19397 11839 19431
rect 1593 19329 1627 19363
rect 3157 19329 3191 19363
rect 4537 19329 4571 19363
rect 9689 19329 9723 19363
rect 13001 19329 13035 19363
rect 4997 19261 5031 19295
rect 5089 19261 5123 19295
rect 5641 19261 5675 19295
rect 6193 19261 6227 19295
rect 6653 19261 6687 19295
rect 7113 19261 7147 19295
rect 7665 19261 7699 19295
rect 7849 19261 7883 19295
rect 10885 19261 10919 19295
rect 14657 19261 14691 19295
rect 16773 19329 16807 19363
rect 18061 19329 18095 19363
rect 19763 19329 19797 19363
rect 24409 19329 24443 19363
rect 15209 19261 15243 19295
rect 16957 19261 16991 19295
rect 17417 19261 17451 19295
rect 17693 19261 17727 19295
rect 18153 19261 18187 19295
rect 19676 19261 19710 19295
rect 20085 19261 20119 19295
rect 1685 19193 1719 19227
rect 2237 19193 2271 19227
rect 3249 19193 3283 19227
rect 8861 19193 8895 19227
rect 9321 19193 9355 19227
rect 14933 19193 14967 19227
rect 15571 19193 15605 19227
rect 16405 19193 16439 19227
rect 2973 19125 3007 19159
rect 5181 19125 5215 19159
rect 6929 19125 6963 19159
rect 9229 19125 9263 19159
rect 13369 19125 13403 19159
rect 14289 19125 14323 19159
rect 17141 19125 17175 19159
rect 2053 18921 2087 18955
rect 5089 18921 5123 18955
rect 10333 18921 10367 18955
rect 16957 18921 16991 18955
rect 2513 18853 2547 18887
rect 3065 18853 3099 18887
rect 4261 18853 4295 18887
rect 6187 18853 6221 18887
rect 7941 18853 7975 18887
rect 8033 18853 8067 18887
rect 12903 18853 12937 18887
rect 15485 18853 15519 18887
rect 18429 18853 18463 18887
rect 5825 18785 5859 18819
rect 7573 18785 7607 18819
rect 8180 18785 8214 18819
rect 8769 18785 8803 18819
rect 9689 18785 9723 18819
rect 11069 18785 11103 18819
rect 11253 18785 11287 18819
rect 13461 18785 13495 18819
rect 16865 18785 16899 18819
rect 17325 18785 17359 18819
rect 19073 18785 19107 18819
rect 2421 18717 2455 18751
rect 3433 18717 3467 18751
rect 4169 18717 4203 18751
rect 4445 18717 4479 18751
rect 5733 18717 5767 18751
rect 8401 18717 8435 18751
rect 10057 18717 10091 18751
rect 12541 18717 12575 18751
rect 13737 18717 13771 18751
rect 15393 18717 15427 18751
rect 15669 18717 15703 18751
rect 6745 18649 6779 18683
rect 11437 18649 11471 18683
rect 12357 18649 12391 18683
rect 1593 18581 1627 18615
rect 7021 18581 7055 18615
rect 8309 18581 8343 18615
rect 9321 18581 9355 18615
rect 9827 18581 9861 18615
rect 9965 18581 9999 18615
rect 10793 18581 10827 18615
rect 11805 18581 11839 18615
rect 14381 18581 14415 18615
rect 18153 18581 18187 18615
rect 2421 18377 2455 18411
rect 2881 18377 2915 18411
rect 4169 18377 4203 18411
rect 5825 18377 5859 18411
rect 10498 18377 10532 18411
rect 10977 18377 11011 18411
rect 12909 18377 12943 18411
rect 15393 18377 15427 18411
rect 16865 18377 16899 18411
rect 17325 18377 17359 18411
rect 19073 18377 19107 18411
rect 4721 18309 4755 18343
rect 6193 18309 6227 18343
rect 10609 18309 10643 18343
rect 12587 18309 12621 18343
rect 12725 18309 12759 18343
rect 18705 18309 18739 18343
rect 3157 18241 3191 18275
rect 3433 18241 3467 18275
rect 8125 18241 8159 18275
rect 10701 18241 10735 18275
rect 12817 18241 12851 18275
rect 14381 18241 14415 18275
rect 14841 18241 14875 18275
rect 15945 18241 15979 18275
rect 18153 18241 18187 18275
rect 19625 18241 19659 18275
rect 4905 18173 4939 18207
rect 6837 18173 6871 18207
rect 7297 18173 7331 18207
rect 8861 18173 8895 18207
rect 11805 18173 11839 18207
rect 13369 18173 13403 18207
rect 1501 18105 1535 18139
rect 1593 18105 1627 18139
rect 2145 18105 2179 18139
rect 3249 18105 3283 18139
rect 9505 18105 9539 18139
rect 10333 18105 10367 18139
rect 11437 18105 11471 18139
rect 12449 18105 12483 18139
rect 14197 18105 14231 18139
rect 14473 18105 14507 18139
rect 16037 18105 16071 18139
rect 16589 18105 16623 18139
rect 17877 18105 17911 18139
rect 18245 18105 18279 18139
rect 5273 18037 5307 18071
rect 6561 18037 6595 18071
rect 6929 18037 6963 18071
rect 8585 18037 8619 18071
rect 9873 18037 9907 18071
rect 10149 18037 10183 18071
rect 12265 18037 12299 18071
rect 13553 18037 13587 18071
rect 15761 18037 15795 18071
rect 3157 17833 3191 17867
rect 4721 17833 4755 17867
rect 5733 17833 5767 17867
rect 6009 17833 6043 17867
rect 8493 17833 8527 17867
rect 13093 17833 13127 17867
rect 13461 17833 13495 17867
rect 13737 17833 13771 17867
rect 15117 17833 15151 17867
rect 15853 17833 15887 17867
rect 16773 17833 16807 17867
rect 2145 17765 2179 17799
rect 5175 17765 5209 17799
rect 10241 17765 10275 17799
rect 10977 17765 11011 17799
rect 18337 17765 18371 17799
rect 7481 17697 7515 17731
rect 10388 17697 10422 17731
rect 12081 17697 12115 17731
rect 12541 17697 12575 17731
rect 13277 17697 13311 17731
rect 13645 17697 13679 17731
rect 14105 17697 14139 17731
rect 15301 17697 15335 17731
rect 19717 17697 19751 17731
rect 2053 17629 2087 17663
rect 2697 17629 2731 17663
rect 4813 17629 4847 17663
rect 8125 17629 8159 17663
rect 10609 17629 10643 17663
rect 12817 17629 12851 17663
rect 6929 17561 6963 17595
rect 10517 17561 10551 17595
rect 11253 17561 11287 17595
rect 11621 17561 11655 17595
rect 16405 17629 16439 17663
rect 18245 17629 18279 17663
rect 18705 17629 18739 17663
rect 15485 17561 15519 17595
rect 19901 17561 19935 17595
rect 1685 17493 1719 17527
rect 3525 17493 3559 17527
rect 4261 17493 4295 17527
rect 8769 17493 8803 17527
rect 9505 17493 9539 17527
rect 9965 17493 9999 17527
rect 13277 17493 13311 17527
rect 17325 17493 17359 17527
rect 1685 17289 1719 17323
rect 2513 17289 2547 17323
rect 4169 17289 4203 17323
rect 4905 17289 4939 17323
rect 6561 17289 6595 17323
rect 8953 17289 8987 17323
rect 9965 17289 9999 17323
rect 10885 17289 10919 17323
rect 11253 17289 11287 17323
rect 12725 17289 12759 17323
rect 13001 17289 13035 17323
rect 14565 17289 14599 17323
rect 16773 17289 16807 17323
rect 18337 17289 18371 17323
rect 19073 17289 19107 17323
rect 3617 17221 3651 17255
rect 7757 17221 7791 17255
rect 8815 17221 8849 17255
rect 9137 17221 9171 17255
rect 11989 17221 12023 17255
rect 3065 17153 3099 17187
rect 4537 17153 4571 17187
rect 9045 17153 9079 17187
rect 10977 17153 11011 17187
rect 11713 17153 11747 17187
rect 14933 17221 14967 17255
rect 16037 17221 16071 17255
rect 2053 17085 2087 17119
rect 5457 17085 5491 17119
rect 5641 17085 5675 17119
rect 5917 17085 5951 17119
rect 6285 17085 6319 17119
rect 6837 17085 6871 17119
rect 8677 17085 8711 17119
rect 10756 17085 10790 17119
rect 12449 17085 12483 17119
rect 12725 17085 12759 17119
rect 13645 17085 13679 17119
rect 16957 17085 16991 17119
rect 17509 17085 17543 17119
rect 17877 17085 17911 17119
rect 18153 17085 18187 17119
rect 3157 17017 3191 17051
rect 7158 17017 7192 17051
rect 8585 17017 8619 17051
rect 10241 17017 10275 17051
rect 10609 17017 10643 17051
rect 13966 17017 14000 17051
rect 15485 17017 15519 17051
rect 15577 17017 15611 17051
rect 2881 16949 2915 16983
rect 8033 16949 8067 16983
rect 12633 16949 12667 16983
rect 13461 16949 13495 16983
rect 15301 16949 15335 16983
rect 16405 16949 16439 16983
rect 17095 16949 17129 16983
rect 19717 16949 19751 16983
rect 3065 16745 3099 16779
rect 6193 16745 6227 16779
rect 6745 16745 6779 16779
rect 7665 16745 7699 16779
rect 10333 16745 10367 16779
rect 11161 16745 11195 16779
rect 13001 16745 13035 16779
rect 13553 16745 13587 16779
rect 14657 16745 14691 16779
rect 2145 16677 2179 16711
rect 4997 16677 5031 16711
rect 7113 16677 7147 16711
rect 9137 16677 9171 16711
rect 10793 16677 10827 16711
rect 13737 16677 13771 16711
rect 13829 16677 13863 16711
rect 16773 16677 16807 16711
rect 18153 16677 18187 16711
rect 4261 16609 4295 16643
rect 5825 16609 5859 16643
rect 7573 16609 7607 16643
rect 8033 16609 8067 16643
rect 9689 16609 9723 16643
rect 11989 16609 12023 16643
rect 12449 16609 12483 16643
rect 15301 16609 15335 16643
rect 18797 16609 18831 16643
rect 2053 16541 2087 16575
rect 2513 16541 2547 16575
rect 3709 16541 3743 16575
rect 4408 16541 4442 16575
rect 4629 16541 4663 16575
rect 10057 16541 10091 16575
rect 12725 16541 12759 16575
rect 14381 16541 14415 16575
rect 15761 16541 15795 16575
rect 16681 16541 16715 16575
rect 16957 16541 16991 16575
rect 17601 16541 17635 16575
rect 11805 16473 11839 16507
rect 1777 16405 1811 16439
rect 3433 16405 3467 16439
rect 4537 16405 4571 16439
rect 5365 16405 5399 16439
rect 5641 16405 5675 16439
rect 7481 16405 7515 16439
rect 8769 16405 8803 16439
rect 9827 16405 9861 16439
rect 9965 16405 9999 16439
rect 11529 16405 11563 16439
rect 15485 16405 15519 16439
rect 4353 16201 4387 16235
rect 8309 16201 8343 16235
rect 10517 16201 10551 16235
rect 15945 16201 15979 16235
rect 17049 16201 17083 16235
rect 18245 16201 18279 16235
rect 18889 16201 18923 16235
rect 6193 16133 6227 16167
rect 7849 16133 7883 16167
rect 9045 16133 9079 16167
rect 13921 16133 13955 16167
rect 15669 16133 15703 16167
rect 3433 16065 3467 16099
rect 3709 16065 3743 16099
rect 4813 16065 4847 16099
rect 8401 16065 8435 16099
rect 8916 16065 8950 16099
rect 9137 16065 9171 16099
rect 9229 16065 9263 16099
rect 13001 16065 13035 16099
rect 14289 16065 14323 16099
rect 16497 16065 16531 16099
rect 17325 16065 17359 16099
rect 1777 15997 1811 16031
rect 5457 15997 5491 16031
rect 5733 15997 5767 16031
rect 7113 15997 7147 16031
rect 7389 15997 7423 16031
rect 1685 15929 1719 15963
rect 3525 15929 3559 15963
rect 5917 15929 5951 15963
rect 6653 15929 6687 15963
rect 10793 15997 10827 16031
rect 11253 15997 11287 16031
rect 11529 15997 11563 16031
rect 14749 15997 14783 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 8585 15929 8619 15963
rect 8769 15929 8803 15963
rect 9781 15929 9815 15963
rect 11989 15929 12023 15963
rect 13322 15929 13356 15963
rect 15070 15929 15104 15963
rect 2789 15861 2823 15895
rect 3157 15861 3191 15895
rect 6929 15861 6963 15895
rect 8401 15861 8435 15895
rect 10241 15861 10275 15895
rect 12909 15861 12943 15895
rect 14565 15861 14599 15895
rect 1409 15657 1443 15691
rect 4629 15657 4663 15691
rect 6469 15657 6503 15691
rect 7941 15657 7975 15691
rect 8217 15657 8251 15691
rect 8585 15657 8619 15691
rect 13093 15657 13127 15691
rect 13553 15657 13587 15691
rect 14749 15657 14783 15691
rect 2605 15589 2639 15623
rect 5267 15589 5301 15623
rect 6193 15589 6227 15623
rect 6974 15589 7008 15623
rect 8953 15589 8987 15623
rect 9413 15589 9447 15623
rect 9689 15589 9723 15623
rect 12817 15589 12851 15623
rect 13829 15589 13863 15623
rect 16129 15589 16163 15623
rect 16681 15589 16715 15623
rect 17509 15589 17543 15623
rect 4353 15521 4387 15555
rect 6653 15521 6687 15555
rect 8401 15521 8435 15555
rect 10793 15521 10827 15555
rect 12081 15521 12115 15555
rect 12541 15521 12575 15555
rect 17601 15521 17635 15555
rect 2513 15453 2547 15487
rect 2881 15453 2915 15487
rect 4905 15453 4939 15487
rect 10057 15453 10091 15487
rect 10425 15453 10459 15487
rect 13737 15453 13771 15487
rect 14381 15453 14415 15487
rect 16037 15453 16071 15487
rect 7573 15385 7607 15419
rect 1961 15317 1995 15351
rect 2329 15317 2363 15351
rect 5825 15317 5859 15351
rect 9827 15317 9861 15351
rect 9965 15317 9999 15351
rect 11253 15317 11287 15351
rect 11897 15317 11931 15351
rect 1593 15113 1627 15147
rect 5641 15113 5675 15147
rect 6653 15113 6687 15147
rect 7941 15113 7975 15147
rect 8309 15113 8343 15147
rect 10517 15113 10551 15147
rect 16313 15113 16347 15147
rect 17601 15113 17635 15147
rect 2145 15045 2179 15079
rect 5273 15045 5307 15079
rect 8907 15045 8941 15079
rect 9045 15045 9079 15079
rect 12173 15045 12207 15079
rect 15577 15045 15611 15079
rect 2513 14977 2547 15011
rect 2605 14977 2639 15011
rect 4537 14977 4571 15011
rect 8677 14977 8711 15011
rect 9137 14977 9171 15011
rect 13737 14977 13771 15011
rect 14565 14977 14599 15011
rect 14841 14977 14875 15011
rect 1409 14909 1443 14943
rect 2973 14909 3007 14943
rect 3709 14909 3743 14943
rect 6837 14909 6871 14943
rect 7389 14909 7423 14943
rect 10701 14909 10735 14943
rect 11161 14909 11195 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 15945 14909 15979 14943
rect 16129 14909 16163 14943
rect 4261 14841 4295 14875
rect 4353 14841 4387 14875
rect 5733 14841 5767 14875
rect 8769 14841 8803 14875
rect 10333 14841 10367 14875
rect 13185 14841 13219 14875
rect 14657 14841 14691 14875
rect 4077 14773 4111 14807
rect 6285 14773 6319 14807
rect 6929 14773 6963 14807
rect 9413 14773 9447 14807
rect 9873 14773 9907 14807
rect 11437 14773 11471 14807
rect 11805 14773 11839 14807
rect 14289 14773 14323 14807
rect 1685 14569 1719 14603
rect 2973 14569 3007 14603
rect 7113 14569 7147 14603
rect 8033 14569 8067 14603
rect 8953 14569 8987 14603
rect 9321 14569 9355 14603
rect 10517 14569 10551 14603
rect 11345 14569 11379 14603
rect 12173 14569 12207 14603
rect 12909 14569 12943 14603
rect 14657 14569 14691 14603
rect 16405 14569 16439 14603
rect 2053 14501 2087 14535
rect 5549 14501 5583 14535
rect 6555 14501 6589 14535
rect 7481 14501 7515 14535
rect 7849 14501 7883 14535
rect 13782 14501 13816 14535
rect 15577 14501 15611 14535
rect 4721 14433 4755 14467
rect 6193 14433 6227 14467
rect 8217 14433 8251 14467
rect 8493 14433 8527 14467
rect 9689 14433 9723 14467
rect 10241 14433 10275 14467
rect 11529 14433 11563 14467
rect 12449 14433 12483 14467
rect 13461 14433 13495 14467
rect 16957 14433 16991 14467
rect 1961 14365 1995 14399
rect 2421 14365 2455 14399
rect 4077 14365 4111 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 13277 14297 13311 14331
rect 17095 14297 17129 14331
rect 3249 14229 3283 14263
rect 5273 14229 5307 14263
rect 9873 14229 9907 14263
rect 12633 14229 12667 14263
rect 14381 14229 14415 14263
rect 4169 14025 4203 14059
rect 10885 14025 10919 14059
rect 11897 14025 11931 14059
rect 12265 14025 12299 14059
rect 14565 14025 14599 14059
rect 7757 13957 7791 13991
rect 8999 13957 9033 13991
rect 9137 13957 9171 13991
rect 9965 13957 9999 13991
rect 10590 13957 10624 13991
rect 10701 13957 10735 13991
rect 15761 13957 15795 13991
rect 17141 13957 17175 13991
rect 1593 13889 1627 13923
rect 2513 13889 2547 13923
rect 3433 13889 3467 13923
rect 8769 13889 8803 13923
rect 9229 13889 9263 13923
rect 10793 13889 10827 13923
rect 15025 13889 15059 13923
rect 16681 13889 16715 13923
rect 5089 13821 5123 13855
rect 5181 13821 5215 13855
rect 5641 13821 5675 13855
rect 6837 13821 6871 13855
rect 8401 13821 8435 13855
rect 8861 13821 8895 13855
rect 10425 13821 10459 13855
rect 12817 13821 12851 13855
rect 1685 13753 1719 13787
rect 2237 13753 2271 13787
rect 3157 13753 3191 13787
rect 3249 13753 3283 13787
rect 7158 13753 7192 13787
rect 12725 13753 12759 13787
rect 13179 13753 13213 13787
rect 14013 13753 14047 13787
rect 15209 13753 15243 13787
rect 15301 13753 15335 13787
rect 16497 13753 16531 13787
rect 2973 13685 3007 13719
rect 5457 13685 5491 13719
rect 6193 13685 6227 13719
rect 6561 13685 6595 13719
rect 9505 13685 9539 13719
rect 10333 13685 10367 13719
rect 11529 13685 11563 13719
rect 13737 13685 13771 13719
rect 16129 13685 16163 13719
rect 2605 13481 2639 13515
rect 6101 13481 6135 13515
rect 6285 13481 6319 13515
rect 7297 13481 7331 13515
rect 9137 13481 9171 13515
rect 10701 13481 10735 13515
rect 11161 13481 11195 13515
rect 13461 13481 13495 13515
rect 1777 13413 1811 13447
rect 4445 13413 4479 13447
rect 10425 13413 10459 13447
rect 12633 13413 12667 13447
rect 12909 13413 12943 13447
rect 13829 13413 13863 13447
rect 14381 13413 14415 13447
rect 16037 13413 16071 13447
rect 6469 13345 6503 13379
rect 6653 13345 6687 13379
rect 8125 13345 8159 13379
rect 8585 13345 8619 13379
rect 9965 13345 9999 13379
rect 11897 13345 11931 13379
rect 12357 13345 12391 13379
rect 15393 13345 15427 13379
rect 1685 13277 1719 13311
rect 1961 13277 1995 13311
rect 2973 13277 3007 13311
rect 4353 13277 4387 13311
rect 4629 13277 4663 13311
rect 8677 13277 8711 13311
rect 13737 13277 13771 13311
rect 7849 13141 7883 13175
rect 9413 13141 9447 13175
rect 2605 12937 2639 12971
rect 6285 12937 6319 12971
rect 8125 12937 8159 12971
rect 10885 12937 10919 12971
rect 11253 12937 11287 12971
rect 11989 12937 12023 12971
rect 13645 12937 13679 12971
rect 15393 12937 15427 12971
rect 4537 12869 4571 12903
rect 5917 12869 5951 12903
rect 12633 12869 12667 12903
rect 1593 12801 1627 12835
rect 1961 12801 1995 12835
rect 2973 12801 3007 12835
rect 4169 12801 4203 12835
rect 4997 12801 5031 12835
rect 6653 12801 6687 12835
rect 8677 12801 8711 12835
rect 10977 12801 11011 12835
rect 11621 12801 11655 12835
rect 13737 12801 13771 12835
rect 7113 12733 7147 12767
rect 7665 12733 7699 12767
rect 9597 12733 9631 12767
rect 10756 12733 10790 12767
rect 12449 12733 12483 12767
rect 12909 12733 12943 12767
rect 13829 12733 13863 12767
rect 1685 12665 1719 12699
rect 3525 12665 3559 12699
rect 3617 12665 3651 12699
rect 7849 12665 7883 12699
rect 8998 12665 9032 12699
rect 10609 12665 10643 12699
rect 3249 12597 3283 12631
rect 4905 12597 4939 12631
rect 5365 12597 5399 12631
rect 8493 12597 8527 12631
rect 9965 12597 9999 12631
rect 10517 12597 10551 12631
rect 1409 12393 1443 12427
rect 2237 12393 2271 12427
rect 3525 12393 3559 12427
rect 4077 12393 4111 12427
rect 4537 12393 4571 12427
rect 5089 12393 5123 12427
rect 6653 12393 6687 12427
rect 7757 12393 7791 12427
rect 9045 12393 9079 12427
rect 11069 12393 11103 12427
rect 11897 12393 11931 12427
rect 12357 12393 12391 12427
rect 13093 12393 13127 12427
rect 13829 12393 13863 12427
rect 3157 12325 3191 12359
rect 5819 12325 5853 12359
rect 8170 12325 8204 12359
rect 9873 12325 9907 12359
rect 11253 12325 11287 12359
rect 12817 12325 12851 12359
rect 3065 12257 3099 12291
rect 5457 12257 5491 12291
rect 7849 12257 7883 12291
rect 13001 12257 13035 12291
rect 9781 12189 9815 12223
rect 10057 12189 10091 12223
rect 11621 12189 11655 12223
rect 9413 12121 9447 12155
rect 14105 12121 14139 12155
rect 1961 12053 1995 12087
rect 6377 12053 6411 12087
rect 7113 12053 7147 12087
rect 8769 12053 8803 12087
rect 10701 12053 10735 12087
rect 11391 12053 11425 12087
rect 11529 12053 11563 12087
rect 1961 11849 1995 11883
rect 2605 11849 2639 11883
rect 6193 11849 6227 11883
rect 7941 11849 7975 11883
rect 10793 11849 10827 11883
rect 11437 11849 11471 11883
rect 9137 11781 9171 11815
rect 12817 11781 12851 11815
rect 3617 11713 3651 11747
rect 4261 11713 4295 11747
rect 5457 11713 5491 11747
rect 7113 11713 7147 11747
rect 8493 11713 8527 11747
rect 9781 11713 9815 11747
rect 10057 11713 10091 11747
rect 2145 11645 2179 11679
rect 11253 11645 11287 11679
rect 11713 11645 11747 11679
rect 12081 11645 12115 11679
rect 3433 11577 3467 11611
rect 3702 11577 3736 11611
rect 5181 11577 5215 11611
rect 5273 11577 5307 11611
rect 8217 11577 8251 11611
rect 8309 11577 8343 11611
rect 9873 11577 9907 11611
rect 4629 11509 4663 11543
rect 4997 11509 5031 11543
rect 9597 11509 9631 11543
rect 11069 11509 11103 11543
rect 13277 11509 13311 11543
rect 1685 11305 1719 11339
rect 2697 11305 2731 11339
rect 5457 11305 5491 11339
rect 6929 11305 6963 11339
rect 7665 11305 7699 11339
rect 8769 11305 8803 11339
rect 9505 11305 9539 11339
rect 11345 11305 11379 11339
rect 4353 11237 4387 11271
rect 7941 11237 7975 11271
rect 8493 11237 8527 11271
rect 9689 11237 9723 11271
rect 2881 11169 2915 11203
rect 4997 11169 5031 11203
rect 6745 11169 6779 11203
rect 9781 11169 9815 11203
rect 7849 11101 7883 11135
rect 7297 11033 7331 11067
rect 3525 10965 3559 10999
rect 1593 10761 1627 10795
rect 2651 10761 2685 10795
rect 4077 10761 4111 10795
rect 4445 10761 4479 10795
rect 5687 10761 5721 10795
rect 8861 10761 8895 10795
rect 9597 10761 9631 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 3663 10693 3697 10727
rect 4675 10693 4709 10727
rect 2329 10625 2363 10659
rect 7021 10625 7055 10659
rect 7757 10625 7791 10659
rect 7849 10625 7883 10659
rect 1409 10557 1443 10591
rect 2548 10557 2582 10591
rect 2973 10557 3007 10591
rect 3592 10557 3626 10591
rect 4261 10557 4295 10591
rect 4572 10557 4606 10591
rect 4997 10557 5031 10591
rect 5584 10557 5618 10591
rect 6009 10557 6043 10591
rect 8493 10557 8527 10591
rect 9413 10557 9447 10591
rect 9873 10557 9907 10591
rect 10425 10557 10459 10591
rect 4169 10421 4203 10455
rect 10977 10421 11011 10455
rect 2559 10217 2593 10251
rect 4215 10217 4249 10251
rect 8585 10217 8619 10251
rect 1547 10149 1581 10183
rect 1460 10081 1494 10115
rect 2488 10081 2522 10115
rect 4112 10081 4146 10115
rect 7573 10081 7607 10115
rect 8125 10081 8159 10115
rect 7941 10013 7975 10047
rect 1961 9877 1995 9911
rect 1547 9673 1581 9707
rect 2329 9673 2363 9707
rect 2559 9673 2593 9707
rect 3617 9673 3651 9707
rect 4169 9673 4203 9707
rect 3157 9605 3191 9639
rect 3249 9605 3283 9639
rect 4583 9605 4617 9639
rect 1476 9469 1510 9503
rect 1869 9469 1903 9503
rect 2488 9469 2522 9503
rect 2881 9469 2915 9503
rect 3157 9469 3191 9503
rect 3468 9469 3502 9503
rect 4512 9469 4546 9503
rect 4905 9469 4939 9503
rect 7389 9469 7423 9503
rect 7113 9333 7147 9367
rect 7757 9333 7791 9367
rect 8309 9333 8343 9367
rect 1547 9129 1581 9163
rect 2559 9129 2593 9163
rect 7849 9061 7883 9095
rect 8401 9061 8435 9095
rect 1444 8993 1478 9027
rect 1961 8993 1995 9027
rect 2488 8993 2522 9027
rect 8033 8993 8067 9027
rect 7297 8857 7331 8891
rect 1869 8585 1903 8619
rect 2237 8585 2271 8619
rect 2697 8585 2731 8619
rect 3249 8585 3283 8619
rect 8217 8585 8251 8619
rect 1685 8517 1719 8551
rect 2881 8517 2915 8551
rect 1476 8381 1510 8415
rect 2456 8381 2490 8415
rect 7941 8245 7975 8279
rect 1409 7905 1443 7939
rect 1547 7769 1581 7803
rect 1593 7497 1627 7531
rect 1409 6817 1443 6851
rect 1547 6749 1581 6783
rect 1593 6409 1627 6443
rect 1444 5729 1478 5763
rect 1547 5661 1581 5695
rect 1593 5321 1627 5355
rect 1444 4641 1478 4675
rect 1547 4573 1581 4607
rect 1593 4233 1627 4267
rect 1593 3689 1627 3723
rect 1444 3553 1478 3587
rect 2237 3145 2271 3179
rect 1444 2941 1478 2975
rect 1869 2941 1903 2975
rect 1547 2805 1581 2839
rect 2559 2601 2593 2635
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 2456 2465 2490 2499
rect 2881 2465 2915 2499
rect 1547 2397 1581 2431
<< metal1 >>
rect 2498 26188 2504 26240
rect 2556 26228 2562 26240
rect 18230 26228 18236 26240
rect 2556 26200 18236 26228
rect 2556 26188 2562 26200
rect 18230 26188 18236 26200
rect 18288 26188 18294 26240
rect 1486 26120 1492 26172
rect 1544 26160 1550 26172
rect 16574 26160 16580 26172
rect 1544 26132 16580 26160
rect 1544 26120 1550 26132
rect 16574 26120 16580 26132
rect 16632 26120 16638 26172
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 106 25440 112 25492
rect 164 25480 170 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 164 25452 4261 25480
rect 164 25440 170 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 4249 25443 4307 25449
rect 4525 25483 4583 25489
rect 4525 25449 4537 25483
rect 4571 25480 4583 25483
rect 4709 25483 4767 25489
rect 4709 25480 4721 25483
rect 4571 25452 4721 25480
rect 4571 25449 4583 25452
rect 4525 25443 4583 25449
rect 4709 25449 4721 25452
rect 4755 25480 4767 25483
rect 12345 25483 12403 25489
rect 12345 25480 12357 25483
rect 4755 25452 12357 25480
rect 4755 25449 4767 25452
rect 4709 25443 4767 25449
rect 12345 25449 12357 25452
rect 12391 25449 12403 25483
rect 12345 25443 12403 25449
rect 15473 25483 15531 25489
rect 15473 25449 15485 25483
rect 15519 25480 15531 25483
rect 15654 25480 15660 25492
rect 15519 25452 15660 25480
rect 15519 25449 15531 25452
rect 15473 25443 15531 25449
rect 15654 25440 15660 25452
rect 15712 25480 15718 25492
rect 17034 25480 17040 25492
rect 15712 25452 17040 25480
rect 15712 25440 15718 25452
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 2866 25372 2872 25424
rect 2924 25412 2930 25424
rect 18463 25415 18521 25421
rect 18463 25412 18475 25415
rect 2924 25384 18475 25412
rect 2924 25372 2930 25384
rect 18463 25381 18475 25384
rect 18509 25381 18521 25415
rect 18463 25375 18521 25381
rect 2498 25344 2504 25356
rect 2459 25316 2504 25344
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4525 25347 4583 25353
rect 4525 25344 4537 25347
rect 4111 25316 4537 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4525 25313 4537 25316
rect 4571 25313 4583 25347
rect 4525 25307 4583 25313
rect 5813 25347 5871 25353
rect 5813 25313 5825 25347
rect 5859 25344 5871 25347
rect 6086 25344 6092 25356
rect 5859 25316 6092 25344
rect 5859 25313 5871 25316
rect 5813 25307 5871 25313
rect 6086 25304 6092 25316
rect 6144 25304 6150 25356
rect 8294 25344 8300 25356
rect 8255 25316 8300 25344
rect 8294 25304 8300 25316
rect 8352 25304 8358 25356
rect 9858 25344 9864 25356
rect 9819 25316 9864 25344
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 11400 25347 11458 25353
rect 11400 25313 11412 25347
rect 11446 25344 11458 25347
rect 11790 25344 11796 25356
rect 11446 25316 11796 25344
rect 11446 25313 11458 25316
rect 11400 25307 11458 25313
rect 11790 25304 11796 25316
rect 11848 25304 11854 25356
rect 12894 25344 12900 25356
rect 12855 25316 12900 25344
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 13906 25344 13912 25356
rect 13867 25316 13912 25344
rect 13906 25304 13912 25316
rect 13964 25304 13970 25356
rect 16574 25344 16580 25356
rect 16535 25316 16580 25344
rect 16574 25304 16580 25316
rect 16632 25304 16638 25356
rect 18230 25344 18236 25356
rect 18191 25316 18236 25344
rect 18230 25304 18236 25316
rect 18288 25304 18294 25356
rect 19334 25344 19340 25356
rect 19295 25316 19340 25344
rect 19334 25304 19340 25316
rect 19392 25304 19398 25356
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 2406 25276 2412 25288
rect 2367 25248 2412 25276
rect 2406 25236 2412 25248
rect 2464 25236 2470 25288
rect 5166 25276 5172 25288
rect 5127 25248 5172 25276
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 7742 25276 7748 25288
rect 7703 25248 7748 25276
rect 7742 25236 7748 25248
rect 7800 25236 7806 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 15470 25276 15476 25288
rect 12391 25248 15476 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 15470 25236 15476 25248
rect 15528 25236 15534 25288
rect 16715 25211 16773 25217
rect 16715 25208 16727 25211
rect 4126 25180 16727 25208
rect 3050 25100 3056 25152
rect 3108 25140 3114 25152
rect 4126 25140 4154 25180
rect 16715 25177 16727 25180
rect 16761 25177 16773 25211
rect 16715 25171 16773 25177
rect 10042 25140 10048 25152
rect 3108 25112 4154 25140
rect 10003 25112 10048 25140
rect 3108 25100 3114 25112
rect 10042 25100 10048 25112
rect 10100 25100 10106 25152
rect 11471 25143 11529 25149
rect 11471 25109 11483 25143
rect 11517 25140 11529 25143
rect 11882 25140 11888 25152
rect 11517 25112 11888 25140
rect 11517 25109 11529 25112
rect 11471 25103 11529 25109
rect 11882 25100 11888 25112
rect 11940 25100 11946 25152
rect 13035 25143 13093 25149
rect 13035 25109 13047 25143
rect 13081 25140 13093 25143
rect 13722 25140 13728 25152
rect 13081 25112 13728 25140
rect 13081 25109 13093 25112
rect 13035 25103 13093 25109
rect 13722 25100 13728 25112
rect 13780 25100 13786 25152
rect 13814 25100 13820 25152
rect 13872 25140 13878 25152
rect 14047 25143 14105 25149
rect 14047 25140 14059 25143
rect 13872 25112 14059 25140
rect 13872 25100 13878 25112
rect 14047 25109 14059 25112
rect 14093 25109 14105 25143
rect 14047 25103 14105 25109
rect 15703 25143 15761 25149
rect 15703 25109 15715 25143
rect 15749 25140 15761 25143
rect 15838 25140 15844 25152
rect 15749 25112 15844 25140
rect 15749 25109 15761 25112
rect 15703 25103 15761 25109
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 18598 25100 18604 25152
rect 18656 25140 18662 25152
rect 19475 25143 19533 25149
rect 19475 25140 19487 25143
rect 18656 25112 19487 25140
rect 18656 25100 18662 25112
rect 19475 25109 19487 25112
rect 19521 25109 19533 25143
rect 19475 25103 19533 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 5077 24939 5135 24945
rect 5077 24905 5089 24939
rect 5123 24936 5135 24939
rect 5166 24936 5172 24948
rect 5123 24908 5172 24936
rect 5123 24905 5135 24908
rect 5077 24899 5135 24905
rect 5166 24896 5172 24908
rect 5224 24896 5230 24948
rect 9858 24936 9864 24948
rect 9819 24908 9864 24936
rect 9858 24896 9864 24908
rect 9916 24896 9922 24948
rect 11790 24936 11796 24948
rect 11751 24908 11796 24936
rect 11790 24896 11796 24908
rect 11848 24896 11854 24948
rect 12894 24896 12900 24948
rect 12952 24936 12958 24948
rect 13449 24939 13507 24945
rect 13449 24936 13461 24939
rect 12952 24908 13461 24936
rect 12952 24896 12958 24908
rect 13449 24905 13461 24908
rect 13495 24905 13507 24939
rect 13449 24899 13507 24905
rect 13906 24896 13912 24948
rect 13964 24936 13970 24948
rect 14461 24939 14519 24945
rect 14461 24936 14473 24939
rect 13964 24908 14473 24936
rect 13964 24896 13970 24908
rect 14461 24905 14473 24908
rect 14507 24905 14519 24939
rect 14826 24936 14832 24948
rect 14787 24908 14832 24936
rect 14461 24899 14519 24905
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 15654 24936 15660 24948
rect 15615 24908 15660 24936
rect 15654 24896 15660 24908
rect 15712 24896 15718 24948
rect 16574 24936 16580 24948
rect 16535 24908 16580 24936
rect 16574 24896 16580 24908
rect 16632 24896 16638 24948
rect 18230 24896 18236 24948
rect 18288 24936 18294 24948
rect 18509 24939 18567 24945
rect 18509 24936 18521 24939
rect 18288 24908 18521 24936
rect 18288 24896 18294 24908
rect 18509 24905 18521 24908
rect 18555 24905 18567 24939
rect 18509 24899 18567 24905
rect 5350 24828 5356 24880
rect 5408 24868 5414 24880
rect 18598 24868 18604 24880
rect 5408 24840 18604 24868
rect 5408 24828 5414 24840
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 1394 24760 1400 24812
rect 1452 24800 1458 24812
rect 1946 24800 1952 24812
rect 1452 24772 1952 24800
rect 1452 24760 1458 24772
rect 1946 24760 1952 24772
rect 2004 24760 2010 24812
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24800 4767 24803
rect 6086 24800 6092 24812
rect 4755 24772 6092 24800
rect 4755 24769 4767 24772
rect 4709 24763 4767 24769
rect 6086 24760 6092 24772
rect 6144 24760 6150 24812
rect 9766 24760 9772 24812
rect 9824 24800 9830 24812
rect 9824 24772 14964 24800
rect 9824 24760 9830 24772
rect 3513 24735 3571 24741
rect 3513 24701 3525 24735
rect 3559 24732 3571 24735
rect 4246 24732 4252 24744
rect 3559 24704 4252 24732
rect 3559 24701 3571 24704
rect 3513 24695 3571 24701
rect 4246 24692 4252 24704
rect 4304 24692 4310 24744
rect 6546 24692 6552 24744
rect 6604 24732 6610 24744
rect 6641 24735 6699 24741
rect 6641 24732 6653 24735
rect 6604 24704 6653 24732
rect 6604 24692 6610 24704
rect 6641 24701 6653 24704
rect 6687 24732 6699 24735
rect 6917 24735 6975 24741
rect 6917 24732 6929 24735
rect 6687 24704 6929 24732
rect 6687 24701 6699 24704
rect 6641 24695 6699 24701
rect 6917 24701 6929 24704
rect 6963 24701 6975 24735
rect 8478 24732 8484 24744
rect 8391 24704 8484 24732
rect 6917 24695 6975 24701
rect 8478 24692 8484 24704
rect 8536 24732 8542 24744
rect 8665 24735 8723 24741
rect 8665 24732 8677 24735
rect 8536 24704 8677 24732
rect 8536 24692 8542 24704
rect 8665 24701 8677 24704
rect 8711 24701 8723 24735
rect 8665 24695 8723 24701
rect 10689 24735 10747 24741
rect 10689 24701 10701 24735
rect 10735 24732 10747 24735
rect 10870 24732 10876 24744
rect 10735 24704 10876 24732
rect 10735 24701 10747 24704
rect 10689 24695 10747 24701
rect 10870 24692 10876 24704
rect 10928 24692 10934 24744
rect 12250 24732 12256 24744
rect 12163 24704 12256 24732
rect 12250 24692 12256 24704
rect 12308 24732 12314 24744
rect 12529 24735 12587 24741
rect 12529 24732 12541 24735
rect 12308 24704 12541 24732
rect 12308 24692 12314 24704
rect 12529 24701 12541 24704
rect 12575 24701 12587 24735
rect 12529 24695 12587 24701
rect 14052 24735 14110 24741
rect 14052 24701 14064 24735
rect 14098 24732 14110 24735
rect 14826 24732 14832 24744
rect 14098 24704 14832 24732
rect 14098 24701 14110 24704
rect 14052 24695 14110 24701
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 1765 24667 1823 24673
rect 1765 24633 1777 24667
rect 1811 24664 1823 24667
rect 2041 24667 2099 24673
rect 2041 24664 2053 24667
rect 1811 24636 2053 24664
rect 1811 24633 1823 24636
rect 1765 24627 1823 24633
rect 2041 24633 2053 24636
rect 2087 24664 2099 24667
rect 2222 24664 2228 24676
rect 2087 24636 2228 24664
rect 2087 24633 2099 24636
rect 2041 24627 2099 24633
rect 2222 24624 2228 24636
rect 2280 24624 2286 24676
rect 2590 24664 2596 24676
rect 2551 24636 2596 24664
rect 2590 24624 2596 24636
rect 2648 24624 2654 24676
rect 5258 24664 5264 24676
rect 5219 24636 5264 24664
rect 5258 24624 5264 24636
rect 5316 24624 5322 24676
rect 5353 24667 5411 24673
rect 5353 24633 5365 24667
rect 5399 24633 5411 24667
rect 5353 24627 5411 24633
rect 5905 24667 5963 24673
rect 5905 24633 5917 24667
rect 5951 24664 5963 24667
rect 6454 24664 6460 24676
rect 5951 24636 6460 24664
rect 5951 24633 5963 24636
rect 5905 24627 5963 24633
rect 2498 24556 2504 24608
rect 2556 24596 2562 24608
rect 2869 24599 2927 24605
rect 2869 24596 2881 24599
rect 2556 24568 2881 24596
rect 2556 24556 2562 24568
rect 2869 24565 2881 24568
rect 2915 24565 2927 24599
rect 3878 24596 3884 24608
rect 3839 24568 3884 24596
rect 2869 24559 2927 24565
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5368 24596 5396 24627
rect 6454 24624 6460 24636
rect 6512 24624 6518 24676
rect 6822 24664 6828 24676
rect 6783 24636 6828 24664
rect 6822 24624 6828 24636
rect 6880 24624 6886 24676
rect 10778 24664 10784 24676
rect 10739 24636 10784 24664
rect 10778 24624 10784 24636
rect 10836 24624 10842 24676
rect 12434 24664 12440 24676
rect 12395 24636 12440 24664
rect 12434 24624 12440 24636
rect 12492 24624 12498 24676
rect 14139 24667 14197 24673
rect 14139 24633 14151 24667
rect 14185 24664 14197 24667
rect 14550 24664 14556 24676
rect 14185 24636 14556 24664
rect 14185 24633 14197 24636
rect 14139 24627 14197 24633
rect 14550 24624 14556 24636
rect 14608 24624 14614 24676
rect 14936 24664 14964 24772
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 19199 24803 19257 24809
rect 19199 24800 19211 24803
rect 15528 24772 19211 24800
rect 15528 24760 15534 24772
rect 19199 24769 19211 24772
rect 19245 24769 19257 24803
rect 19199 24763 19257 24769
rect 15841 24735 15899 24741
rect 15841 24701 15853 24735
rect 15887 24732 15899 24735
rect 15930 24732 15936 24744
rect 15887 24704 15936 24732
rect 15887 24701 15899 24704
rect 15841 24695 15899 24701
rect 15930 24692 15936 24704
rect 15988 24692 15994 24744
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 18084 24735 18142 24741
rect 18084 24732 18096 24735
rect 18012 24704 18096 24732
rect 18012 24692 18018 24704
rect 18084 24701 18096 24704
rect 18130 24732 18142 24735
rect 18877 24735 18935 24741
rect 18877 24732 18889 24735
rect 18130 24704 18889 24732
rect 18130 24701 18142 24704
rect 18084 24695 18142 24701
rect 18877 24701 18889 24704
rect 18923 24701 18935 24735
rect 18877 24695 18935 24701
rect 18966 24692 18972 24744
rect 19024 24732 19030 24744
rect 19096 24735 19154 24741
rect 19096 24732 19108 24735
rect 19024 24704 19108 24732
rect 19024 24692 19030 24704
rect 19096 24701 19108 24704
rect 19142 24732 19154 24735
rect 19889 24735 19947 24741
rect 19889 24732 19901 24735
rect 19142 24704 19901 24732
rect 19142 24701 19154 24704
rect 19096 24695 19154 24701
rect 19889 24701 19901 24704
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 17126 24664 17132 24676
rect 14936 24636 17132 24664
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 18690 24624 18696 24676
rect 18748 24664 18754 24676
rect 19334 24664 19340 24676
rect 18748 24636 19340 24664
rect 18748 24624 18754 24636
rect 19334 24624 19340 24636
rect 19392 24664 19398 24676
rect 19521 24667 19579 24673
rect 19521 24664 19533 24667
rect 19392 24636 19533 24664
rect 19392 24624 19398 24636
rect 19521 24633 19533 24636
rect 19567 24633 19579 24667
rect 19521 24627 19579 24633
rect 5224 24568 5396 24596
rect 7929 24599 7987 24605
rect 5224 24556 5230 24568
rect 7929 24565 7941 24599
rect 7975 24596 7987 24599
rect 8294 24596 8300 24608
rect 7975 24568 8300 24596
rect 7975 24565 7987 24568
rect 7929 24559 7987 24565
rect 8294 24556 8300 24568
rect 8352 24556 8358 24608
rect 8846 24596 8852 24608
rect 8807 24568 8852 24596
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 16071 24599 16129 24605
rect 16071 24565 16083 24599
rect 16117 24596 16129 24599
rect 16482 24596 16488 24608
rect 16117 24568 16488 24596
rect 16117 24565 16129 24568
rect 16071 24559 16129 24565
rect 16482 24556 16488 24568
rect 16540 24556 16546 24608
rect 16942 24596 16948 24608
rect 16903 24568 16948 24596
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 18187 24599 18245 24605
rect 18187 24596 18199 24599
rect 17092 24568 18199 24596
rect 17092 24556 17098 24568
rect 18187 24565 18199 24568
rect 18233 24565 18245 24599
rect 18187 24559 18245 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1946 24392 1952 24404
rect 1907 24364 1952 24392
rect 1946 24352 1952 24364
rect 2004 24352 2010 24404
rect 4338 24352 4344 24404
rect 4396 24392 4402 24404
rect 6822 24392 6828 24404
rect 4396 24364 6828 24392
rect 4396 24352 4402 24364
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 11882 24392 11888 24404
rect 11843 24364 11888 24392
rect 11882 24352 11888 24364
rect 11940 24392 11946 24404
rect 18509 24395 18567 24401
rect 11940 24364 12204 24392
rect 11940 24352 11946 24364
rect 2314 24324 2320 24336
rect 2275 24296 2320 24324
rect 2314 24284 2320 24296
rect 2372 24284 2378 24336
rect 4246 24324 4252 24336
rect 4159 24296 4252 24324
rect 4246 24284 4252 24296
rect 4304 24324 4310 24336
rect 4982 24324 4988 24336
rect 4304 24296 4988 24324
rect 4304 24284 4310 24296
rect 4982 24284 4988 24296
rect 5040 24284 5046 24336
rect 5813 24327 5871 24333
rect 5813 24293 5825 24327
rect 5859 24324 5871 24327
rect 6086 24324 6092 24336
rect 5859 24296 6092 24324
rect 5859 24293 5871 24296
rect 5813 24287 5871 24293
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 6365 24327 6423 24333
rect 6365 24293 6377 24327
rect 6411 24324 6423 24327
rect 6454 24324 6460 24336
rect 6411 24296 6460 24324
rect 6411 24293 6423 24296
rect 6365 24287 6423 24293
rect 6454 24284 6460 24296
rect 6512 24284 6518 24336
rect 8205 24327 8263 24333
rect 8205 24293 8217 24327
rect 8251 24324 8263 24327
rect 8294 24324 8300 24336
rect 8251 24296 8300 24324
rect 8251 24293 8263 24296
rect 8205 24287 8263 24293
rect 8294 24284 8300 24296
rect 8352 24284 8358 24336
rect 9858 24284 9864 24336
rect 9916 24324 9922 24336
rect 12176 24333 12204 24364
rect 18509 24361 18521 24395
rect 18555 24392 18567 24395
rect 21174 24392 21180 24404
rect 18555 24364 21180 24392
rect 18555 24361 18567 24364
rect 18509 24355 18567 24361
rect 21174 24352 21180 24364
rect 21232 24352 21238 24404
rect 10137 24327 10195 24333
rect 10137 24324 10149 24327
rect 9916 24296 10149 24324
rect 9916 24284 9922 24296
rect 10137 24293 10149 24296
rect 10183 24293 10195 24327
rect 10137 24287 10195 24293
rect 12161 24327 12219 24333
rect 12161 24293 12173 24327
rect 12207 24293 12219 24327
rect 12161 24287 12219 24293
rect 12250 24284 12256 24336
rect 12308 24324 12314 24336
rect 15746 24324 15752 24336
rect 12308 24296 12353 24324
rect 15463 24296 15752 24324
rect 12308 24284 12314 24296
rect 14090 24256 14096 24268
rect 14051 24228 14096 24256
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 15463 24265 15491 24296
rect 15746 24284 15752 24296
rect 15804 24324 15810 24336
rect 18046 24324 18052 24336
rect 15804 24296 18052 24324
rect 15804 24284 15810 24296
rect 18046 24284 18052 24296
rect 18104 24284 18110 24336
rect 15448 24259 15506 24265
rect 15448 24225 15460 24259
rect 15494 24225 15506 24259
rect 15448 24219 15506 24225
rect 16715 24259 16773 24265
rect 16715 24225 16727 24259
rect 16761 24256 16773 24259
rect 18325 24259 18383 24265
rect 18325 24256 18337 24259
rect 16761 24228 18337 24256
rect 16761 24225 16773 24228
rect 16715 24219 16773 24225
rect 18325 24225 18337 24228
rect 18371 24256 18383 24259
rect 19058 24256 19064 24268
rect 18371 24228 19064 24256
rect 18371 24225 18383 24228
rect 18325 24219 18383 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 19493 24256 19499 24268
rect 19454 24228 19499 24256
rect 19493 24216 19499 24228
rect 19551 24216 19557 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24157 2283 24191
rect 2590 24188 2596 24200
rect 2551 24160 2596 24188
rect 2225 24151 2283 24157
rect 2130 24080 2136 24132
rect 2188 24120 2194 24132
rect 2240 24120 2268 24151
rect 2590 24148 2596 24160
rect 2648 24148 2654 24200
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4212 24160 4257 24188
rect 4212 24148 4218 24160
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4672 24160 4813 24188
rect 4672 24148 4678 24160
rect 4801 24157 4813 24160
rect 4847 24188 4859 24191
rect 5721 24191 5779 24197
rect 5721 24188 5733 24191
rect 4847 24160 5733 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 5721 24157 5733 24160
rect 5767 24188 5779 24191
rect 6362 24188 6368 24200
rect 5767 24160 6368 24188
rect 5767 24157 5779 24160
rect 5721 24151 5779 24157
rect 6362 24148 6368 24160
rect 6420 24148 6426 24200
rect 8113 24191 8171 24197
rect 8113 24157 8125 24191
rect 8159 24157 8171 24191
rect 8386 24188 8392 24200
rect 8347 24160 8392 24188
rect 8113 24151 8171 24157
rect 3145 24123 3203 24129
rect 3145 24120 3157 24123
rect 2188 24092 3157 24120
rect 2188 24080 2194 24092
rect 3145 24089 3157 24092
rect 3191 24089 3203 24123
rect 3145 24083 3203 24089
rect 7929 24123 7987 24129
rect 7929 24089 7941 24123
rect 7975 24120 7987 24123
rect 8128 24120 8156 24151
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 10045 24191 10103 24197
rect 10045 24188 10057 24191
rect 9824 24160 10057 24188
rect 9824 24148 9830 24160
rect 10045 24157 10057 24160
rect 10091 24157 10103 24191
rect 10686 24188 10692 24200
rect 10647 24160 10692 24188
rect 10045 24151 10103 24157
rect 10686 24148 10692 24160
rect 10744 24148 10750 24200
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 13081 24191 13139 24197
rect 13081 24188 13093 24191
rect 12851 24160 13093 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 13081 24157 13093 24160
rect 13127 24188 13139 24191
rect 13170 24188 13176 24200
rect 13127 24160 13176 24188
rect 13127 24157 13139 24160
rect 13081 24151 13139 24157
rect 13170 24148 13176 24160
rect 13228 24148 13234 24200
rect 14366 24188 14372 24200
rect 14327 24160 14372 24188
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 8570 24120 8576 24132
rect 7975 24092 8576 24120
rect 7975 24089 7987 24092
rect 7929 24083 7987 24089
rect 8570 24080 8576 24092
rect 8628 24080 8634 24132
rect 17862 24080 17868 24132
rect 17920 24120 17926 24132
rect 19567 24123 19625 24129
rect 19567 24120 19579 24123
rect 17920 24092 19579 24120
rect 17920 24080 17926 24092
rect 19567 24089 19579 24092
rect 19613 24089 19625 24123
rect 19567 24083 19625 24089
rect 5258 24052 5264 24064
rect 5171 24024 5264 24052
rect 5258 24012 5264 24024
rect 5316 24052 5322 24064
rect 6822 24052 6828 24064
rect 5316 24024 6828 24052
rect 5316 24012 5322 24024
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 14642 24012 14648 24064
rect 14700 24052 14706 24064
rect 15519 24055 15577 24061
rect 15519 24052 15531 24055
rect 14700 24024 15531 24052
rect 14700 24012 14706 24024
rect 15519 24021 15531 24024
rect 15565 24021 15577 24055
rect 15930 24052 15936 24064
rect 15891 24024 15936 24052
rect 15519 24015 15577 24021
rect 15930 24012 15936 24024
rect 15988 24012 15994 24064
rect 16390 24012 16396 24064
rect 16448 24052 16454 24064
rect 16485 24055 16543 24061
rect 16485 24052 16497 24055
rect 16448 24024 16497 24052
rect 16448 24012 16454 24024
rect 16485 24021 16497 24024
rect 16531 24021 16543 24055
rect 19242 24052 19248 24064
rect 19203 24024 19248 24052
rect 16485 24015 16543 24021
rect 19242 24012 19248 24024
rect 19300 24012 19306 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2314 23808 2320 23860
rect 2372 23848 2378 23860
rect 2590 23848 2596 23860
rect 2372 23820 2596 23848
rect 2372 23808 2378 23820
rect 2590 23808 2596 23820
rect 2648 23808 2654 23860
rect 3789 23851 3847 23857
rect 3789 23817 3801 23851
rect 3835 23848 3847 23851
rect 3878 23848 3884 23860
rect 3835 23820 3884 23848
rect 3835 23817 3847 23820
rect 3789 23811 3847 23817
rect 3878 23808 3884 23820
rect 3936 23808 3942 23860
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 5629 23851 5687 23857
rect 5629 23848 5641 23851
rect 5592 23820 5641 23848
rect 5592 23808 5598 23820
rect 5629 23817 5641 23820
rect 5675 23817 5687 23851
rect 6362 23848 6368 23860
rect 6323 23820 6368 23848
rect 5629 23811 5687 23817
rect 6362 23808 6368 23820
rect 6420 23808 6426 23860
rect 8757 23851 8815 23857
rect 8757 23817 8769 23851
rect 8803 23848 8815 23851
rect 8846 23848 8852 23860
rect 8803 23820 8852 23848
rect 8803 23817 8815 23820
rect 8757 23811 8815 23817
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9858 23848 9864 23860
rect 9819 23820 9864 23848
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 10689 23851 10747 23857
rect 10689 23817 10701 23851
rect 10735 23848 10747 23851
rect 10778 23848 10784 23860
rect 10735 23820 10784 23848
rect 10735 23817 10747 23820
rect 10689 23811 10747 23817
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 12161 23851 12219 23857
rect 12161 23817 12173 23851
rect 12207 23848 12219 23851
rect 12250 23848 12256 23860
rect 12207 23820 12256 23848
rect 12207 23817 12219 23820
rect 12161 23811 12219 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 14090 23848 14096 23860
rect 14051 23820 14096 23848
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 14366 23808 14372 23860
rect 14424 23848 14430 23860
rect 14461 23851 14519 23857
rect 14461 23848 14473 23851
rect 14424 23820 14473 23848
rect 14424 23808 14430 23820
rect 14461 23817 14473 23820
rect 14507 23817 14519 23851
rect 15746 23848 15752 23860
rect 15707 23820 15752 23848
rect 14461 23811 14519 23817
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 18782 23848 18788 23860
rect 17083 23820 18788 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 19058 23848 19064 23860
rect 19019 23820 19064 23848
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 19429 23851 19487 23857
rect 19429 23817 19441 23851
rect 19475 23848 19487 23851
rect 22186 23848 22192 23860
rect 19475 23820 22192 23848
rect 19475 23817 19487 23820
rect 19429 23811 19487 23817
rect 22186 23808 22192 23820
rect 22244 23808 22250 23860
rect 24949 23851 25007 23857
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 27338 23848 27344 23860
rect 24995 23820 27344 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 27338 23808 27344 23820
rect 27396 23808 27402 23860
rect 18325 23783 18383 23789
rect 14384 23752 15056 23780
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 1854 23712 1860 23724
rect 1719 23684 1860 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 2130 23712 2136 23724
rect 2091 23684 2136 23712
rect 2130 23672 2136 23684
rect 2188 23712 2194 23724
rect 2314 23712 2320 23724
rect 2188 23684 2320 23712
rect 2188 23672 2194 23684
rect 2314 23672 2320 23684
rect 2372 23672 2378 23724
rect 3421 23715 3479 23721
rect 3421 23681 3433 23715
rect 3467 23712 3479 23715
rect 4154 23712 4160 23724
rect 3467 23684 4160 23712
rect 3467 23681 3479 23684
rect 3421 23675 3479 23681
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 4614 23712 4620 23724
rect 4575 23684 4620 23712
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23712 8079 23715
rect 8110 23712 8116 23724
rect 8067 23684 8116 23712
rect 8067 23681 8079 23684
rect 8021 23675 8079 23681
rect 8110 23672 8116 23684
rect 8168 23712 8174 23724
rect 8386 23712 8392 23724
rect 8168 23684 8392 23712
rect 8168 23672 8174 23684
rect 8386 23672 8392 23684
rect 8444 23672 8450 23724
rect 9214 23712 9220 23724
rect 9175 23684 9220 23712
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 11330 23712 11336 23724
rect 10704 23684 11336 23712
rect 5433 23647 5491 23653
rect 5433 23644 5445 23647
rect 5368 23616 5445 23644
rect 1762 23536 1768 23588
rect 1820 23576 1826 23588
rect 2958 23576 2964 23588
rect 1820 23548 1865 23576
rect 2919 23548 2964 23576
rect 1820 23536 1826 23548
rect 2958 23536 2964 23548
rect 3016 23576 3022 23588
rect 3973 23579 4031 23585
rect 3973 23576 3985 23579
rect 3016 23548 3985 23576
rect 3016 23536 3022 23548
rect 3973 23545 3985 23548
rect 4019 23545 4031 23579
rect 3973 23539 4031 23545
rect 4065 23579 4123 23585
rect 4065 23545 4077 23579
rect 4111 23545 4123 23579
rect 4065 23539 4123 23545
rect 3878 23468 3884 23520
rect 3936 23508 3942 23520
rect 4080 23508 4108 23539
rect 4982 23508 4988 23520
rect 3936 23480 4108 23508
rect 4943 23480 4988 23508
rect 3936 23468 3942 23480
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 5368 23517 5396 23616
rect 5433 23613 5445 23616
rect 5479 23613 5491 23647
rect 5433 23607 5491 23613
rect 7374 23576 7380 23588
rect 7335 23548 7380 23576
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 7469 23579 7527 23585
rect 7469 23545 7481 23579
rect 7515 23576 7527 23579
rect 7742 23576 7748 23588
rect 7515 23548 7748 23576
rect 7515 23545 7527 23548
rect 7469 23539 7527 23545
rect 5353 23511 5411 23517
rect 5353 23477 5365 23511
rect 5399 23508 5411 23511
rect 5534 23508 5540 23520
rect 5399 23480 5540 23508
rect 5399 23477 5411 23480
rect 5353 23471 5411 23477
rect 5534 23468 5540 23480
rect 5592 23468 5598 23520
rect 6086 23508 6092 23520
rect 6047 23480 6092 23508
rect 6086 23468 6092 23480
rect 6144 23468 6150 23520
rect 7193 23511 7251 23517
rect 7193 23477 7205 23511
rect 7239 23508 7251 23511
rect 7484 23508 7512 23539
rect 7742 23536 7748 23548
rect 7800 23536 7806 23588
rect 8389 23579 8447 23585
rect 8389 23576 8401 23579
rect 7944 23548 8401 23576
rect 7944 23520 7972 23548
rect 8389 23545 8401 23548
rect 8435 23576 8447 23579
rect 8941 23579 8999 23585
rect 8941 23576 8953 23579
rect 8435 23548 8953 23576
rect 8435 23545 8447 23548
rect 8389 23539 8447 23545
rect 8941 23545 8953 23548
rect 8987 23545 8999 23579
rect 8941 23539 8999 23545
rect 9033 23579 9091 23585
rect 9033 23545 9045 23579
rect 9079 23545 9091 23579
rect 9033 23539 9091 23545
rect 10321 23579 10379 23585
rect 10321 23545 10333 23579
rect 10367 23576 10379 23579
rect 10704 23576 10732 23684
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 12710 23672 12716 23724
rect 12768 23712 12774 23724
rect 13170 23712 13176 23724
rect 12768 23684 13176 23712
rect 12768 23672 12774 23684
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23712 13875 23715
rect 14384 23712 14412 23752
rect 13863 23684 14412 23712
rect 13863 23681 13875 23684
rect 13817 23675 13875 23681
rect 14458 23672 14464 23724
rect 14516 23712 14522 23724
rect 15028 23721 15056 23752
rect 18325 23749 18337 23783
rect 18371 23780 18383 23783
rect 20070 23780 20076 23792
rect 18371 23752 20076 23780
rect 18371 23749 18383 23752
rect 18325 23743 18383 23749
rect 20070 23740 20076 23752
rect 20128 23740 20134 23792
rect 23845 23783 23903 23789
rect 23845 23749 23857 23783
rect 23891 23780 23903 23783
rect 25038 23780 25044 23792
rect 23891 23752 25044 23780
rect 23891 23749 23903 23752
rect 23845 23743 23903 23749
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 14516 23684 14749 23712
rect 14516 23672 14522 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 15013 23715 15071 23721
rect 15013 23681 15025 23715
rect 15059 23712 15071 23715
rect 16390 23712 16396 23724
rect 15059 23684 16396 23712
rect 15059 23681 15071 23684
rect 15013 23675 15071 23681
rect 16390 23672 16396 23684
rect 16448 23712 16454 23724
rect 16577 23715 16635 23721
rect 16577 23712 16589 23715
rect 16448 23684 16589 23712
rect 16448 23672 16454 23684
rect 16577 23681 16589 23684
rect 16623 23681 16635 23715
rect 16577 23675 16635 23681
rect 19518 23672 19524 23724
rect 19576 23712 19582 23724
rect 19797 23715 19855 23721
rect 19797 23712 19809 23715
rect 19576 23684 19809 23712
rect 19576 23672 19582 23684
rect 19797 23681 19809 23684
rect 19843 23681 19855 23715
rect 19797 23675 19855 23681
rect 19996 23684 20116 23712
rect 16482 23604 16488 23656
rect 16540 23644 16546 23656
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 16540 23616 16865 23644
rect 16540 23604 16546 23616
rect 16853 23613 16865 23616
rect 16899 23644 16911 23647
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16899 23616 17417 23644
rect 16899 23613 16911 23616
rect 16853 23607 16911 23613
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 18138 23644 18144 23656
rect 18051 23616 18144 23644
rect 17405 23607 17463 23613
rect 18138 23604 18144 23616
rect 18196 23644 18202 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18196 23616 18705 23644
rect 18196 23604 18202 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 19242 23644 19248 23656
rect 19203 23616 19248 23644
rect 18693 23607 18751 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 10873 23579 10931 23585
rect 10873 23576 10885 23579
rect 10367 23548 10885 23576
rect 10367 23545 10379 23548
rect 10321 23539 10379 23545
rect 10873 23545 10885 23548
rect 10919 23545 10931 23579
rect 10873 23539 10931 23545
rect 10965 23579 11023 23585
rect 10965 23545 10977 23579
rect 11011 23545 11023 23579
rect 11514 23576 11520 23588
rect 11475 23548 11520 23576
rect 10965 23539 11023 23545
rect 7239 23480 7512 23508
rect 7239 23477 7251 23480
rect 7193 23471 7251 23477
rect 7926 23468 7932 23520
rect 7984 23468 7990 23520
rect 8846 23468 8852 23520
rect 8904 23508 8910 23520
rect 9048 23508 9076 23539
rect 8904 23480 9076 23508
rect 8904 23468 8910 23480
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 10980 23508 11008 23539
rect 11514 23536 11520 23548
rect 11572 23536 11578 23588
rect 13265 23579 13323 23585
rect 13265 23545 13277 23579
rect 13311 23576 13323 23579
rect 13311 23548 13814 23576
rect 13311 23545 13323 23548
rect 13265 23539 13323 23545
rect 10836 23480 11008 23508
rect 12989 23511 13047 23517
rect 10836 23468 10842 23480
rect 12989 23477 13001 23511
rect 13035 23508 13047 23511
rect 13280 23508 13308 23539
rect 13035 23480 13308 23508
rect 13786 23508 13814 23548
rect 14366 23536 14372 23588
rect 14424 23576 14430 23588
rect 14829 23579 14887 23585
rect 14829 23576 14841 23579
rect 14424 23548 14841 23576
rect 14424 23536 14430 23548
rect 14829 23545 14841 23548
rect 14875 23545 14887 23579
rect 14829 23539 14887 23545
rect 14918 23536 14924 23588
rect 14976 23576 14982 23588
rect 19996 23576 20024 23684
rect 20088 23644 20116 23684
rect 20384 23647 20442 23653
rect 20384 23644 20396 23647
rect 20088 23616 20396 23644
rect 20384 23613 20396 23616
rect 20430 23644 20442 23647
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20430 23616 20821 23644
rect 20430 23613 20442 23616
rect 20384 23607 20442 23613
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 20809 23607 20867 23613
rect 21412 23647 21470 23653
rect 21412 23613 21424 23647
rect 21458 23644 21470 23647
rect 21726 23644 21732 23656
rect 21458 23616 21732 23644
rect 21458 23613 21470 23616
rect 21412 23607 21470 23613
rect 21726 23604 21732 23616
rect 21784 23644 21790 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21784 23616 21833 23644
rect 21784 23604 21790 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 22152 23616 23673 23644
rect 22152 23604 22158 23616
rect 23661 23613 23673 23616
rect 23707 23644 23719 23647
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23707 23616 24225 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 24765 23647 24823 23653
rect 24765 23613 24777 23647
rect 24811 23613 24823 23647
rect 24765 23607 24823 23613
rect 14976 23548 20024 23576
rect 14976 23536 14982 23548
rect 20070 23536 20076 23588
rect 20128 23576 20134 23588
rect 21499 23579 21557 23585
rect 21499 23576 21511 23579
rect 20128 23548 21511 23576
rect 20128 23536 20134 23548
rect 21499 23545 21511 23548
rect 21545 23545 21557 23579
rect 21499 23539 21557 23545
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 24780 23576 24808 23607
rect 25317 23579 25375 23585
rect 25317 23576 25329 23579
rect 23532 23548 25329 23576
rect 23532 23536 23538 23548
rect 25317 23545 25329 23548
rect 25363 23545 25375 23579
rect 25317 23539 25375 23545
rect 14090 23508 14096 23520
rect 13786 23480 14096 23508
rect 13035 23477 13047 23480
rect 12989 23471 13047 23477
rect 14090 23468 14096 23480
rect 14148 23468 14154 23520
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 20487 23511 20545 23517
rect 20487 23508 20499 23511
rect 20036 23480 20499 23508
rect 20036 23468 20042 23480
rect 20487 23477 20499 23480
rect 20533 23477 20545 23511
rect 20487 23471 20545 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2222 23304 2228 23316
rect 2183 23276 2228 23304
rect 2222 23264 2228 23276
rect 2280 23264 2286 23316
rect 3142 23264 3148 23316
rect 3200 23304 3206 23316
rect 4249 23307 4307 23313
rect 4249 23304 4261 23307
rect 3200 23276 4261 23304
rect 3200 23264 3206 23276
rect 4249 23273 4261 23276
rect 4295 23273 4307 23307
rect 4249 23267 4307 23273
rect 14458 23264 14464 23316
rect 14516 23304 14522 23316
rect 14737 23307 14795 23313
rect 14737 23304 14749 23307
rect 14516 23276 14749 23304
rect 14516 23264 14522 23276
rect 14737 23273 14749 23276
rect 14783 23304 14795 23307
rect 16942 23304 16948 23316
rect 14783 23276 16948 23304
rect 14783 23273 14795 23276
rect 14737 23267 14795 23273
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 17359 23307 17417 23313
rect 17359 23273 17371 23307
rect 17405 23304 17417 23307
rect 18138 23304 18144 23316
rect 17405 23276 18144 23304
rect 17405 23273 17417 23276
rect 17359 23267 17417 23273
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 18371 23307 18429 23313
rect 18371 23273 18383 23307
rect 18417 23304 18429 23307
rect 19242 23304 19248 23316
rect 18417 23276 19248 23304
rect 18417 23273 18429 23276
rect 18371 23267 18429 23273
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 5899 23239 5957 23245
rect 5899 23205 5911 23239
rect 5945 23236 5957 23239
rect 6270 23236 6276 23248
rect 5945 23208 6276 23236
rect 5945 23205 5957 23208
rect 5899 23199 5957 23205
rect 6270 23196 6276 23208
rect 6328 23196 6334 23248
rect 8202 23236 8208 23248
rect 8163 23208 8208 23236
rect 8202 23196 8208 23208
rect 8260 23236 8266 23248
rect 8478 23236 8484 23248
rect 8260 23208 8484 23236
rect 8260 23196 8266 23208
rect 8478 23196 8484 23208
rect 8536 23196 8542 23248
rect 8757 23239 8815 23245
rect 8757 23205 8769 23239
rect 8803 23236 8815 23239
rect 9214 23236 9220 23248
rect 8803 23208 9220 23236
rect 8803 23205 8815 23208
rect 8757 23199 8815 23205
rect 9214 23196 9220 23208
rect 9272 23196 9278 23248
rect 10597 23239 10655 23245
rect 10597 23205 10609 23239
rect 10643 23236 10655 23239
rect 10870 23236 10876 23248
rect 10643 23208 10876 23236
rect 10643 23205 10655 23208
rect 10597 23199 10655 23205
rect 10870 23196 10876 23208
rect 10928 23196 10934 23248
rect 11149 23239 11207 23245
rect 11149 23205 11161 23239
rect 11195 23236 11207 23239
rect 11514 23236 11520 23248
rect 11195 23208 11520 23236
rect 11195 23205 11207 23208
rect 11149 23199 11207 23205
rect 11514 23196 11520 23208
rect 11572 23196 11578 23248
rect 12161 23239 12219 23245
rect 12161 23205 12173 23239
rect 12207 23236 12219 23239
rect 12434 23236 12440 23248
rect 12207 23208 12440 23236
rect 12207 23205 12219 23208
rect 12161 23199 12219 23205
rect 12434 23196 12440 23208
rect 12492 23196 12498 23248
rect 12710 23236 12716 23248
rect 12671 23208 12716 23236
rect 12710 23196 12716 23208
rect 12768 23196 12774 23248
rect 13817 23239 13875 23245
rect 13817 23205 13829 23239
rect 13863 23236 13875 23239
rect 14182 23236 14188 23248
rect 13863 23208 14188 23236
rect 13863 23205 13875 23208
rect 13817 23199 13875 23205
rect 14182 23196 14188 23208
rect 14240 23196 14246 23248
rect 2590 23168 2596 23180
rect 2551 23140 2596 23168
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 4065 23171 4123 23177
rect 4065 23137 4077 23171
rect 4111 23168 4123 23171
rect 4522 23168 4528 23180
rect 4111 23140 4528 23168
rect 4111 23137 4123 23140
rect 4065 23131 4123 23137
rect 4522 23128 4528 23140
rect 4580 23128 4586 23180
rect 14918 23168 14924 23180
rect 14660 23140 14924 23168
rect 3602 23060 3608 23112
rect 3660 23100 3666 23112
rect 5537 23103 5595 23109
rect 3660 23072 4154 23100
rect 3660 23060 3666 23072
rect 4126 23032 4154 23072
rect 5537 23069 5549 23103
rect 5583 23100 5595 23103
rect 5994 23100 6000 23112
rect 5583 23072 6000 23100
rect 5583 23069 5595 23072
rect 5537 23063 5595 23069
rect 5994 23060 6000 23072
rect 6052 23060 6058 23112
rect 8110 23100 8116 23112
rect 8023 23072 8116 23100
rect 8110 23060 8116 23072
rect 8168 23100 8174 23112
rect 9582 23100 9588 23112
rect 8168 23072 9588 23100
rect 8168 23060 8174 23072
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23100 10563 23103
rect 10686 23100 10692 23112
rect 10551 23072 10692 23100
rect 10551 23069 10563 23072
rect 10505 23063 10563 23069
rect 10686 23060 10692 23072
rect 10744 23100 10750 23112
rect 11425 23103 11483 23109
rect 11425 23100 11437 23103
rect 10744 23072 11437 23100
rect 10744 23060 10750 23072
rect 11425 23069 11437 23072
rect 11471 23069 11483 23103
rect 11425 23063 11483 23069
rect 11882 23060 11888 23112
rect 11940 23100 11946 23112
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 11940 23072 12081 23100
rect 11940 23060 11946 23072
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 13722 23100 13728 23112
rect 13683 23072 13728 23100
rect 12069 23063 12127 23069
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 14660 23100 14688 23140
rect 14918 23128 14924 23140
rect 14976 23128 14982 23180
rect 15654 23168 15660 23180
rect 15615 23140 15660 23168
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 17218 23168 17224 23180
rect 17179 23140 17224 23168
rect 17218 23128 17224 23140
rect 17276 23128 17282 23180
rect 18268 23171 18326 23177
rect 18268 23137 18280 23171
rect 18314 23137 18326 23171
rect 18268 23131 18326 23137
rect 19312 23171 19370 23177
rect 19312 23137 19324 23171
rect 19358 23168 19370 23171
rect 19886 23168 19892 23180
rect 19358 23140 19892 23168
rect 19358 23137 19370 23140
rect 19312 23131 19370 23137
rect 14200 23072 14688 23100
rect 6825 23035 6883 23041
rect 6825 23032 6837 23035
rect 4126 23004 6837 23032
rect 6825 23001 6837 23004
rect 6871 23032 6883 23035
rect 7190 23032 7196 23044
rect 6871 23004 7196 23032
rect 6871 23001 6883 23004
rect 6825 22995 6883 23001
rect 7190 22992 7196 23004
rect 7248 22992 7254 23044
rect 8938 22992 8944 23044
rect 8996 23032 9002 23044
rect 14200 23032 14228 23072
rect 14826 23060 14832 23112
rect 14884 23100 14890 23112
rect 15289 23103 15347 23109
rect 15289 23100 15301 23103
rect 14884 23072 15301 23100
rect 14884 23060 14890 23072
rect 15289 23069 15301 23072
rect 15335 23069 15347 23103
rect 15289 23063 15347 23069
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 18283 23100 18311 23131
rect 19886 23128 19892 23140
rect 19944 23128 19950 23180
rect 18874 23100 18880 23112
rect 16724 23072 18880 23100
rect 16724 23060 16730 23072
rect 18874 23060 18880 23072
rect 18932 23060 18938 23112
rect 8996 23004 14228 23032
rect 8996 22992 9002 23004
rect 14274 22992 14280 23044
rect 14332 23032 14338 23044
rect 14332 23004 14377 23032
rect 14332 22992 14338 23004
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 1854 22924 1860 22976
rect 1912 22964 1918 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 1912 22936 3065 22964
rect 1912 22924 1918 22936
rect 3053 22933 3065 22936
rect 3099 22964 3111 22967
rect 3326 22964 3332 22976
rect 3099 22936 3332 22964
rect 3099 22933 3111 22936
rect 3053 22927 3111 22933
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 5074 22964 5080 22976
rect 5035 22936 5080 22964
rect 5074 22924 5080 22936
rect 5132 22924 5138 22976
rect 5258 22924 5264 22976
rect 5316 22964 5322 22976
rect 6457 22967 6515 22973
rect 6457 22964 6469 22967
rect 5316 22936 6469 22964
rect 5316 22924 5322 22936
rect 6457 22933 6469 22936
rect 6503 22933 6515 22967
rect 7374 22964 7380 22976
rect 7335 22936 7380 22964
rect 6457 22927 6515 22933
rect 7374 22924 7380 22936
rect 7432 22924 7438 22976
rect 7929 22967 7987 22973
rect 7929 22933 7941 22967
rect 7975 22964 7987 22967
rect 8294 22964 8300 22976
rect 7975 22936 8300 22964
rect 7975 22933 7987 22936
rect 7929 22927 7987 22933
rect 8294 22924 8300 22936
rect 8352 22964 8358 22976
rect 8754 22964 8760 22976
rect 8352 22936 8760 22964
rect 8352 22924 8358 22936
rect 8754 22924 8760 22936
rect 8812 22924 8818 22976
rect 9766 22924 9772 22976
rect 9824 22964 9830 22976
rect 9953 22967 10011 22973
rect 9953 22964 9965 22967
rect 9824 22936 9965 22964
rect 9824 22924 9830 22936
rect 9953 22933 9965 22936
rect 9999 22933 10011 22967
rect 12986 22964 12992 22976
rect 12947 22936 12992 22964
rect 9953 22927 10011 22933
rect 12986 22924 12992 22936
rect 13044 22924 13050 22976
rect 16390 22964 16396 22976
rect 16351 22936 16396 22964
rect 16390 22924 16396 22936
rect 16448 22924 16454 22976
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 19383 22967 19441 22973
rect 19383 22964 19395 22967
rect 18104 22936 19395 22964
rect 18104 22924 18110 22936
rect 19383 22933 19395 22936
rect 19429 22933 19441 22967
rect 19383 22927 19441 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2590 22720 2596 22772
rect 2648 22760 2654 22772
rect 2961 22763 3019 22769
rect 2961 22760 2973 22763
rect 2648 22732 2973 22760
rect 2648 22720 2654 22732
rect 2961 22729 2973 22732
rect 3007 22760 3019 22763
rect 5258 22760 5264 22772
rect 3007 22732 5264 22760
rect 3007 22729 3019 22732
rect 2961 22723 3019 22729
rect 5258 22720 5264 22732
rect 5316 22720 5322 22772
rect 5905 22763 5963 22769
rect 5905 22729 5917 22763
rect 5951 22760 5963 22763
rect 6086 22760 6092 22772
rect 5951 22732 6092 22760
rect 5951 22729 5963 22732
rect 5905 22723 5963 22729
rect 6086 22720 6092 22732
rect 6144 22720 6150 22772
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8202 22760 8208 22772
rect 7975 22732 8208 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8202 22720 8208 22732
rect 8260 22760 8266 22772
rect 9309 22763 9367 22769
rect 9309 22760 9321 22763
rect 8260 22732 9321 22760
rect 8260 22720 8266 22732
rect 9309 22729 9321 22732
rect 9355 22729 9367 22763
rect 9582 22760 9588 22772
rect 9543 22732 9588 22760
rect 9309 22723 9367 22729
rect 9582 22720 9588 22732
rect 9640 22720 9646 22772
rect 10042 22760 10048 22772
rect 10003 22732 10048 22760
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 12069 22763 12127 22769
rect 12069 22729 12081 22763
rect 12115 22760 12127 22763
rect 12434 22760 12440 22772
rect 12115 22732 12440 22760
rect 12115 22729 12127 22732
rect 12069 22723 12127 22729
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 13817 22763 13875 22769
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 14090 22760 14096 22772
rect 13863 22732 14096 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 14182 22720 14188 22772
rect 14240 22760 14246 22772
rect 15654 22760 15660 22772
rect 14240 22732 15660 22760
rect 14240 22720 14246 22732
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 17218 22760 17224 22772
rect 16361 22732 17224 22760
rect 2866 22692 2872 22704
rect 1964 22664 2872 22692
rect 1964 22633 1992 22664
rect 2866 22652 2872 22664
rect 2924 22652 2930 22704
rect 4890 22652 4896 22704
rect 4948 22692 4954 22704
rect 11517 22695 11575 22701
rect 11517 22692 11529 22695
rect 4948 22664 11529 22692
rect 4948 22652 4954 22664
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22593 2007 22627
rect 2314 22624 2320 22636
rect 2275 22596 2320 22624
rect 1949 22587 2007 22593
rect 2314 22584 2320 22596
rect 2372 22584 2378 22636
rect 10244 22633 10272 22664
rect 11517 22661 11529 22664
rect 11563 22661 11575 22695
rect 11517 22655 11575 22661
rect 11606 22652 11612 22704
rect 11664 22692 11670 22704
rect 16361 22692 16389 22732
rect 17218 22720 17224 22732
rect 17276 22760 17282 22772
rect 17313 22763 17371 22769
rect 17313 22760 17325 22763
rect 17276 22732 17325 22760
rect 17276 22720 17282 22732
rect 17313 22729 17325 22732
rect 17359 22729 17371 22763
rect 18874 22760 18880 22772
rect 18835 22732 18880 22760
rect 17313 22723 17371 22729
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 19058 22720 19064 22772
rect 19116 22760 19122 22772
rect 19199 22763 19257 22769
rect 19199 22760 19211 22763
rect 19116 22732 19211 22760
rect 19116 22720 19122 22732
rect 19199 22729 19211 22732
rect 19245 22729 19257 22763
rect 19886 22760 19892 22772
rect 19847 22732 19892 22760
rect 19199 22723 19257 22729
rect 19886 22720 19892 22732
rect 19944 22720 19950 22772
rect 11664 22664 16389 22692
rect 11664 22652 11670 22664
rect 16482 22652 16488 22704
rect 16540 22692 16546 22704
rect 16540 22664 19334 22692
rect 16540 22652 16546 22664
rect 6457 22627 6515 22633
rect 6457 22593 6469 22627
rect 6503 22624 6515 22627
rect 10229 22627 10287 22633
rect 6503 22596 6868 22624
rect 6503 22593 6515 22596
rect 6457 22587 6515 22593
rect 3329 22559 3387 22565
rect 3329 22525 3341 22559
rect 3375 22556 3387 22559
rect 3694 22556 3700 22568
rect 3375 22528 3700 22556
rect 3375 22525 3387 22528
rect 3329 22519 3387 22525
rect 3694 22516 3700 22528
rect 3752 22516 3758 22568
rect 3881 22559 3939 22565
rect 3881 22525 3893 22559
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 4798 22556 4804 22568
rect 4203 22528 4804 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 1765 22491 1823 22497
rect 1765 22457 1777 22491
rect 1811 22488 1823 22491
rect 2041 22491 2099 22497
rect 2041 22488 2053 22491
rect 1811 22460 2053 22488
rect 1811 22457 1823 22460
rect 1765 22451 1823 22457
rect 2041 22457 2053 22460
rect 2087 22488 2099 22491
rect 2314 22488 2320 22500
rect 2087 22460 2320 22488
rect 2087 22457 2099 22460
rect 2041 22451 2099 22457
rect 2314 22448 2320 22460
rect 2372 22448 2378 22500
rect 3602 22448 3608 22500
rect 3660 22488 3666 22500
rect 3896 22488 3924 22519
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 4985 22559 5043 22565
rect 4985 22525 4997 22559
rect 5031 22556 5043 22559
rect 5074 22556 5080 22568
rect 5031 22528 5080 22556
rect 5031 22525 5043 22528
rect 4985 22519 5043 22525
rect 5074 22516 5080 22528
rect 5132 22556 5138 22568
rect 6840 22565 6868 22596
rect 10229 22593 10241 22627
rect 10275 22593 10287 22627
rect 10686 22624 10692 22636
rect 10647 22596 10692 22624
rect 10229 22587 10287 22593
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 14274 22584 14280 22636
rect 14332 22624 14338 22636
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14332 22596 15025 22624
rect 14332 22584 14338 22596
rect 15013 22593 15025 22596
rect 15059 22624 15071 22627
rect 15470 22624 15476 22636
rect 15059 22596 15476 22624
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 15470 22584 15476 22596
rect 15528 22584 15534 22636
rect 16666 22624 16672 22636
rect 16627 22596 16672 22624
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 19306 22624 19334 22664
rect 20073 22627 20131 22633
rect 20073 22624 20085 22627
rect 19306 22596 20085 22624
rect 20073 22593 20085 22596
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 6825 22559 6883 22565
rect 5132 22528 6684 22556
rect 5132 22516 5138 22528
rect 3660 22460 3924 22488
rect 5347 22491 5405 22497
rect 3660 22448 3666 22460
rect 5347 22457 5359 22491
rect 5393 22457 5405 22491
rect 5347 22451 5405 22457
rect 4522 22420 4528 22432
rect 4483 22392 4528 22420
rect 4522 22380 4528 22392
rect 4580 22380 4586 22432
rect 4893 22423 4951 22429
rect 4893 22389 4905 22423
rect 4939 22420 4951 22423
rect 5074 22420 5080 22432
rect 4939 22392 5080 22420
rect 4939 22389 4951 22392
rect 4893 22383 4951 22389
rect 5074 22380 5080 22392
rect 5132 22420 5138 22432
rect 5368 22420 5396 22451
rect 5442 22448 5448 22500
rect 5500 22488 5506 22500
rect 6457 22491 6515 22497
rect 6457 22488 6469 22491
rect 5500 22460 6469 22488
rect 5500 22448 5506 22460
rect 6457 22457 6469 22460
rect 6503 22488 6515 22491
rect 6549 22491 6607 22497
rect 6549 22488 6561 22491
rect 6503 22460 6561 22488
rect 6503 22457 6515 22460
rect 6457 22451 6515 22457
rect 6549 22457 6561 22460
rect 6595 22457 6607 22491
rect 6549 22451 6607 22457
rect 6270 22420 6276 22432
rect 5132 22392 6276 22420
rect 5132 22380 5138 22392
rect 6270 22380 6276 22392
rect 6328 22380 6334 22432
rect 6656 22420 6684 22528
rect 6825 22525 6837 22559
rect 6871 22525 6883 22559
rect 6825 22519 6883 22525
rect 7190 22516 7196 22568
rect 7248 22556 7254 22568
rect 7285 22559 7343 22565
rect 7285 22556 7297 22559
rect 7248 22528 7297 22556
rect 7248 22516 7254 22528
rect 7285 22525 7297 22528
rect 7331 22525 7343 22559
rect 7285 22519 7343 22525
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22556 8447 22559
rect 9030 22556 9036 22568
rect 8435 22528 9036 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 9030 22516 9036 22528
rect 9088 22516 9094 22568
rect 12250 22516 12256 22568
rect 12308 22556 12314 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12308 22528 12909 22556
rect 12308 22516 12314 22528
rect 12897 22525 12909 22528
rect 12943 22556 12955 22559
rect 12986 22556 12992 22568
rect 12943 22528 12992 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 12986 22516 12992 22528
rect 13044 22516 13050 22568
rect 18116 22559 18174 22565
rect 18116 22525 18128 22559
rect 18162 22556 18174 22559
rect 18506 22556 18512 22568
rect 18162 22528 18512 22556
rect 18162 22525 18174 22528
rect 18116 22519 18174 22525
rect 18506 22516 18512 22528
rect 18564 22516 18570 22568
rect 19128 22559 19186 22565
rect 19128 22525 19140 22559
rect 19174 22556 19186 22559
rect 19518 22556 19524 22568
rect 19174 22528 19524 22556
rect 19174 22525 19186 22528
rect 19128 22519 19186 22525
rect 19518 22516 19524 22528
rect 19576 22516 19582 22568
rect 8297 22491 8355 22497
rect 8297 22457 8309 22491
rect 8343 22488 8355 22491
rect 8751 22491 8809 22497
rect 8751 22488 8763 22491
rect 8343 22460 8763 22488
rect 8343 22457 8355 22460
rect 8297 22451 8355 22457
rect 8751 22457 8763 22460
rect 8797 22488 8809 22491
rect 8846 22488 8852 22500
rect 8797 22460 8852 22488
rect 8797 22457 8809 22460
rect 8751 22451 8809 22457
rect 8846 22448 8852 22460
rect 8904 22448 8910 22500
rect 10321 22491 10379 22497
rect 10321 22457 10333 22491
rect 10367 22457 10379 22491
rect 14734 22488 14740 22500
rect 14695 22460 14740 22488
rect 10321 22451 10379 22457
rect 6917 22423 6975 22429
rect 6917 22420 6929 22423
rect 6656 22392 6929 22420
rect 6917 22389 6929 22392
rect 6963 22389 6975 22423
rect 6917 22383 6975 22389
rect 10042 22380 10048 22432
rect 10100 22420 10106 22432
rect 10336 22420 10364 22451
rect 14734 22448 14740 22460
rect 14792 22448 14798 22500
rect 14826 22448 14832 22500
rect 14884 22488 14890 22500
rect 16390 22488 16396 22500
rect 14884 22460 14929 22488
rect 16351 22460 16396 22488
rect 14884 22448 14890 22460
rect 16390 22448 16396 22460
rect 16448 22448 16454 22500
rect 16482 22448 16488 22500
rect 16540 22488 16546 22500
rect 16540 22460 16585 22488
rect 16540 22448 16546 22460
rect 10100 22392 10364 22420
rect 10100 22380 10106 22392
rect 10870 22380 10876 22432
rect 10928 22420 10934 22432
rect 11238 22420 11244 22432
rect 10928 22392 11244 22420
rect 10928 22380 10934 22392
rect 11238 22380 11244 22392
rect 11296 22380 11302 22432
rect 12802 22420 12808 22432
rect 12715 22392 12808 22420
rect 12802 22380 12808 22392
rect 12860 22420 12866 22432
rect 13265 22423 13323 22429
rect 13265 22420 13277 22423
rect 12860 22392 13277 22420
rect 12860 22380 12866 22392
rect 13265 22389 13277 22392
rect 13311 22389 13323 22423
rect 13265 22383 13323 22389
rect 14553 22423 14611 22429
rect 14553 22389 14565 22423
rect 14599 22420 14611 22423
rect 14844 22420 14872 22448
rect 14599 22392 14872 22420
rect 16209 22423 16267 22429
rect 14599 22389 14611 22392
rect 14553 22383 14611 22389
rect 16209 22389 16221 22423
rect 16255 22420 16267 22423
rect 16500 22420 16528 22448
rect 16255 22392 16528 22420
rect 16255 22389 16267 22392
rect 16209 22383 16267 22389
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 18187 22423 18245 22429
rect 18187 22420 18199 22423
rect 16632 22392 18199 22420
rect 16632 22380 16638 22392
rect 18187 22389 18199 22392
rect 18233 22389 18245 22423
rect 19518 22420 19524 22432
rect 19479 22392 19524 22420
rect 18187 22383 18245 22389
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 2866 22216 2872 22228
rect 2823 22188 2872 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 2866 22176 2872 22188
rect 2924 22176 2930 22228
rect 4982 22176 4988 22228
rect 5040 22216 5046 22228
rect 5721 22219 5779 22225
rect 5721 22216 5733 22219
rect 5040 22188 5733 22216
rect 5040 22176 5046 22188
rect 5721 22185 5733 22188
rect 5767 22185 5779 22219
rect 5721 22179 5779 22185
rect 6825 22219 6883 22225
rect 6825 22185 6837 22219
rect 6871 22216 6883 22219
rect 7926 22216 7932 22228
rect 6871 22188 7932 22216
rect 6871 22185 6883 22188
rect 6825 22179 6883 22185
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 8754 22216 8760 22228
rect 8715 22188 8760 22216
rect 8754 22176 8760 22188
rect 8812 22176 8818 22228
rect 11238 22216 11244 22228
rect 11199 22188 11244 22216
rect 11238 22176 11244 22188
rect 11296 22176 11302 22228
rect 12158 22176 12164 22228
rect 12216 22216 12222 22228
rect 12989 22219 13047 22225
rect 12989 22216 13001 22219
rect 12216 22188 13001 22216
rect 12216 22176 12222 22188
rect 12989 22185 13001 22188
rect 13035 22185 13047 22219
rect 13722 22216 13728 22228
rect 13683 22188 13728 22216
rect 12989 22179 13047 22185
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 14734 22216 14740 22228
rect 14695 22188 14740 22216
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 15470 22216 15476 22228
rect 15431 22188 15476 22216
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 22649 22219 22707 22225
rect 22649 22185 22661 22219
rect 22695 22216 22707 22219
rect 24210 22216 24216 22228
rect 22695 22188 24216 22216
rect 22695 22185 22707 22188
rect 22649 22179 22707 22185
rect 24210 22176 24216 22188
rect 24268 22176 24274 22228
rect 1670 22148 1676 22160
rect 1631 22120 1676 22148
rect 1670 22108 1676 22120
rect 1728 22108 1734 22160
rect 5160 22108 5166 22160
rect 5218 22148 5224 22160
rect 5218 22120 5263 22148
rect 5218 22108 5224 22120
rect 6270 22108 6276 22160
rect 6328 22148 6334 22160
rect 6454 22148 6460 22160
rect 6328 22120 6460 22148
rect 6328 22108 6334 22120
rect 6454 22108 6460 22120
rect 6512 22148 6518 22160
rect 8018 22148 8024 22160
rect 6512 22120 8024 22148
rect 6512 22108 6518 22120
rect 8018 22108 8024 22120
rect 8076 22148 8082 22160
rect 8199 22151 8257 22157
rect 8199 22148 8211 22151
rect 8076 22120 8211 22148
rect 8076 22108 8082 22120
rect 8199 22117 8211 22120
rect 8245 22148 8257 22151
rect 8846 22148 8852 22160
rect 8245 22120 8852 22148
rect 8245 22117 8257 22120
rect 8199 22111 8257 22117
rect 8846 22108 8852 22120
rect 8904 22148 8910 22160
rect 10410 22148 10416 22160
rect 8904 22120 10416 22148
rect 8904 22108 8910 22120
rect 10410 22108 10416 22120
rect 10468 22148 10474 22160
rect 10683 22151 10741 22157
rect 10683 22148 10695 22151
rect 10468 22120 10695 22148
rect 10468 22108 10474 22120
rect 10683 22117 10695 22120
rect 10729 22148 10741 22151
rect 12431 22151 12489 22157
rect 12431 22148 12443 22151
rect 10729 22120 12443 22148
rect 10729 22117 10741 22120
rect 10683 22111 10741 22117
rect 12431 22117 12443 22120
rect 12477 22148 12489 22151
rect 12802 22148 12808 22160
rect 12477 22120 12808 22148
rect 12477 22117 12489 22120
rect 12431 22111 12489 22117
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 15488 22148 15516 22176
rect 15749 22151 15807 22157
rect 15749 22148 15761 22151
rect 15488 22120 15761 22148
rect 15749 22117 15761 22120
rect 15795 22117 15807 22151
rect 15749 22111 15807 22117
rect 15841 22151 15899 22157
rect 15841 22117 15853 22151
rect 15887 22148 15899 22151
rect 15930 22148 15936 22160
rect 15887 22120 15936 22148
rect 15887 22117 15899 22120
rect 15841 22111 15899 22117
rect 15930 22108 15936 22120
rect 15988 22108 15994 22160
rect 16393 22151 16451 22157
rect 16393 22117 16405 22151
rect 16439 22148 16451 22151
rect 16666 22148 16672 22160
rect 16439 22120 16672 22148
rect 16439 22117 16451 22120
rect 16393 22111 16451 22117
rect 16666 22108 16672 22120
rect 16724 22108 16730 22160
rect 2314 22080 2320 22092
rect 2275 22052 2320 22080
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 9950 22040 9956 22092
rect 10008 22080 10014 22092
rect 11882 22080 11888 22092
rect 10008 22052 11888 22080
rect 10008 22040 10014 22052
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 14090 22040 14096 22092
rect 14148 22080 14154 22092
rect 14252 22083 14310 22089
rect 14252 22080 14264 22083
rect 14148 22052 14264 22080
rect 14148 22040 14154 22052
rect 14252 22049 14264 22052
rect 14298 22080 14310 22083
rect 15562 22080 15568 22092
rect 14298 22052 15568 22080
rect 14298 22049 14310 22052
rect 14252 22043 14310 22049
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 17126 22040 17132 22092
rect 17184 22080 17190 22092
rect 17256 22083 17314 22089
rect 17256 22080 17268 22083
rect 17184 22052 17268 22080
rect 17184 22040 17190 22052
rect 17256 22049 17268 22052
rect 17302 22049 17314 22083
rect 17256 22043 17314 22049
rect 18300 22083 18358 22089
rect 18300 22049 18312 22083
rect 18346 22080 18358 22083
rect 18414 22080 18420 22092
rect 18346 22052 18420 22080
rect 18346 22049 18358 22052
rect 18300 22043 18358 22049
rect 18414 22040 18420 22052
rect 18472 22040 18478 22092
rect 19312 22083 19370 22089
rect 19312 22049 19324 22083
rect 19358 22080 19370 22083
rect 19518 22080 19524 22092
rect 19358 22052 19524 22080
rect 19358 22049 19370 22052
rect 19312 22043 19370 22049
rect 19518 22040 19524 22052
rect 19576 22040 19582 22092
rect 21358 22080 21364 22092
rect 21319 22052 21364 22080
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 22462 22080 22468 22092
rect 22423 22052 22468 22080
rect 22462 22040 22468 22052
rect 22520 22040 22526 22092
rect 4798 22012 4804 22024
rect 4759 21984 4804 22012
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 7926 22012 7932 22024
rect 7883 21984 7932 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 7926 21972 7932 21984
rect 7984 21972 7990 22024
rect 10321 22015 10379 22021
rect 10321 22012 10333 22015
rect 10152 21984 10333 22012
rect 1854 21904 1860 21956
rect 1912 21944 1918 21956
rect 5350 21944 5356 21956
rect 1912 21916 5356 21944
rect 1912 21904 1918 21916
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 10152 21888 10180 21984
rect 10321 21981 10333 21984
rect 10367 21981 10379 22015
rect 10321 21975 10379 21981
rect 12069 22015 12127 22021
rect 12069 21981 12081 22015
rect 12115 22012 12127 22015
rect 12158 22012 12164 22024
rect 12115 21984 12164 22012
rect 12115 21981 12127 21984
rect 12069 21975 12127 21981
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 14734 22012 14740 22024
rect 12676 21984 14740 22012
rect 12676 21972 12682 21984
rect 14734 21972 14740 21984
rect 14792 21972 14798 22024
rect 12894 21904 12900 21956
rect 12952 21944 12958 21956
rect 13265 21947 13323 21953
rect 13265 21944 13277 21947
rect 12952 21916 13277 21944
rect 12952 21904 12958 21916
rect 13265 21913 13277 21916
rect 13311 21913 13323 21947
rect 13265 21907 13323 21913
rect 21545 21947 21603 21953
rect 21545 21913 21557 21947
rect 21591 21944 21603 21947
rect 23198 21944 23204 21956
rect 21591 21916 23204 21944
rect 21591 21913 21603 21916
rect 21545 21907 21603 21913
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 3513 21879 3571 21885
rect 3513 21845 3525 21879
rect 3559 21876 3571 21879
rect 3602 21876 3608 21888
rect 3559 21848 3608 21876
rect 3559 21845 3571 21848
rect 3513 21839 3571 21845
rect 3602 21836 3608 21848
rect 3660 21836 3666 21888
rect 5994 21876 6000 21888
rect 5955 21848 6000 21876
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 10134 21876 10140 21888
rect 10095 21848 10140 21876
rect 10134 21836 10140 21848
rect 10192 21836 10198 21888
rect 13630 21836 13636 21888
rect 13688 21876 13694 21888
rect 14323 21879 14381 21885
rect 14323 21876 14335 21879
rect 13688 21848 14335 21876
rect 13688 21836 13694 21848
rect 14323 21845 14335 21848
rect 14369 21845 14381 21879
rect 14323 21839 14381 21845
rect 15562 21836 15568 21888
rect 15620 21876 15626 21888
rect 17359 21879 17417 21885
rect 17359 21876 17371 21879
rect 15620 21848 17371 21876
rect 15620 21836 15626 21848
rect 17359 21845 17371 21848
rect 17405 21845 17417 21879
rect 17359 21839 17417 21845
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 18371 21879 18429 21885
rect 18371 21876 18383 21879
rect 17552 21848 18383 21876
rect 17552 21836 17558 21848
rect 18371 21845 18383 21848
rect 18417 21845 18429 21879
rect 18371 21839 18429 21845
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 19383 21879 19441 21885
rect 19383 21876 19395 21879
rect 18564 21848 19395 21876
rect 18564 21836 18570 21848
rect 19383 21845 19395 21848
rect 19429 21845 19441 21879
rect 19383 21839 19441 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2682 21632 2688 21684
rect 2740 21672 2746 21684
rect 3881 21675 3939 21681
rect 3881 21672 3893 21675
rect 2740 21644 3893 21672
rect 2740 21632 2746 21644
rect 3881 21641 3893 21644
rect 3927 21641 3939 21675
rect 3881 21635 3939 21641
rect 4798 21632 4804 21684
rect 4856 21672 4862 21684
rect 6181 21675 6239 21681
rect 6181 21672 6193 21675
rect 4856 21644 6193 21672
rect 4856 21632 4862 21644
rect 6181 21641 6193 21644
rect 6227 21641 6239 21675
rect 6181 21635 6239 21641
rect 7929 21675 7987 21681
rect 7929 21641 7941 21675
rect 7975 21672 7987 21675
rect 8018 21672 8024 21684
rect 7975 21644 8024 21672
rect 7975 21641 7987 21644
rect 7929 21635 7987 21641
rect 8018 21632 8024 21644
rect 8076 21632 8082 21684
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 9907 21675 9965 21681
rect 9907 21672 9919 21675
rect 9824 21644 9919 21672
rect 9824 21632 9830 21644
rect 9907 21641 9919 21644
rect 9953 21641 9965 21675
rect 10410 21672 10416 21684
rect 10371 21644 10416 21672
rect 9907 21635 9965 21641
rect 10410 21632 10416 21644
rect 10468 21672 10474 21684
rect 10686 21672 10692 21684
rect 10468 21644 10692 21672
rect 10468 21632 10474 21644
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 12161 21675 12219 21681
rect 12161 21641 12173 21675
rect 12207 21672 12219 21675
rect 12802 21672 12808 21684
rect 12207 21644 12808 21672
rect 12207 21641 12219 21644
rect 12161 21635 12219 21641
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 13817 21675 13875 21681
rect 13817 21641 13829 21675
rect 13863 21672 13875 21675
rect 14182 21672 14188 21684
rect 13863 21644 14188 21672
rect 13863 21641 13875 21644
rect 13817 21635 13875 21641
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 16482 21632 16488 21684
rect 16540 21672 16546 21684
rect 16669 21675 16727 21681
rect 16669 21672 16681 21675
rect 16540 21644 16681 21672
rect 16540 21632 16546 21644
rect 16669 21641 16681 21644
rect 16715 21641 16727 21675
rect 16669 21635 16727 21641
rect 17126 21632 17132 21684
rect 17184 21672 17190 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 17184 21644 17417 21672
rect 17184 21632 17190 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 1762 21564 1768 21616
rect 1820 21604 1826 21616
rect 2314 21604 2320 21616
rect 1820 21576 2320 21604
rect 1820 21564 1826 21576
rect 2314 21564 2320 21576
rect 2372 21604 2378 21616
rect 5905 21607 5963 21613
rect 5905 21604 5917 21607
rect 2372 21576 5917 21604
rect 2372 21564 2378 21576
rect 5905 21573 5917 21576
rect 5951 21573 5963 21607
rect 5905 21567 5963 21573
rect 9677 21607 9735 21613
rect 9677 21573 9689 21607
rect 9723 21604 9735 21607
rect 10962 21604 10968 21616
rect 9723 21576 10968 21604
rect 9723 21573 9735 21576
rect 9677 21567 9735 21573
rect 6638 21536 6644 21548
rect 4126 21508 6644 21536
rect 3605 21471 3663 21477
rect 3605 21437 3617 21471
rect 3651 21468 3663 21471
rect 3697 21471 3755 21477
rect 3697 21468 3709 21471
rect 3651 21440 3709 21468
rect 3651 21437 3663 21440
rect 3605 21431 3663 21437
rect 3697 21437 3709 21440
rect 3743 21468 3755 21471
rect 4126 21468 4154 21508
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 6822 21536 6828 21548
rect 6783 21508 6828 21536
rect 6822 21496 6828 21508
rect 6880 21496 6886 21548
rect 8404 21508 9352 21536
rect 3743 21440 4154 21468
rect 4985 21471 5043 21477
rect 3743 21437 3755 21440
rect 3697 21431 3755 21437
rect 4985 21437 4997 21471
rect 5031 21468 5043 21471
rect 5626 21468 5632 21480
rect 5031 21440 5632 21468
rect 5031 21437 5043 21440
rect 4985 21431 5043 21437
rect 5626 21428 5632 21440
rect 5684 21468 5690 21480
rect 8404 21477 8432 21508
rect 6549 21471 6607 21477
rect 6549 21468 6561 21471
rect 5684 21440 6561 21468
rect 5684 21428 5690 21440
rect 6549 21437 6561 21440
rect 6595 21437 6607 21471
rect 6549 21431 6607 21437
rect 8389 21471 8447 21477
rect 8389 21437 8401 21471
rect 8435 21437 8447 21471
rect 8389 21431 8447 21437
rect 8478 21428 8484 21480
rect 8536 21468 8542 21480
rect 8665 21471 8723 21477
rect 8665 21468 8677 21471
rect 8536 21440 8677 21468
rect 8536 21428 8542 21440
rect 8665 21437 8677 21440
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 1673 21403 1731 21409
rect 1673 21369 1685 21403
rect 1719 21400 1731 21403
rect 2222 21400 2228 21412
rect 1719 21372 2228 21400
rect 1719 21369 1731 21372
rect 1673 21363 1731 21369
rect 2222 21360 2228 21372
rect 2280 21360 2286 21412
rect 2314 21360 2320 21412
rect 2372 21400 2378 21412
rect 2866 21400 2872 21412
rect 2372 21372 2417 21400
rect 2827 21372 2872 21400
rect 2372 21360 2378 21372
rect 2866 21360 2872 21372
rect 2924 21360 2930 21412
rect 4525 21403 4583 21409
rect 4525 21369 4537 21403
rect 4571 21400 4583 21403
rect 4893 21403 4951 21409
rect 4893 21400 4905 21403
rect 4571 21372 4905 21400
rect 4571 21369 4583 21372
rect 4525 21363 4583 21369
rect 4893 21369 4905 21372
rect 4939 21400 4951 21403
rect 5074 21400 5080 21412
rect 4939 21372 5080 21400
rect 4939 21369 4951 21372
rect 4893 21363 4951 21369
rect 5074 21360 5080 21372
rect 5132 21400 5138 21412
rect 5306 21403 5364 21409
rect 5306 21400 5318 21403
rect 5132 21372 5318 21400
rect 5132 21360 5138 21372
rect 5306 21369 5318 21372
rect 5352 21369 5364 21403
rect 5306 21363 5364 21369
rect 7561 21403 7619 21409
rect 7561 21369 7573 21403
rect 7607 21400 7619 21403
rect 8496 21400 8524 21428
rect 9324 21409 9352 21508
rect 9851 21477 9879 21576
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 14090 21604 14096 21616
rect 14051 21576 14096 21604
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 19199 21607 19257 21613
rect 19199 21573 19211 21607
rect 19245 21604 19257 21607
rect 22462 21604 22468 21616
rect 19245 21576 22468 21604
rect 19245 21573 19257 21576
rect 19199 21567 19257 21573
rect 22462 21564 22468 21576
rect 22520 21564 22526 21616
rect 18187 21539 18245 21545
rect 18187 21505 18199 21539
rect 18233 21536 18245 21539
rect 21358 21536 21364 21548
rect 18233 21508 21364 21536
rect 18233 21505 18245 21508
rect 18187 21499 18245 21505
rect 21358 21496 21364 21508
rect 21416 21496 21422 21548
rect 9836 21471 9894 21477
rect 9836 21437 9848 21471
rect 9882 21437 9894 21471
rect 10870 21468 10876 21480
rect 10831 21440 10876 21468
rect 9836 21431 9894 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 10962 21428 10968 21480
rect 11020 21468 11026 21480
rect 11241 21471 11299 21477
rect 11241 21468 11253 21471
rect 11020 21440 11253 21468
rect 11020 21428 11026 21440
rect 11241 21437 11253 21440
rect 11287 21437 11299 21471
rect 12894 21468 12900 21480
rect 12855 21440 12900 21468
rect 11241 21431 11299 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 14642 21468 14648 21480
rect 14603 21440 14648 21468
rect 14642 21428 14648 21440
rect 14700 21428 14706 21480
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21468 15623 21471
rect 15930 21468 15936 21480
rect 15611 21440 15936 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 15930 21428 15936 21440
rect 15988 21468 15994 21480
rect 16301 21471 16359 21477
rect 16301 21468 16313 21471
rect 15988 21440 16313 21468
rect 15988 21428 15994 21440
rect 16301 21437 16313 21440
rect 16347 21468 16359 21471
rect 16485 21471 16543 21477
rect 16485 21468 16497 21471
rect 16347 21440 16497 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16485 21437 16497 21440
rect 16531 21437 16543 21471
rect 16485 21431 16543 21437
rect 18100 21471 18158 21477
rect 18100 21437 18112 21471
rect 18146 21437 18158 21471
rect 18100 21431 18158 21437
rect 7607 21372 8524 21400
rect 9309 21403 9367 21409
rect 7607 21369 7619 21372
rect 7561 21363 7619 21369
rect 9309 21369 9321 21403
rect 9355 21400 9367 21403
rect 10888 21400 10916 21428
rect 9355 21372 10916 21400
rect 11517 21403 11575 21409
rect 9355 21369 9367 21372
rect 9309 21363 9367 21369
rect 11517 21369 11529 21403
rect 11563 21400 11575 21403
rect 12158 21400 12164 21412
rect 11563 21372 12164 21400
rect 11563 21369 11575 21372
rect 11517 21363 11575 21369
rect 12158 21360 12164 21372
rect 12216 21360 12222 21412
rect 12802 21360 12808 21412
rect 12860 21400 12866 21412
rect 13218 21403 13276 21409
rect 13218 21400 13230 21403
rect 12860 21372 13230 21400
rect 12860 21360 12866 21372
rect 13218 21369 13230 21372
rect 13264 21400 13276 21403
rect 14461 21403 14519 21409
rect 14461 21400 14473 21403
rect 13264 21372 14473 21400
rect 13264 21369 13276 21372
rect 13218 21363 13276 21369
rect 14461 21369 14473 21372
rect 14507 21400 14519 21403
rect 14966 21403 15024 21409
rect 14966 21400 14978 21403
rect 14507 21372 14978 21400
rect 14507 21369 14519 21372
rect 14461 21363 14519 21369
rect 14966 21369 14978 21372
rect 15012 21400 15024 21403
rect 15286 21400 15292 21412
rect 15012 21372 15292 21400
rect 15012 21369 15024 21372
rect 14966 21363 15024 21369
rect 15286 21360 15292 21372
rect 15344 21360 15350 21412
rect 18115 21400 18143 21431
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 19096 21471 19154 21477
rect 19096 21468 19108 21471
rect 18840 21440 19108 21468
rect 18840 21428 18846 21440
rect 19096 21437 19108 21440
rect 19142 21468 19154 21471
rect 19889 21471 19947 21477
rect 19889 21468 19901 21471
rect 19142 21440 19901 21468
rect 19142 21437 19154 21440
rect 19096 21431 19154 21437
rect 19889 21437 19901 21440
rect 19935 21437 19947 21471
rect 19889 21431 19947 21437
rect 18322 21400 18328 21412
rect 18115 21372 18328 21400
rect 18322 21360 18328 21372
rect 18380 21400 18386 21412
rect 18877 21403 18935 21409
rect 18877 21400 18889 21403
rect 18380 21372 18889 21400
rect 18380 21360 18386 21372
rect 18877 21369 18889 21372
rect 18923 21369 18935 21403
rect 18877 21363 18935 21369
rect 2041 21335 2099 21341
rect 2041 21301 2053 21335
rect 2087 21332 2099 21335
rect 2332 21332 2360 21360
rect 2087 21304 2360 21332
rect 2087 21301 2099 21304
rect 2041 21295 2099 21301
rect 7926 21292 7932 21344
rect 7984 21332 7990 21344
rect 8297 21335 8355 21341
rect 8297 21332 8309 21335
rect 7984 21304 8309 21332
rect 7984 21292 7990 21304
rect 8297 21301 8309 21304
rect 8343 21301 8355 21335
rect 18506 21332 18512 21344
rect 18467 21304 18512 21332
rect 8297 21295 8355 21301
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 19518 21332 19524 21344
rect 19479 21304 19524 21332
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1762 21128 1768 21140
rect 1723 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 2314 21088 2320 21140
rect 2372 21128 2378 21140
rect 2501 21131 2559 21137
rect 2501 21128 2513 21131
rect 2372 21100 2513 21128
rect 2372 21088 2378 21100
rect 2501 21097 2513 21100
rect 2547 21097 2559 21131
rect 4246 21128 4252 21140
rect 4207 21100 4252 21128
rect 2501 21091 2559 21097
rect 4246 21088 4252 21100
rect 4304 21088 4310 21140
rect 5626 21128 5632 21140
rect 5587 21100 5632 21128
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 7926 21128 7932 21140
rect 7887 21100 7932 21128
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 9858 21088 9864 21140
rect 9916 21128 9922 21140
rect 10597 21131 10655 21137
rect 10597 21128 10609 21131
rect 9916 21100 10609 21128
rect 9916 21088 9922 21100
rect 10597 21097 10609 21100
rect 10643 21097 10655 21131
rect 10597 21091 10655 21097
rect 10870 21088 10876 21140
rect 10928 21128 10934 21140
rect 10965 21131 11023 21137
rect 10965 21128 10977 21131
rect 10928 21100 10977 21128
rect 10928 21088 10934 21100
rect 10965 21097 10977 21100
rect 11011 21128 11023 21131
rect 11011 21100 12388 21128
rect 11011 21097 11023 21100
rect 10965 21091 11023 21097
rect 3694 21020 3700 21072
rect 3752 21060 3758 21072
rect 5074 21060 5080 21072
rect 3752 21032 5080 21060
rect 3752 21020 3758 21032
rect 5074 21020 5080 21032
rect 5132 21020 5138 21072
rect 6270 21060 6276 21072
rect 5828 21032 6276 21060
rect 2869 20995 2927 21001
rect 2869 20961 2881 20995
rect 2915 20992 2927 20995
rect 3234 20992 3240 21004
rect 2915 20964 3240 20992
rect 2915 20961 2927 20964
rect 2869 20955 2927 20961
rect 3234 20952 3240 20964
rect 3292 20952 3298 21004
rect 4065 20995 4123 21001
rect 4065 20961 4077 20995
rect 4111 20961 4123 20995
rect 4065 20955 4123 20961
rect 3786 20884 3792 20936
rect 3844 20924 3850 20936
rect 4080 20924 4108 20955
rect 5166 20952 5172 21004
rect 5224 20992 5230 21004
rect 5828 21001 5856 21032
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 8757 21063 8815 21069
rect 8757 21029 8769 21063
rect 8803 21060 8815 21063
rect 9030 21060 9036 21072
rect 8803 21032 9036 21060
rect 8803 21029 8815 21032
rect 8757 21023 8815 21029
rect 9030 21020 9036 21032
rect 9088 21020 9094 21072
rect 10039 21063 10097 21069
rect 10039 21029 10051 21063
rect 10085 21060 10097 21063
rect 10686 21060 10692 21072
rect 10085 21032 10692 21060
rect 10085 21029 10097 21032
rect 10039 21023 10097 21029
rect 10686 21020 10692 21032
rect 10744 21020 10750 21072
rect 12250 21060 12256 21072
rect 12211 21032 12256 21060
rect 12250 21020 12256 21032
rect 12308 21020 12314 21072
rect 12360 21060 12388 21100
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 13173 21131 13231 21137
rect 13173 21128 13185 21131
rect 12952 21100 13185 21128
rect 12952 21088 12958 21100
rect 13173 21097 13185 21100
rect 13219 21097 13231 21131
rect 13173 21091 13231 21097
rect 17310 21060 17316 21072
rect 12360 21032 13400 21060
rect 17271 21032 17316 21060
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5224 20964 5825 20992
rect 5224 20952 5230 20964
rect 5813 20961 5825 20964
rect 5859 20961 5871 20995
rect 6086 20992 6092 21004
rect 6047 20964 6092 20992
rect 5813 20955 5871 20961
rect 6086 20952 6092 20964
rect 6144 20952 6150 21004
rect 6362 20992 6368 21004
rect 6323 20964 6368 20992
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 8294 20992 8300 21004
rect 8255 20964 8300 20992
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 8478 20992 8484 21004
rect 8439 20964 8484 20992
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 11790 20992 11796 21004
rect 11751 20964 11796 20992
rect 11790 20952 11796 20964
rect 11848 20952 11854 21004
rect 11977 20995 12035 21001
rect 11977 20961 11989 20995
rect 12023 20961 12035 20995
rect 11977 20955 12035 20961
rect 3844 20896 4108 20924
rect 5445 20927 5503 20933
rect 3844 20884 3850 20896
rect 5445 20893 5457 20927
rect 5491 20924 5503 20927
rect 6104 20924 6132 20952
rect 9674 20924 9680 20936
rect 5491 20896 6132 20924
rect 9635 20896 9680 20924
rect 5491 20893 5503 20896
rect 5445 20887 5503 20893
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 11992 20924 12020 20955
rect 12158 20952 12164 21004
rect 12216 20992 12222 21004
rect 13372 21001 13400 21032
rect 17310 21020 17316 21032
rect 17368 21020 17374 21072
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12216 20964 12909 20992
rect 12216 20952 12222 20964
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 13357 20995 13415 21001
rect 13357 20961 13369 20995
rect 13403 20992 13415 20995
rect 13446 20992 13452 21004
rect 13403 20964 13452 20992
rect 13403 20961 13415 20964
rect 13357 20955 13415 20961
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 13541 20995 13599 21001
rect 13541 20961 13553 20995
rect 13587 20961 13599 20995
rect 15470 20992 15476 21004
rect 15431 20964 15476 20992
rect 13541 20955 13599 20961
rect 13556 20924 13584 20955
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 19058 20992 19064 21004
rect 19019 20964 19064 20992
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 11256 20896 12020 20924
rect 12912 20896 13584 20924
rect 4893 20791 4951 20797
rect 4893 20757 4905 20791
rect 4939 20788 4951 20791
rect 5442 20788 5448 20800
rect 4939 20760 5448 20788
rect 4939 20757 4951 20760
rect 4893 20751 4951 20757
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 6914 20788 6920 20800
rect 6875 20760 6920 20788
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 9490 20788 9496 20800
rect 9451 20760 9496 20788
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11256 20797 11284 20896
rect 12912 20800 12940 20896
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14516 20896 15301 20924
rect 14516 20884 14522 20896
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 17218 20924 17224 20936
rect 17179 20896 17224 20924
rect 15289 20887 15347 20893
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 18230 20884 18236 20936
rect 18288 20924 18294 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18288 20896 18705 20924
rect 18288 20884 18294 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 17773 20859 17831 20865
rect 17773 20825 17785 20859
rect 17819 20856 17831 20859
rect 18782 20856 18788 20868
rect 17819 20828 18788 20856
rect 17819 20825 17831 20828
rect 17773 20819 17831 20825
rect 18782 20816 18788 20828
rect 18840 20816 18846 20868
rect 11241 20791 11299 20797
rect 11241 20788 11253 20791
rect 11020 20760 11253 20788
rect 11020 20748 11026 20760
rect 11241 20757 11253 20760
rect 11287 20757 11299 20791
rect 11241 20751 11299 20757
rect 12621 20791 12679 20797
rect 12621 20757 12633 20791
rect 12667 20788 12679 20791
rect 12894 20788 12900 20800
rect 12667 20760 12900 20788
rect 12667 20757 12679 20760
rect 12621 20751 12679 20757
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13170 20748 13176 20800
rect 13228 20788 13234 20800
rect 14642 20788 14648 20800
rect 13228 20760 14648 20788
rect 13228 20748 13234 20760
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 16482 20788 16488 20800
rect 16443 20760 16488 20788
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 18138 20788 18144 20800
rect 18099 20760 18144 20788
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 3878 20584 3884 20596
rect 3839 20556 3884 20584
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 5905 20587 5963 20593
rect 5905 20553 5917 20587
rect 5951 20584 5963 20587
rect 5994 20584 6000 20596
rect 5951 20556 6000 20584
rect 5951 20553 5963 20556
rect 5905 20547 5963 20553
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 6270 20584 6276 20596
rect 6183 20556 6276 20584
rect 6270 20544 6276 20556
rect 6328 20584 6334 20596
rect 9398 20584 9404 20596
rect 6328 20556 9404 20584
rect 6328 20544 6334 20556
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 10413 20587 10471 20593
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 10686 20584 10692 20596
rect 10459 20556 10692 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 14369 20587 14427 20593
rect 14369 20553 14381 20587
rect 14415 20584 14427 20587
rect 14642 20584 14648 20596
rect 14415 20556 14648 20584
rect 14415 20553 14427 20556
rect 14369 20547 14427 20553
rect 14642 20544 14648 20556
rect 14700 20584 14706 20596
rect 15470 20584 15476 20596
rect 14700 20556 15476 20584
rect 14700 20544 14706 20556
rect 15470 20544 15476 20556
rect 15528 20544 15534 20596
rect 16482 20584 16488 20596
rect 16395 20556 16488 20584
rect 3142 20516 3148 20528
rect 2240 20488 3148 20516
rect 2240 20457 2268 20488
rect 3142 20476 3148 20488
rect 3200 20476 3206 20528
rect 7745 20519 7803 20525
rect 7745 20516 7757 20519
rect 5920 20488 7757 20516
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20417 2283 20451
rect 2866 20448 2872 20460
rect 2827 20420 2872 20448
rect 2225 20411 2283 20417
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 3234 20448 3240 20460
rect 3007 20420 3240 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 3234 20408 3240 20420
rect 3292 20448 3298 20460
rect 5920 20448 5948 20488
rect 7745 20485 7757 20488
rect 7791 20485 7803 20519
rect 7745 20479 7803 20485
rect 9309 20519 9367 20525
rect 9309 20485 9321 20519
rect 9355 20516 9367 20519
rect 11790 20516 11796 20528
rect 9355 20488 11796 20516
rect 9355 20485 9367 20488
rect 9309 20479 9367 20485
rect 3292 20420 5948 20448
rect 3292 20408 3298 20420
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6512 20420 6561 20448
rect 6512 20408 6518 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 3697 20383 3755 20389
rect 3697 20380 3709 20383
rect 3528 20352 3709 20380
rect 1673 20315 1731 20321
rect 1673 20281 1685 20315
rect 1719 20312 1731 20315
rect 2041 20315 2099 20321
rect 2041 20312 2053 20315
rect 1719 20284 2053 20312
rect 1719 20281 1731 20284
rect 1673 20275 1731 20281
rect 2041 20281 2053 20284
rect 2087 20312 2099 20315
rect 2317 20315 2375 20321
rect 2317 20312 2329 20315
rect 2087 20284 2329 20312
rect 2087 20281 2099 20284
rect 2041 20275 2099 20281
rect 2317 20281 2329 20284
rect 2363 20281 2375 20315
rect 2317 20275 2375 20281
rect 2332 20244 2360 20275
rect 2866 20272 2872 20324
rect 2924 20312 2930 20324
rect 3528 20321 3556 20352
rect 3697 20349 3709 20352
rect 3743 20349 3755 20383
rect 3697 20343 3755 20349
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 5077 20383 5135 20389
rect 5077 20380 5089 20383
rect 4755 20352 5089 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 5077 20349 5089 20352
rect 5123 20380 5135 20383
rect 5166 20380 5172 20392
rect 5123 20352 5172 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5500 20352 5641 20380
rect 5500 20340 5506 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 5813 20383 5871 20389
rect 5813 20349 5825 20383
rect 5859 20380 5871 20383
rect 5902 20380 5908 20392
rect 5859 20352 5908 20380
rect 5859 20349 5871 20352
rect 5813 20343 5871 20349
rect 3513 20315 3571 20321
rect 3513 20312 3525 20315
rect 2924 20284 3525 20312
rect 2924 20272 2930 20284
rect 3513 20281 3525 20284
rect 3559 20281 3571 20315
rect 3513 20275 3571 20281
rect 4341 20315 4399 20321
rect 4341 20281 4353 20315
rect 4387 20312 4399 20315
rect 5828 20312 5856 20343
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6564 20312 6592 20411
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 6914 20380 6920 20392
rect 6871 20352 6920 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 8294 20380 8300 20392
rect 8159 20352 8300 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 8294 20340 8300 20352
rect 8352 20380 8358 20392
rect 9416 20389 9444 20488
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 10134 20448 10140 20460
rect 10095 20420 10140 20448
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 11330 20448 11336 20460
rect 11291 20420 11336 20448
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 13170 20448 13176 20460
rect 13131 20420 13176 20448
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 14550 20448 14556 20460
rect 14511 20420 14556 20448
rect 14550 20408 14556 20420
rect 14608 20408 14614 20460
rect 14826 20448 14832 20460
rect 14787 20420 14832 20448
rect 14826 20408 14832 20420
rect 14884 20408 14890 20460
rect 16408 20448 16436 20556
rect 16482 20544 16488 20556
rect 16540 20584 16546 20596
rect 16540 20556 16620 20584
rect 16540 20544 16546 20556
rect 16592 20516 16620 20556
rect 17310 20544 17316 20596
rect 17368 20584 17374 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17368 20556 17509 20584
rect 17368 20544 17374 20556
rect 17497 20553 17509 20556
rect 17543 20584 17555 20587
rect 19058 20584 19064 20596
rect 17543 20556 19064 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 16592 20488 19748 20516
rect 16474 20451 16532 20457
rect 16474 20448 16486 20451
rect 16408 20420 16486 20448
rect 16474 20417 16486 20420
rect 16520 20417 16532 20451
rect 18138 20448 18144 20460
rect 18051 20420 18144 20448
rect 16474 20411 16532 20417
rect 18138 20408 18144 20420
rect 18196 20448 18202 20460
rect 19613 20451 19671 20457
rect 19613 20448 19625 20451
rect 18196 20420 19625 20448
rect 18196 20408 18202 20420
rect 19613 20417 19625 20420
rect 19659 20417 19671 20451
rect 19720 20448 19748 20488
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 19720 20420 20637 20448
rect 19613 20411 19671 20417
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 8352 20352 9413 20380
rect 8352 20340 8358 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 9858 20380 9864 20392
rect 9548 20352 9864 20380
rect 9548 20340 9554 20352
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12176 20352 12449 20380
rect 6638 20312 6644 20324
rect 4387 20284 5856 20312
rect 6551 20284 6644 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 6638 20272 6644 20284
rect 6696 20312 6702 20324
rect 7146 20315 7204 20321
rect 7146 20312 7158 20315
rect 6696 20284 7158 20312
rect 6696 20272 6702 20284
rect 7146 20281 7158 20284
rect 7192 20281 7204 20315
rect 7146 20275 7204 20281
rect 8941 20315 8999 20321
rect 8941 20281 8953 20315
rect 8987 20312 8999 20315
rect 9674 20312 9680 20324
rect 8987 20284 9680 20312
rect 8987 20281 8999 20284
rect 8941 20275 8999 20281
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 2961 20247 3019 20253
rect 2961 20244 2973 20247
rect 2332 20216 2973 20244
rect 2961 20213 2973 20216
rect 3007 20213 3019 20247
rect 3142 20244 3148 20256
rect 3103 20216 3148 20244
rect 2961 20207 3019 20213
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 8478 20244 8484 20256
rect 8439 20216 8484 20244
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 10962 20204 10968 20256
rect 11020 20244 11026 20256
rect 11149 20247 11207 20253
rect 11149 20244 11161 20247
rect 11020 20216 11161 20244
rect 11020 20204 11026 20216
rect 11149 20213 11161 20216
rect 11195 20213 11207 20247
rect 11790 20244 11796 20256
rect 11751 20216 11796 20244
rect 11149 20207 11207 20213
rect 11790 20204 11796 20216
rect 11848 20244 11854 20256
rect 12176 20253 12204 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 12894 20380 12900 20392
rect 12855 20352 12900 20380
rect 12437 20343 12495 20349
rect 12894 20340 12900 20352
rect 12952 20380 12958 20392
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 12952 20352 13829 20380
rect 12952 20340 12958 20352
rect 13817 20349 13829 20352
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 14642 20312 14648 20324
rect 14603 20284 14648 20312
rect 14642 20272 14648 20284
rect 14700 20272 14706 20324
rect 16301 20315 16359 20321
rect 16301 20281 16313 20315
rect 16347 20312 16359 20315
rect 16577 20315 16635 20321
rect 16577 20312 16589 20315
rect 16347 20284 16589 20312
rect 16347 20281 16359 20284
rect 16301 20275 16359 20281
rect 16577 20281 16589 20284
rect 16623 20312 16635 20315
rect 16850 20312 16856 20324
rect 16623 20284 16856 20312
rect 16623 20281 16635 20284
rect 16577 20275 16635 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 17129 20315 17187 20321
rect 17129 20281 17141 20315
rect 17175 20312 17187 20315
rect 18138 20312 18144 20324
rect 17175 20284 18144 20312
rect 17175 20281 17187 20284
rect 17129 20275 17187 20281
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 18230 20272 18236 20324
rect 18288 20312 18294 20324
rect 18782 20312 18788 20324
rect 18288 20284 18333 20312
rect 18743 20284 18788 20312
rect 18288 20272 18294 20284
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 11848 20216 12173 20244
rect 11848 20204 11854 20216
rect 12161 20213 12173 20216
rect 12207 20213 12219 20247
rect 13538 20244 13544 20256
rect 13499 20216 13544 20244
rect 12161 20207 12219 20213
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 17865 20247 17923 20253
rect 17865 20213 17877 20247
rect 17911 20244 17923 20247
rect 18248 20244 18276 20272
rect 17911 20216 18276 20244
rect 17911 20213 17923 20216
rect 17865 20207 17923 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2222 20000 2228 20052
rect 2280 20040 2286 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2280 20012 2973 20040
rect 2280 20000 2286 20012
rect 2961 20009 2973 20012
rect 3007 20009 3019 20043
rect 2961 20003 3019 20009
rect 5905 20043 5963 20049
rect 5905 20009 5917 20043
rect 5951 20040 5963 20043
rect 5994 20040 6000 20052
rect 5951 20012 6000 20040
rect 5951 20009 5963 20012
rect 5905 20003 5963 20009
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 9769 20043 9827 20049
rect 9769 20040 9781 20043
rect 9732 20012 9781 20040
rect 9732 20000 9738 20012
rect 9769 20009 9781 20012
rect 9815 20009 9827 20043
rect 9769 20003 9827 20009
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14608 20012 14657 20040
rect 14608 20000 14614 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 17310 20040 17316 20052
rect 16991 20012 17316 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 17310 20000 17316 20012
rect 17368 20000 17374 20052
rect 24581 20043 24639 20049
rect 24581 20009 24593 20043
rect 24627 20040 24639 20043
rect 26326 20040 26332 20052
rect 24627 20012 26332 20040
rect 24627 20009 24639 20012
rect 24581 20003 24639 20009
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 1670 19932 1676 19984
rect 1728 19972 1734 19984
rect 2501 19975 2559 19981
rect 2501 19972 2513 19975
rect 1728 19944 2513 19972
rect 1728 19932 1734 19944
rect 2501 19941 2513 19944
rect 2547 19972 2559 19975
rect 3050 19972 3056 19984
rect 2547 19944 3056 19972
rect 2547 19941 2559 19944
rect 2501 19935 2559 19941
rect 3050 19932 3056 19944
rect 3108 19932 3114 19984
rect 4249 19975 4307 19981
rect 4249 19941 4261 19975
rect 4295 19972 4307 19975
rect 4338 19972 4344 19984
rect 4295 19944 4344 19972
rect 4295 19941 4307 19944
rect 4249 19935 4307 19941
rect 4338 19932 4344 19944
rect 4396 19932 4402 19984
rect 4798 19972 4804 19984
rect 4759 19944 4804 19972
rect 4798 19932 4804 19944
rect 4856 19932 4862 19984
rect 5074 19932 5080 19984
rect 5132 19972 5138 19984
rect 5629 19975 5687 19981
rect 5629 19972 5641 19975
rect 5132 19944 5641 19972
rect 5132 19932 5138 19944
rect 5629 19941 5641 19944
rect 5675 19972 5687 19975
rect 6362 19972 6368 19984
rect 5675 19944 6368 19972
rect 5675 19941 5687 19944
rect 5629 19935 5687 19941
rect 6362 19932 6368 19944
rect 6420 19972 6426 19984
rect 7929 19975 7987 19981
rect 6420 19944 6684 19972
rect 6420 19932 6426 19944
rect 2038 19904 2044 19916
rect 1999 19876 2044 19904
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 6086 19904 6092 19916
rect 6047 19876 6092 19904
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 6656 19913 6684 19944
rect 7929 19941 7941 19975
rect 7975 19972 7987 19975
rect 10870 19972 10876 19984
rect 7975 19944 8616 19972
rect 7975 19941 7987 19944
rect 7929 19935 7987 19941
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 7098 19904 7104 19916
rect 6687 19876 7104 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 8294 19904 8300 19916
rect 8255 19876 8300 19904
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8588 19913 8616 19944
rect 9784 19944 10876 19972
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19904 8631 19907
rect 8754 19904 8760 19916
rect 8619 19876 8760 19904
rect 8619 19873 8631 19876
rect 8573 19867 8631 19873
rect 8754 19864 8760 19876
rect 8812 19864 8818 19916
rect 9784 19913 9812 19944
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 13817 19975 13875 19981
rect 13817 19941 13829 19975
rect 13863 19972 13875 19975
rect 14182 19972 14188 19984
rect 13863 19944 14188 19972
rect 13863 19941 13875 19944
rect 13817 19935 13875 19941
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 15286 19932 15292 19984
rect 15344 19972 15350 19984
rect 16346 19975 16404 19981
rect 16346 19972 16358 19975
rect 15344 19944 16358 19972
rect 15344 19932 15350 19944
rect 16346 19941 16358 19944
rect 16392 19941 16404 19975
rect 17954 19972 17960 19984
rect 17915 19944 17960 19972
rect 16346 19935 16404 19941
rect 17954 19932 17960 19944
rect 18012 19972 18018 19984
rect 18785 19975 18843 19981
rect 18785 19972 18797 19975
rect 18012 19944 18797 19972
rect 18012 19932 18018 19944
rect 18785 19941 18797 19944
rect 18831 19941 18843 19975
rect 18785 19935 18843 19941
rect 9769 19907 9827 19913
rect 9769 19873 9781 19907
rect 9815 19873 9827 19907
rect 9769 19867 9827 19873
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9916 19876 10149 19904
rect 9916 19864 9922 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 11790 19904 11796 19916
rect 11751 19876 11796 19904
rect 10137 19867 10195 19873
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 12158 19904 12164 19916
rect 12119 19876 12164 19904
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 19334 19904 19340 19916
rect 19295 19876 19340 19904
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 24210 19864 24216 19916
rect 24268 19904 24274 19916
rect 24397 19907 24455 19913
rect 24397 19904 24409 19907
rect 24268 19876 24409 19904
rect 24268 19864 24274 19876
rect 24397 19873 24409 19876
rect 24443 19873 24455 19907
rect 24397 19867 24455 19873
rect 2130 19836 2136 19848
rect 2091 19808 2136 19836
rect 2130 19796 2136 19808
rect 2188 19796 2194 19848
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4522 19836 4528 19848
rect 4203 19808 4528 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 5902 19796 5908 19848
rect 5960 19836 5966 19848
rect 6733 19839 6791 19845
rect 6733 19836 6745 19839
rect 5960 19808 6745 19836
rect 5960 19796 5966 19808
rect 6733 19805 6745 19808
rect 6779 19836 6791 19839
rect 8662 19836 8668 19848
rect 6779 19808 7328 19836
rect 8623 19808 8668 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 3234 19728 3240 19780
rect 3292 19768 3298 19780
rect 3786 19768 3792 19780
rect 3292 19740 3792 19768
rect 3292 19728 3298 19740
rect 3786 19728 3792 19740
rect 3844 19728 3850 19780
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 5166 19700 5172 19712
rect 5127 19672 5172 19700
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 7300 19709 7328 19808
rect 8662 19796 8668 19808
rect 8720 19796 8726 19848
rect 12437 19839 12495 19845
rect 12437 19805 12449 19839
rect 12483 19836 12495 19839
rect 13078 19836 13084 19848
rect 12483 19808 13084 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 13587 19808 13737 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13725 19805 13737 19808
rect 13771 19836 13783 19839
rect 13814 19836 13820 19848
rect 13771 19808 13820 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13814 19796 13820 19808
rect 13872 19796 13878 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 15654 19836 15660 19848
rect 14415 19808 15660 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16022 19836 16028 19848
rect 15983 19808 16028 19836
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19805 17923 19839
rect 18322 19836 18328 19848
rect 18283 19808 18328 19836
rect 17865 19799 17923 19805
rect 15672 19768 15700 19796
rect 17589 19771 17647 19777
rect 17589 19768 17601 19771
rect 15672 19740 17601 19768
rect 17589 19737 17601 19740
rect 17635 19768 17647 19771
rect 17880 19768 17908 19799
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 17635 19740 17908 19768
rect 17635 19737 17647 19740
rect 17589 19731 17647 19737
rect 7285 19703 7343 19709
rect 7285 19669 7297 19703
rect 7331 19700 7343 19703
rect 7926 19700 7932 19712
rect 7331 19672 7932 19700
rect 7331 19669 7343 19672
rect 7285 19663 7343 19669
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 9398 19700 9404 19712
rect 9359 19672 9404 19700
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 12986 19700 12992 19712
rect 12947 19672 12992 19700
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 14826 19660 14832 19712
rect 14884 19700 14890 19712
rect 17218 19700 17224 19712
rect 14884 19672 17224 19700
rect 14884 19660 14890 19672
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 19518 19700 19524 19712
rect 19479 19672 19524 19700
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 4157 19499 4215 19505
rect 4157 19465 4169 19499
rect 4203 19496 4215 19499
rect 4338 19496 4344 19508
rect 4203 19468 4344 19496
rect 4203 19465 4215 19468
rect 4157 19459 4215 19465
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 8294 19496 8300 19508
rect 8255 19468 8300 19496
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 9398 19456 9404 19508
rect 9456 19505 9462 19508
rect 9456 19499 9505 19505
rect 9456 19465 9459 19499
rect 9493 19465 9505 19499
rect 9456 19459 9505 19465
rect 9456 19456 9462 19459
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9916 19468 9965 19496
rect 9916 19456 9922 19468
rect 9953 19465 9965 19468
rect 9999 19496 10011 19499
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 9999 19468 10701 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 10689 19465 10701 19468
rect 10735 19465 10747 19499
rect 12158 19496 12164 19508
rect 12119 19468 12164 19496
rect 10689 19459 10747 19465
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 12802 19496 12808 19508
rect 12763 19468 12808 19496
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19496 13967 19499
rect 14642 19496 14648 19508
rect 13955 19468 14648 19496
rect 13955 19465 13967 19468
rect 13909 19459 13967 19465
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 14921 19499 14979 19505
rect 14921 19465 14933 19499
rect 14967 19496 14979 19499
rect 15105 19499 15163 19505
rect 15105 19496 15117 19499
rect 14967 19468 15117 19496
rect 14967 19465 14979 19468
rect 14921 19459 14979 19465
rect 15105 19465 15117 19468
rect 15151 19496 15163 19499
rect 15286 19496 15292 19508
rect 15151 19468 15292 19496
rect 15151 19465 15163 19468
rect 15105 19459 15163 19465
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 16117 19499 16175 19505
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 16163 19468 17693 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 17681 19465 17693 19468
rect 17727 19496 17739 19499
rect 17773 19499 17831 19505
rect 17773 19496 17785 19499
rect 17727 19468 17785 19496
rect 17727 19465 17739 19468
rect 17681 19459 17739 19465
rect 17773 19465 17785 19468
rect 17819 19496 17831 19499
rect 17954 19496 17960 19508
rect 17819 19468 17960 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 19334 19496 19340 19508
rect 19295 19468 19340 19496
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 2593 19431 2651 19437
rect 2593 19428 2605 19431
rect 2096 19400 2605 19428
rect 2096 19388 2102 19400
rect 2593 19397 2605 19400
rect 2639 19428 2651 19431
rect 3510 19428 3516 19440
rect 2639 19400 3516 19428
rect 2639 19397 2651 19400
rect 2593 19391 2651 19397
rect 3510 19388 3516 19400
rect 3568 19388 3574 19440
rect 3697 19431 3755 19437
rect 3697 19397 3709 19431
rect 3743 19428 3755 19431
rect 4798 19428 4804 19440
rect 3743 19400 4804 19428
rect 3743 19397 3755 19400
rect 3697 19391 3755 19397
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 9582 19428 9588 19440
rect 9543 19400 9588 19428
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 10413 19431 10471 19437
rect 10413 19397 10425 19431
rect 10459 19428 10471 19431
rect 10870 19428 10876 19440
rect 10459 19400 10876 19428
rect 10459 19397 10471 19400
rect 10413 19391 10471 19397
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 11790 19428 11796 19440
rect 11703 19400 11796 19428
rect 11790 19388 11796 19400
rect 11848 19428 11854 19440
rect 19518 19428 19524 19440
rect 11848 19400 19524 19428
rect 11848 19388 11854 19400
rect 19518 19388 19524 19400
rect 19576 19388 19582 19440
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 1670 19360 1676 19372
rect 1627 19332 1676 19360
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19360 3203 19363
rect 3418 19360 3424 19372
rect 3191 19332 3424 19360
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 4522 19360 4528 19372
rect 4435 19332 4528 19360
rect 4522 19320 4528 19332
rect 4580 19360 4586 19372
rect 9677 19363 9735 19369
rect 4580 19332 8064 19360
rect 4580 19320 4586 19332
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19292 5043 19295
rect 5074 19292 5080 19304
rect 5031 19264 5080 19292
rect 5031 19261 5043 19264
rect 4985 19255 5043 19261
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5166 19252 5172 19304
rect 5224 19292 5230 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5224 19264 5641 19292
rect 5224 19252 5230 19264
rect 5629 19261 5641 19264
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 1673 19227 1731 19233
rect 1673 19193 1685 19227
rect 1719 19224 1731 19227
rect 2038 19224 2044 19236
rect 1719 19196 2044 19224
rect 1719 19193 1731 19196
rect 1673 19187 1731 19193
rect 2038 19184 2044 19196
rect 2096 19184 2102 19236
rect 2222 19224 2228 19236
rect 2183 19196 2228 19224
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 3237 19227 3295 19233
rect 3237 19193 3249 19227
rect 3283 19193 3295 19227
rect 5644 19224 5672 19255
rect 6086 19252 6092 19304
rect 6144 19292 6150 19304
rect 6181 19295 6239 19301
rect 6181 19292 6193 19295
rect 6144 19264 6193 19292
rect 6144 19252 6150 19264
rect 6181 19261 6193 19264
rect 6227 19292 6239 19295
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 6227 19264 6653 19292
rect 6227 19261 6239 19264
rect 6181 19255 6239 19261
rect 6641 19261 6653 19264
rect 6687 19292 6699 19295
rect 7101 19295 7159 19301
rect 7101 19292 7113 19295
rect 6687 19264 7113 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7101 19261 7113 19264
rect 7147 19261 7159 19295
rect 7650 19292 7656 19304
rect 7611 19264 7656 19292
rect 7101 19255 7159 19261
rect 7116 19224 7144 19255
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 7837 19295 7895 19301
rect 7837 19261 7849 19295
rect 7883 19292 7895 19295
rect 7926 19292 7932 19304
rect 7883 19264 7932 19292
rect 7883 19261 7895 19264
rect 7837 19255 7895 19261
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8036 19292 8064 19332
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9858 19360 9864 19372
rect 9723 19332 9864 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 12986 19360 12992 19372
rect 12947 19332 12992 19360
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 16022 19320 16028 19372
rect 16080 19360 16086 19372
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16080 19332 16773 19360
rect 16080 19320 16086 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 16908 19332 18061 19360
rect 16908 19320 16914 19332
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 19751 19363 19809 19369
rect 19751 19329 19763 19363
rect 19797 19360 19809 19363
rect 24210 19360 24216 19372
rect 19797 19332 24216 19360
rect 19797 19329 19809 19332
rect 19751 19323 19809 19329
rect 24210 19320 24216 19332
rect 24268 19360 24274 19372
rect 24397 19363 24455 19369
rect 24397 19360 24409 19363
rect 24268 19332 24409 19360
rect 24268 19320 24274 19332
rect 24397 19329 24409 19332
rect 24443 19329 24455 19363
rect 24397 19323 24455 19329
rect 10873 19295 10931 19301
rect 10873 19292 10885 19295
rect 8036 19264 10885 19292
rect 10873 19261 10885 19264
rect 10919 19261 10931 19295
rect 10873 19255 10931 19261
rect 13078 19252 13084 19304
rect 13136 19292 13142 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 13136 19264 14657 19292
rect 13136 19252 13142 19264
rect 14645 19261 14657 19264
rect 14691 19292 14703 19295
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 14691 19264 15209 19292
rect 14691 19261 14703 19264
rect 14645 19255 14703 19261
rect 15197 19261 15209 19264
rect 15243 19261 15255 19295
rect 16942 19292 16948 19304
rect 16903 19264 16948 19292
rect 15197 19255 15255 19261
rect 16942 19252 16948 19264
rect 17000 19292 17006 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 17000 19264 17417 19292
rect 17000 19252 17006 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 17681 19295 17739 19301
rect 17681 19261 17693 19295
rect 17727 19292 17739 19295
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 17727 19264 18153 19292
rect 17727 19261 17739 19264
rect 17681 19255 17739 19261
rect 18141 19261 18153 19264
rect 18187 19261 18199 19295
rect 18141 19255 18199 19261
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 19664 19295 19722 19301
rect 19664 19292 19676 19295
rect 18748 19264 19676 19292
rect 18748 19252 18754 19264
rect 19664 19261 19676 19264
rect 19710 19292 19722 19295
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 19710 19264 20085 19292
rect 19710 19261 19722 19264
rect 19664 19255 19722 19261
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 8018 19224 8024 19236
rect 5644 19196 7052 19224
rect 7116 19196 8024 19224
rect 3237 19187 3295 19193
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 3252 19156 3280 19187
rect 4798 19156 4804 19168
rect 3007 19128 4804 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5166 19156 5172 19168
rect 5127 19128 5172 19156
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 6914 19156 6920 19168
rect 6875 19128 6920 19156
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7024 19156 7052 19196
rect 8018 19184 8024 19196
rect 8076 19224 8082 19236
rect 8849 19227 8907 19233
rect 8849 19224 8861 19227
rect 8076 19196 8861 19224
rect 8076 19184 8082 19196
rect 8849 19193 8861 19196
rect 8895 19224 8907 19227
rect 9306 19224 9312 19236
rect 8895 19196 9312 19224
rect 8895 19193 8907 19196
rect 8849 19187 8907 19193
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19224 14979 19227
rect 15559 19227 15617 19233
rect 15559 19224 15571 19227
rect 14967 19196 15571 19224
rect 14967 19193 14979 19196
rect 14921 19187 14979 19193
rect 15559 19193 15571 19196
rect 15605 19224 15617 19227
rect 16390 19224 16396 19236
rect 15605 19196 16396 19224
rect 15605 19193 15617 19196
rect 15559 19187 15617 19193
rect 16390 19184 16396 19196
rect 16448 19184 16454 19236
rect 19058 19224 19064 19236
rect 16500 19196 19064 19224
rect 7282 19156 7288 19168
rect 7024 19128 7288 19156
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19156 9275 19159
rect 9858 19156 9864 19168
rect 9263 19128 9864 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9858 19116 9864 19128
rect 9916 19156 9922 19168
rect 10134 19156 10140 19168
rect 9916 19128 10140 19156
rect 9916 19116 9922 19128
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 13354 19156 13360 19168
rect 13315 19128 13360 19156
rect 13354 19116 13360 19128
rect 13412 19116 13418 19168
rect 14274 19156 14280 19168
rect 14187 19128 14280 19156
rect 14274 19116 14280 19128
rect 14332 19156 14338 19168
rect 16500 19156 16528 19196
rect 19058 19184 19064 19196
rect 19116 19184 19122 19236
rect 14332 19128 16528 19156
rect 14332 19116 14338 19128
rect 16850 19116 16856 19168
rect 16908 19156 16914 19168
rect 17129 19159 17187 19165
rect 17129 19156 17141 19159
rect 16908 19128 17141 19156
rect 16908 19116 16914 19128
rect 17129 19125 17141 19128
rect 17175 19125 17187 19159
rect 17129 19119 17187 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2038 18952 2044 18964
rect 1999 18924 2044 18952
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 5074 18952 5080 18964
rect 2188 18924 4154 18952
rect 5035 18924 5080 18952
rect 2188 18912 2194 18924
rect 2406 18844 2412 18896
rect 2464 18884 2470 18896
rect 2501 18887 2559 18893
rect 2501 18884 2513 18887
rect 2464 18856 2513 18884
rect 2464 18844 2470 18856
rect 2501 18853 2513 18856
rect 2547 18853 2559 18887
rect 2501 18847 2559 18853
rect 3053 18887 3111 18893
rect 3053 18853 3065 18887
rect 3099 18884 3111 18887
rect 3418 18884 3424 18896
rect 3099 18856 3424 18884
rect 3099 18853 3111 18856
rect 3053 18847 3111 18853
rect 3418 18844 3424 18856
rect 3476 18844 3482 18896
rect 4126 18884 4154 18924
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 10321 18955 10379 18961
rect 10321 18952 10333 18955
rect 8536 18924 10333 18952
rect 8536 18912 8542 18924
rect 10321 18921 10333 18924
rect 10367 18921 10379 18955
rect 10321 18915 10379 18921
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 16945 18955 17003 18961
rect 16945 18952 16957 18955
rect 13044 18924 16957 18952
rect 13044 18912 13050 18924
rect 16945 18921 16957 18924
rect 16991 18921 17003 18955
rect 16945 18915 17003 18921
rect 4246 18884 4252 18896
rect 4126 18856 4252 18884
rect 4246 18844 4252 18856
rect 4304 18844 4310 18896
rect 6178 18893 6184 18896
rect 6175 18884 6184 18893
rect 6091 18856 6184 18884
rect 6175 18847 6184 18856
rect 6236 18884 6242 18896
rect 6638 18884 6644 18896
rect 6236 18856 6644 18884
rect 6178 18844 6184 18847
rect 6236 18844 6242 18856
rect 6638 18844 6644 18856
rect 6696 18844 6702 18896
rect 7929 18887 7987 18893
rect 7929 18853 7941 18887
rect 7975 18884 7987 18887
rect 8018 18884 8024 18896
rect 7975 18856 8024 18884
rect 7975 18853 7987 18856
rect 7929 18847 7987 18853
rect 8018 18844 8024 18856
rect 8076 18844 8082 18896
rect 9398 18884 9404 18896
rect 8214 18856 9404 18884
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18816 5871 18819
rect 5994 18816 6000 18828
rect 5859 18788 6000 18816
rect 5859 18785 5871 18788
rect 5813 18779 5871 18785
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 8214 18825 8242 18856
rect 9398 18844 9404 18856
rect 9456 18844 9462 18896
rect 12891 18887 12949 18893
rect 12891 18853 12903 18887
rect 12937 18884 12949 18887
rect 13354 18884 13360 18896
rect 12937 18856 13360 18884
rect 12937 18853 12949 18856
rect 12891 18847 12949 18853
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 15470 18884 15476 18896
rect 15383 18856 15476 18884
rect 15470 18844 15476 18856
rect 15528 18884 15534 18896
rect 18417 18887 18475 18893
rect 18417 18884 18429 18887
rect 15528 18856 18429 18884
rect 15528 18844 15534 18856
rect 18417 18853 18429 18856
rect 18463 18853 18475 18887
rect 18417 18847 18475 18853
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 8168 18819 8242 18825
rect 7607 18788 8064 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 3421 18751 3479 18757
rect 3421 18748 3433 18751
rect 2455 18720 3433 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 3421 18717 3433 18720
rect 3467 18748 3479 18751
rect 3786 18748 3792 18760
rect 3467 18720 3792 18748
rect 3467 18717 3479 18720
rect 3421 18711 3479 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 4154 18748 4160 18760
rect 4115 18720 4160 18748
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 4264 18720 4445 18748
rect 2222 18640 2228 18692
rect 2280 18680 2286 18692
rect 3142 18680 3148 18692
rect 2280 18652 3148 18680
rect 2280 18640 2286 18652
rect 3142 18640 3148 18652
rect 3200 18680 3206 18692
rect 4264 18680 4292 18720
rect 4433 18717 4445 18720
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 8036 18748 8064 18788
rect 8168 18785 8180 18819
rect 8214 18788 8242 18819
rect 8754 18816 8760 18828
rect 8715 18788 8760 18816
rect 8214 18785 8226 18788
rect 8168 18779 8226 18785
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9548 18788 9689 18816
rect 9548 18776 9554 18788
rect 9677 18785 9689 18788
rect 9723 18816 9735 18819
rect 11057 18819 11115 18825
rect 11057 18816 11069 18819
rect 9723 18788 11069 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 11057 18785 11069 18788
rect 11103 18785 11115 18819
rect 11057 18779 11115 18785
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18816 11299 18819
rect 11790 18816 11796 18828
rect 11287 18788 11796 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18816 13507 18819
rect 14274 18816 14280 18828
rect 13495 18788 14280 18816
rect 13495 18785 13507 18788
rect 13449 18779 13507 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 16850 18816 16856 18828
rect 16811 18788 16856 18816
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 17310 18816 17316 18828
rect 17271 18788 17316 18816
rect 17310 18776 17316 18788
rect 17368 18776 17374 18828
rect 19058 18816 19064 18828
rect 19019 18788 19064 18816
rect 19058 18776 19064 18788
rect 19116 18776 19122 18828
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 5767 18720 7972 18748
rect 8036 18720 8401 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 7944 18692 7972 18720
rect 8389 18717 8401 18720
rect 8435 18748 8447 18751
rect 9030 18748 9036 18760
rect 8435 18720 9036 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 10134 18748 10140 18760
rect 10091 18720 10140 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18748 12587 18751
rect 13722 18748 13728 18760
rect 12575 18720 13728 18748
rect 12575 18717 12587 18720
rect 12529 18711 12587 18717
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 15378 18748 15384 18760
rect 15339 18720 15384 18748
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15654 18748 15660 18760
rect 15615 18720 15660 18748
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 6733 18683 6791 18689
rect 6733 18680 6745 18683
rect 3200 18652 4292 18680
rect 4632 18652 6745 18680
rect 3200 18640 3206 18652
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 1544 18584 1593 18612
rect 1544 18572 1550 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 4632 18612 4660 18652
rect 6733 18649 6745 18652
rect 6779 18649 6791 18683
rect 6733 18643 6791 18649
rect 7926 18640 7932 18692
rect 7984 18680 7990 18692
rect 11425 18683 11483 18689
rect 11425 18680 11437 18683
rect 7984 18652 11437 18680
rect 7984 18640 7990 18652
rect 11425 18649 11437 18652
rect 11471 18649 11483 18683
rect 11425 18643 11483 18649
rect 11606 18640 11612 18692
rect 11664 18680 11670 18692
rect 12345 18683 12403 18689
rect 12345 18680 12357 18683
rect 11664 18652 12357 18680
rect 11664 18640 11670 18652
rect 12345 18649 12357 18652
rect 12391 18680 12403 18683
rect 12802 18680 12808 18692
rect 12391 18652 12808 18680
rect 12391 18649 12403 18652
rect 12345 18643 12403 18649
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 7006 18612 7012 18624
rect 3568 18584 4660 18612
rect 6967 18584 7012 18612
rect 3568 18572 3574 18584
rect 7006 18572 7012 18584
rect 7064 18612 7070 18624
rect 7650 18612 7656 18624
rect 7064 18584 7656 18612
rect 7064 18572 7070 18584
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 8294 18612 8300 18624
rect 8255 18584 8300 18612
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 8352 18584 9321 18612
rect 8352 18572 8358 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9309 18575 9367 18581
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9674 18612 9680 18624
rect 9456 18584 9680 18612
rect 9456 18572 9462 18584
rect 9674 18572 9680 18584
rect 9732 18612 9738 18624
rect 9815 18615 9873 18621
rect 9815 18612 9827 18615
rect 9732 18584 9827 18612
rect 9732 18572 9738 18584
rect 9815 18581 9827 18584
rect 9861 18581 9873 18615
rect 9950 18612 9956 18624
rect 9911 18584 9956 18612
rect 9815 18575 9873 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10778 18612 10784 18624
rect 10739 18584 10784 18612
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 11790 18612 11796 18624
rect 11751 18584 11796 18612
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 14366 18612 14372 18624
rect 14327 18584 14372 18612
rect 14366 18572 14372 18584
rect 14424 18572 14430 18624
rect 18138 18612 18144 18624
rect 18099 18584 18144 18612
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2406 18408 2412 18420
rect 2367 18380 2412 18408
rect 2406 18368 2412 18380
rect 2464 18368 2470 18420
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 2869 18411 2927 18417
rect 2869 18408 2881 18411
rect 2556 18380 2881 18408
rect 2556 18368 2562 18380
rect 2869 18377 2881 18380
rect 2915 18377 2927 18411
rect 2869 18371 2927 18377
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 4246 18408 4252 18420
rect 4203 18380 4252 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 1486 18136 1492 18148
rect 1447 18108 1492 18136
rect 1486 18096 1492 18108
rect 1544 18096 1550 18148
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18136 1639 18139
rect 1670 18136 1676 18148
rect 1627 18108 1676 18136
rect 1627 18105 1639 18108
rect 1581 18099 1639 18105
rect 1670 18096 1676 18108
rect 1728 18096 1734 18148
rect 2133 18139 2191 18145
rect 2133 18105 2145 18139
rect 2179 18136 2191 18139
rect 2682 18136 2688 18148
rect 2179 18108 2688 18136
rect 2179 18105 2191 18108
rect 2133 18099 2191 18105
rect 2682 18096 2688 18108
rect 2740 18096 2746 18148
rect 2884 18136 2912 18371
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 5813 18411 5871 18417
rect 5813 18408 5825 18411
rect 4856 18380 5825 18408
rect 4856 18368 4862 18380
rect 5813 18377 5825 18380
rect 5859 18408 5871 18411
rect 6546 18408 6552 18420
rect 5859 18380 6552 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10486 18411 10544 18417
rect 10486 18408 10498 18411
rect 9732 18380 10498 18408
rect 9732 18368 9738 18380
rect 10486 18377 10498 18380
rect 10532 18408 10544 18411
rect 10778 18408 10784 18420
rect 10532 18380 10784 18408
rect 10532 18377 10544 18380
rect 10486 18371 10544 18377
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 10962 18408 10968 18420
rect 10923 18380 10968 18408
rect 10962 18368 10968 18380
rect 11020 18368 11026 18420
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 12216 18380 12909 18408
rect 12216 18368 12222 18380
rect 12897 18377 12909 18380
rect 12943 18408 12955 18411
rect 13446 18408 13452 18420
rect 12943 18380 13452 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 15381 18411 15439 18417
rect 15381 18377 15393 18411
rect 15427 18408 15439 18411
rect 15470 18408 15476 18420
rect 15427 18380 15476 18408
rect 15427 18377 15439 18380
rect 15381 18371 15439 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 16850 18408 16856 18420
rect 15764 18380 16856 18408
rect 4709 18343 4767 18349
rect 4709 18309 4721 18343
rect 4755 18340 4767 18343
rect 5258 18340 5264 18352
rect 4755 18312 5264 18340
rect 4755 18309 4767 18312
rect 4709 18303 4767 18309
rect 5258 18300 5264 18312
rect 5316 18340 5322 18352
rect 6178 18340 6184 18352
rect 5316 18312 6184 18340
rect 5316 18300 5322 18312
rect 6178 18300 6184 18312
rect 6236 18300 6242 18352
rect 9490 18300 9496 18352
rect 9548 18340 9554 18352
rect 10318 18340 10324 18352
rect 9548 18312 10324 18340
rect 9548 18300 9554 18312
rect 10318 18300 10324 18312
rect 10376 18300 10382 18352
rect 10597 18343 10655 18349
rect 10597 18309 10609 18343
rect 10643 18340 10655 18343
rect 10643 18312 11008 18340
rect 10643 18309 10655 18312
rect 10597 18303 10655 18309
rect 10980 18284 11008 18312
rect 12526 18300 12532 18352
rect 12584 18349 12590 18352
rect 12584 18343 12633 18349
rect 12584 18309 12587 18343
rect 12621 18309 12633 18343
rect 12584 18303 12633 18309
rect 12713 18343 12771 18349
rect 12713 18309 12725 18343
rect 12759 18309 12771 18343
rect 12713 18303 12771 18309
rect 12584 18300 12590 18303
rect 3142 18272 3148 18284
rect 3103 18244 3148 18272
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 3418 18272 3424 18284
rect 3379 18244 3424 18272
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 7006 18272 7012 18284
rect 6604 18244 7012 18272
rect 6604 18232 6610 18244
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 6840 18213 6868 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8294 18272 8300 18284
rect 8159 18244 8300 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 8294 18232 8300 18244
rect 8352 18272 8358 18284
rect 9582 18272 9588 18284
rect 8352 18244 9588 18272
rect 8352 18232 8358 18244
rect 9582 18232 9588 18244
rect 9640 18272 9646 18284
rect 9950 18272 9956 18284
rect 9640 18244 9956 18272
rect 9640 18232 9646 18244
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 10134 18272 10140 18284
rect 10047 18244 10140 18272
rect 10134 18232 10140 18244
rect 10192 18272 10198 18284
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10192 18244 10701 18272
rect 10192 18232 10198 18244
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 12728 18272 12756 18303
rect 13538 18300 13544 18352
rect 13596 18340 13602 18352
rect 15764 18340 15792 18380
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 19058 18408 19064 18420
rect 19019 18380 19064 18408
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 13596 18312 15792 18340
rect 13596 18300 13602 18312
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 18690 18340 18696 18352
rect 15896 18312 15976 18340
rect 18651 18312 18696 18340
rect 15896 18300 15902 18312
rect 11808 18244 12756 18272
rect 4893 18207 4951 18213
rect 4893 18204 4905 18207
rect 4764 18176 4905 18204
rect 4764 18164 4770 18176
rect 4893 18173 4905 18176
rect 4939 18204 4951 18207
rect 6825 18207 6883 18213
rect 4939 18176 6684 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 3237 18139 3295 18145
rect 3237 18136 3249 18139
rect 2884 18108 3249 18136
rect 3237 18105 3249 18108
rect 3283 18136 3295 18139
rect 4982 18136 4988 18148
rect 3283 18108 4988 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 5258 18068 5264 18080
rect 5219 18040 5264 18068
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 6546 18068 6552 18080
rect 5500 18040 6552 18068
rect 5500 18028 5506 18040
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 6656 18068 6684 18176
rect 6825 18173 6837 18207
rect 6871 18173 6883 18207
rect 7282 18204 7288 18216
rect 7243 18176 7288 18204
rect 6825 18167 6883 18173
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8588 18176 8861 18204
rect 8588 18080 8616 18176
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 9858 18204 9864 18216
rect 8849 18167 8907 18173
rect 9646 18176 9864 18204
rect 9493 18139 9551 18145
rect 9493 18105 9505 18139
rect 9539 18136 9551 18139
rect 9646 18136 9674 18176
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 9539 18108 9674 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 6917 18071 6975 18077
rect 6917 18068 6929 18071
rect 6656 18040 6929 18068
rect 6917 18037 6929 18040
rect 6963 18037 6975 18071
rect 8570 18068 8576 18080
rect 8531 18040 8576 18068
rect 6917 18031 6975 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 10042 18068 10048 18080
rect 9907 18040 10048 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10042 18028 10048 18040
rect 10100 18068 10106 18080
rect 10152 18077 10180 18232
rect 10226 18164 10232 18216
rect 10284 18204 10290 18216
rect 11808 18213 11836 18244
rect 12802 18232 12808 18284
rect 12860 18272 12866 18284
rect 14366 18272 14372 18284
rect 12860 18244 12905 18272
rect 13786 18244 14372 18272
rect 12860 18232 12866 18244
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 10284 18176 11805 18204
rect 10284 18164 10290 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 12526 18204 12532 18216
rect 11793 18167 11851 18173
rect 11900 18176 12532 18204
rect 10318 18136 10324 18148
rect 10231 18108 10324 18136
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 11425 18139 11483 18145
rect 11425 18136 11437 18139
rect 10836 18108 11437 18136
rect 10836 18096 10842 18108
rect 11425 18105 11437 18108
rect 11471 18136 11483 18139
rect 11900 18136 11928 18176
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 12820 18176 13369 18204
rect 12434 18136 12440 18148
rect 11471 18108 11928 18136
rect 11992 18108 12440 18136
rect 11471 18105 11483 18108
rect 11425 18099 11483 18105
rect 10137 18071 10195 18077
rect 10137 18068 10149 18071
rect 10100 18040 10149 18068
rect 10100 18028 10106 18040
rect 10137 18037 10149 18040
rect 10183 18037 10195 18071
rect 10336 18068 10364 18096
rect 11992 18068 12020 18108
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 12544 18136 12572 18164
rect 12820 18136 12848 18176
rect 13357 18173 13369 18176
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 12544 18108 12848 18136
rect 13262 18096 13268 18148
rect 13320 18136 13326 18148
rect 13786 18136 13814 18244
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 15948 18281 15976 18312
rect 18690 18300 18696 18312
rect 18748 18300 18754 18352
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18241 15991 18275
rect 18138 18272 18144 18284
rect 18099 18244 18144 18272
rect 15933 18235 15991 18241
rect 18138 18232 18144 18244
rect 18196 18272 18202 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 18196 18244 19625 18272
rect 18196 18232 18202 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 13320 18108 13814 18136
rect 14185 18139 14243 18145
rect 13320 18096 13326 18108
rect 14185 18105 14197 18139
rect 14231 18136 14243 18139
rect 14458 18136 14464 18148
rect 14231 18108 14464 18136
rect 14231 18105 14243 18108
rect 14185 18099 14243 18105
rect 14458 18096 14464 18108
rect 14516 18096 14522 18148
rect 16025 18139 16083 18145
rect 16025 18105 16037 18139
rect 16071 18105 16083 18139
rect 16574 18136 16580 18148
rect 16535 18108 16580 18136
rect 16025 18099 16083 18105
rect 10336 18040 12020 18068
rect 12253 18071 12311 18077
rect 10137 18031 10195 18037
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 13354 18068 13360 18080
rect 12299 18040 13360 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 13541 18071 13599 18077
rect 13541 18037 13553 18071
rect 13587 18068 13599 18071
rect 15562 18068 15568 18080
rect 13587 18040 15568 18068
rect 13587 18037 13599 18040
rect 13541 18031 13599 18037
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 15746 18068 15752 18080
rect 15659 18040 15752 18068
rect 15746 18028 15752 18040
rect 15804 18068 15810 18080
rect 16040 18068 16068 18099
rect 16574 18096 16580 18108
rect 16632 18096 16638 18148
rect 17865 18139 17923 18145
rect 17865 18105 17877 18139
rect 17911 18136 17923 18139
rect 18230 18136 18236 18148
rect 17911 18108 18236 18136
rect 17911 18105 17923 18108
rect 17865 18099 17923 18105
rect 18230 18096 18236 18108
rect 18288 18096 18294 18148
rect 17586 18068 17592 18080
rect 15804 18040 17592 18068
rect 15804 18028 15810 18040
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3142 17864 3148 17876
rect 3103 17836 3148 17864
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 4706 17864 4712 17876
rect 4667 17836 4712 17864
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 4982 17824 4988 17876
rect 5040 17864 5046 17876
rect 5721 17867 5779 17873
rect 5721 17864 5733 17867
rect 5040 17836 5733 17864
rect 5040 17824 5046 17836
rect 5721 17833 5733 17836
rect 5767 17833 5779 17867
rect 5994 17864 6000 17876
rect 5955 17836 6000 17864
rect 5721 17827 5779 17833
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 8481 17867 8539 17873
rect 8481 17833 8493 17867
rect 8527 17864 8539 17867
rect 9398 17864 9404 17876
rect 8527 17836 9404 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 12492 17836 13093 17864
rect 12492 17824 12498 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13446 17864 13452 17876
rect 13407 17836 13452 17864
rect 13081 17827 13139 17833
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 13722 17864 13728 17876
rect 13683 17836 13728 17864
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 15105 17867 15163 17873
rect 15105 17864 15117 17867
rect 13872 17836 15117 17864
rect 13872 17824 13878 17836
rect 15105 17833 15117 17836
rect 15151 17864 15163 17867
rect 15378 17864 15384 17876
rect 15151 17836 15384 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 15838 17864 15844 17876
rect 15799 17836 15844 17864
rect 15838 17824 15844 17836
rect 15896 17824 15902 17876
rect 16390 17824 16396 17876
rect 16448 17864 16454 17876
rect 16761 17867 16819 17873
rect 16761 17864 16773 17867
rect 16448 17836 16773 17864
rect 16448 17824 16454 17836
rect 16761 17833 16773 17836
rect 16807 17833 16819 17867
rect 19334 17864 19340 17876
rect 16761 17827 16819 17833
rect 18115 17836 19340 17864
rect 2130 17796 2136 17808
rect 2091 17768 2136 17796
rect 2130 17756 2136 17768
rect 2188 17756 2194 17808
rect 5163 17799 5221 17805
rect 5163 17765 5175 17799
rect 5209 17796 5221 17799
rect 5258 17796 5264 17808
rect 5209 17768 5264 17796
rect 5209 17765 5221 17768
rect 5163 17759 5221 17765
rect 5258 17756 5264 17768
rect 5316 17756 5322 17808
rect 9306 17756 9312 17808
rect 9364 17796 9370 17808
rect 10229 17799 10287 17805
rect 10229 17796 10241 17799
rect 9364 17768 10241 17796
rect 9364 17756 9370 17768
rect 10229 17765 10241 17768
rect 10275 17796 10287 17799
rect 10594 17796 10600 17808
rect 10275 17768 10600 17796
rect 10275 17765 10287 17768
rect 10229 17759 10287 17765
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 10965 17799 11023 17805
rect 10965 17765 10977 17799
rect 11011 17796 11023 17799
rect 12894 17796 12900 17808
rect 11011 17768 12900 17796
rect 11011 17765 11023 17768
rect 10965 17759 11023 17765
rect 12894 17756 12900 17768
rect 12952 17756 12958 17808
rect 13464 17796 13492 17824
rect 18115 17796 18143 17836
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 18322 17796 18328 17808
rect 13464 17768 13814 17796
rect 7466 17728 7472 17740
rect 7427 17700 7472 17728
rect 7466 17688 7472 17700
rect 7524 17728 7530 17740
rect 8754 17728 8760 17740
rect 7524 17700 8760 17728
rect 7524 17688 7530 17700
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 10318 17728 10324 17740
rect 10286 17700 10324 17728
rect 10318 17688 10324 17700
rect 10376 17737 10382 17740
rect 10376 17731 10434 17737
rect 10376 17697 10388 17731
rect 10422 17728 10434 17731
rect 10778 17728 10784 17740
rect 10422 17700 10784 17728
rect 10422 17697 10434 17700
rect 10376 17691 10434 17697
rect 10376 17688 10382 17691
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 12032 17700 12081 17728
rect 12032 17688 12038 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12526 17728 12532 17740
rect 12487 17700 12532 17728
rect 12069 17691 12127 17697
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2498 17660 2504 17672
rect 2087 17632 2504 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 2682 17660 2688 17672
rect 2595 17632 2688 17660
rect 2682 17620 2688 17632
rect 2740 17660 2746 17672
rect 3050 17660 3056 17672
rect 2740 17632 3056 17660
rect 2740 17620 2746 17632
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4801 17663 4859 17669
rect 4801 17660 4813 17663
rect 4212 17632 4813 17660
rect 4212 17620 4218 17632
rect 4801 17629 4813 17632
rect 4847 17660 4859 17663
rect 5166 17660 5172 17672
rect 4847 17632 5172 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 6917 17595 6975 17601
rect 6917 17561 6929 17595
rect 6963 17592 6975 17595
rect 7282 17592 7288 17604
rect 6963 17564 7288 17592
rect 6963 17561 6975 17564
rect 6917 17555 6975 17561
rect 7282 17552 7288 17564
rect 7340 17592 7346 17604
rect 7742 17592 7748 17604
rect 7340 17564 7748 17592
rect 7340 17552 7346 17564
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 8128 17592 8156 17623
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10100 17632 10609 17660
rect 10100 17620 10106 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 12084 17660 12112 17691
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 13265 17731 13323 17737
rect 13265 17728 13277 17731
rect 12728 17700 13277 17728
rect 12728 17660 12756 17700
rect 13265 17697 13277 17700
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 13538 17688 13544 17740
rect 13596 17728 13602 17740
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 13596 17700 13645 17728
rect 13596 17688 13602 17700
rect 13633 17697 13645 17700
rect 13679 17697 13691 17731
rect 13786 17728 13814 17768
rect 15304 17768 18143 17796
rect 18283 17768 18328 17796
rect 15304 17740 15332 17768
rect 18322 17756 18328 17768
rect 18380 17756 18386 17808
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 13786 17700 14105 17728
rect 13633 17691 13691 17697
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 15286 17728 15292 17740
rect 15199 17700 15292 17728
rect 14093 17691 14151 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19484 17700 19717 17728
rect 19484 17688 19490 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 12084 17632 12756 17660
rect 12805 17663 12863 17669
rect 10597 17623 10655 17629
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 12851 17632 16405 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 16393 17629 16405 17632
rect 16439 17660 16451 17663
rect 16758 17660 16764 17672
rect 16439 17632 16764 17660
rect 16439 17629 16451 17632
rect 16393 17623 16451 17629
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17660 18291 17663
rect 18414 17660 18420 17672
rect 18279 17632 18420 17660
rect 18279 17629 18291 17632
rect 18233 17623 18291 17629
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 18690 17660 18696 17672
rect 18651 17632 18696 17660
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 9582 17592 9588 17604
rect 8128 17564 9588 17592
rect 9582 17552 9588 17564
rect 9640 17592 9646 17604
rect 10505 17595 10563 17601
rect 9640 17564 10272 17592
rect 9640 17552 9646 17564
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 3510 17524 3516 17536
rect 3471 17496 3516 17524
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 4246 17524 4252 17536
rect 4207 17496 4252 17524
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8720 17496 8769 17524
rect 8720 17484 8726 17496
rect 8757 17493 8769 17496
rect 8803 17493 8815 17527
rect 9490 17524 9496 17536
rect 9451 17496 9496 17524
rect 8757 17487 8815 17493
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 9950 17524 9956 17536
rect 9863 17496 9956 17524
rect 9950 17484 9956 17496
rect 10008 17524 10014 17536
rect 10134 17524 10140 17536
rect 10008 17496 10140 17524
rect 10008 17484 10014 17496
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 10244 17524 10272 17564
rect 10505 17561 10517 17595
rect 10551 17592 10563 17595
rect 10962 17592 10968 17604
rect 10551 17564 10968 17592
rect 10551 17561 10563 17564
rect 10505 17555 10563 17561
rect 10962 17552 10968 17564
rect 11020 17592 11026 17604
rect 11241 17595 11299 17601
rect 11241 17592 11253 17595
rect 11020 17564 11253 17592
rect 11020 17552 11026 17564
rect 11241 17561 11253 17564
rect 11287 17592 11299 17595
rect 11609 17595 11667 17601
rect 11609 17592 11621 17595
rect 11287 17564 11621 17592
rect 11287 17561 11299 17564
rect 11241 17555 11299 17561
rect 11609 17561 11621 17564
rect 11655 17561 11667 17595
rect 11609 17555 11667 17561
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 13814 17592 13820 17604
rect 12952 17564 13820 17592
rect 12952 17552 12958 17564
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 15473 17595 15531 17601
rect 15473 17592 15485 17595
rect 13969 17564 15485 17592
rect 12066 17524 12072 17536
rect 10244 17496 12072 17524
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 13265 17527 13323 17533
rect 13265 17493 13277 17527
rect 13311 17524 13323 17527
rect 13969 17524 13997 17564
rect 15473 17561 15485 17564
rect 15519 17561 15531 17595
rect 15473 17555 15531 17561
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 19889 17595 19947 17601
rect 19889 17592 19901 17595
rect 15620 17564 19901 17592
rect 15620 17552 15626 17564
rect 19889 17561 19901 17564
rect 19935 17561 19947 17595
rect 19889 17555 19947 17561
rect 17310 17524 17316 17536
rect 13311 17496 13997 17524
rect 17271 17496 17316 17524
rect 13311 17493 13323 17496
rect 13265 17487 13323 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 2130 17280 2136 17332
rect 2188 17320 2194 17332
rect 2501 17323 2559 17329
rect 2501 17320 2513 17323
rect 2188 17292 2513 17320
rect 2188 17280 2194 17292
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 2332 17116 2360 17292
rect 2501 17289 2513 17292
rect 2547 17320 2559 17323
rect 2547 17292 3740 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 3712 17264 3740 17292
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4893 17323 4951 17329
rect 4212 17292 4257 17320
rect 4212 17280 4218 17292
rect 4893 17289 4905 17323
rect 4939 17320 4951 17323
rect 5258 17320 5264 17332
rect 4939 17292 5264 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 5258 17280 5264 17292
rect 5316 17320 5322 17332
rect 6178 17320 6184 17332
rect 5316 17292 6184 17320
rect 5316 17280 5322 17292
rect 6178 17280 6184 17292
rect 6236 17320 6242 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6236 17292 6561 17320
rect 6236 17280 6242 17292
rect 6549 17289 6561 17292
rect 6595 17320 6607 17323
rect 7006 17320 7012 17332
rect 6595 17292 7012 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 8941 17323 8999 17329
rect 8941 17320 8953 17323
rect 8628 17292 8953 17320
rect 8628 17280 8634 17292
rect 8941 17289 8953 17292
rect 8987 17289 8999 17323
rect 8941 17283 8999 17289
rect 9953 17323 10011 17329
rect 9953 17289 9965 17323
rect 9999 17320 10011 17323
rect 10318 17320 10324 17332
rect 9999 17292 10324 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 10962 17320 10968 17332
rect 10919 17292 10968 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 12526 17320 12532 17332
rect 11287 17292 12532 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 12713 17323 12771 17329
rect 12713 17289 12725 17323
rect 12759 17320 12771 17323
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 12759 17292 13001 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 12989 17289 13001 17292
rect 13035 17320 13047 17323
rect 13170 17320 13176 17332
rect 13035 17292 13176 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17320 14611 17323
rect 15746 17320 15752 17332
rect 14599 17292 15752 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 16758 17320 16764 17332
rect 16719 17292 16764 17320
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 18230 17280 18236 17332
rect 18288 17320 18294 17332
rect 18325 17323 18383 17329
rect 18325 17320 18337 17323
rect 18288 17292 18337 17320
rect 18288 17280 18294 17292
rect 18325 17289 18337 17292
rect 18371 17289 18383 17323
rect 18325 17283 18383 17289
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 18472 17292 19073 17320
rect 18472 17280 18478 17292
rect 19061 17289 19073 17292
rect 19107 17289 19119 17323
rect 19061 17283 19119 17289
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 3605 17255 3663 17261
rect 3605 17252 3617 17255
rect 2648 17224 3617 17252
rect 2648 17212 2654 17224
rect 3605 17221 3617 17224
rect 3651 17221 3663 17255
rect 3605 17215 3663 17221
rect 3694 17212 3700 17264
rect 3752 17252 3758 17264
rect 7745 17255 7803 17261
rect 7745 17252 7757 17255
rect 3752 17224 7757 17252
rect 3752 17212 3758 17224
rect 7745 17221 7757 17224
rect 7791 17221 7803 17255
rect 7745 17215 7803 17221
rect 8202 17212 8208 17264
rect 8260 17252 8266 17264
rect 8803 17255 8861 17261
rect 8803 17252 8815 17255
rect 8260 17224 8815 17252
rect 8260 17212 8266 17224
rect 8803 17221 8815 17224
rect 8849 17221 8861 17255
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 8803 17215 8861 17221
rect 8910 17224 9137 17252
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17184 3111 17187
rect 3510 17184 3516 17196
rect 3099 17156 3516 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 3510 17144 3516 17156
rect 3568 17144 3574 17196
rect 4525 17187 4583 17193
rect 4525 17153 4537 17187
rect 4571 17184 4583 17187
rect 8018 17184 8024 17196
rect 4571 17156 8024 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 5442 17116 5448 17128
rect 2087 17088 2360 17116
rect 5403 17088 5448 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 5644 17125 5672 17156
rect 8018 17144 8024 17156
rect 8076 17184 8082 17196
rect 8910 17184 8938 17224
rect 9125 17221 9137 17224
rect 9171 17221 9183 17255
rect 10980 17252 11008 17280
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 10980 17224 11989 17252
rect 9125 17215 9183 17221
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 11977 17215 12035 17221
rect 12066 17212 12072 17264
rect 12124 17252 12130 17264
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 12124 17224 14933 17252
rect 12124 17212 12130 17224
rect 14921 17221 14933 17224
rect 14967 17252 14979 17255
rect 15286 17252 15292 17264
rect 14967 17224 15292 17252
rect 14967 17221 14979 17224
rect 14921 17215 14979 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 16025 17255 16083 17261
rect 16025 17221 16037 17255
rect 16071 17252 16083 17255
rect 16574 17252 16580 17264
rect 16071 17224 16580 17252
rect 16071 17221 16083 17224
rect 16025 17215 16083 17221
rect 16574 17212 16580 17224
rect 16632 17252 16638 17264
rect 18432 17252 18460 17280
rect 16632 17224 18460 17252
rect 16632 17212 16638 17224
rect 9030 17184 9036 17196
rect 8076 17156 8938 17184
rect 8991 17156 9036 17184
rect 8076 17144 8082 17156
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 5629 17119 5687 17125
rect 5629 17085 5641 17119
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6273 17119 6331 17125
rect 6273 17116 6285 17119
rect 5951 17088 6285 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6273 17085 6285 17088
rect 6319 17116 6331 17119
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6319 17088 6837 17116
rect 6319 17085 6331 17088
rect 6273 17079 6331 17085
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7650 17076 7656 17128
rect 7708 17116 7714 17128
rect 8662 17116 8668 17128
rect 7708 17088 8668 17116
rect 7708 17076 7714 17088
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 10778 17125 10784 17128
rect 10744 17119 10784 17125
rect 10744 17085 10756 17119
rect 10744 17079 10784 17085
rect 10778 17076 10784 17079
rect 10836 17076 10842 17128
rect 10980 17116 11008 17147
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11296 17156 11713 17184
rect 11296 17144 11302 17156
rect 11701 17153 11713 17156
rect 11747 17184 11759 17187
rect 18230 17184 18236 17196
rect 11747 17156 18236 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 11606 17116 11612 17128
rect 10980 17088 11612 17116
rect 11606 17076 11612 17088
rect 11664 17076 11670 17128
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17116 12495 17119
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12483 17088 12725 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 3145 17051 3203 17057
rect 3145 17017 3157 17051
rect 3191 17017 3203 17051
rect 6730 17048 6736 17060
rect 3145 17011 3203 17017
rect 4126 17020 6736 17048
rect 2869 16983 2927 16989
rect 2869 16949 2881 16983
rect 2915 16980 2927 16983
rect 3160 16980 3188 17011
rect 3510 16980 3516 16992
rect 2915 16952 3516 16980
rect 2915 16949 2927 16952
rect 2869 16943 2927 16949
rect 3510 16940 3516 16952
rect 3568 16980 3574 16992
rect 4126 16980 4154 17020
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 7146 17051 7204 17057
rect 7146 17048 7158 17051
rect 7064 17020 7158 17048
rect 7064 17008 7070 17020
rect 7146 17017 7158 17020
rect 7192 17017 7204 17051
rect 8570 17048 8576 17060
rect 8531 17020 8576 17048
rect 7146 17011 7204 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 10042 17008 10048 17060
rect 10100 17048 10106 17060
rect 10229 17051 10287 17057
rect 10229 17048 10241 17051
rect 10100 17020 10241 17048
rect 10100 17008 10106 17020
rect 10229 17017 10241 17020
rect 10275 17017 10287 17051
rect 10594 17048 10600 17060
rect 10507 17020 10600 17048
rect 10229 17011 10287 17017
rect 10594 17008 10600 17020
rect 10652 17048 10658 17060
rect 11238 17048 11244 17060
rect 10652 17020 11244 17048
rect 10652 17008 10658 17020
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 3568 16952 4154 16980
rect 3568 16940 3574 16952
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 7466 16980 7472 16992
rect 6880 16952 7472 16980
rect 6880 16940 6886 16952
rect 7466 16940 7472 16952
rect 7524 16980 7530 16992
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7524 16952 8033 16980
rect 7524 16940 7530 16952
rect 8021 16949 8033 16952
rect 8067 16949 8079 16983
rect 8021 16943 8079 16949
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 12452 16980 12480 17079
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 13633 17119 13691 17125
rect 13633 17116 13645 17119
rect 12860 17088 13645 17116
rect 12860 17076 12866 17088
rect 13633 17085 13645 17088
rect 13679 17116 13691 17119
rect 14642 17116 14648 17128
rect 13679 17088 14648 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 16942 17116 16948 17128
rect 16903 17088 16948 17116
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 17310 17076 17316 17128
rect 17368 17116 17374 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 17368 17088 17509 17116
rect 17368 17076 17374 17088
rect 17497 17085 17509 17088
rect 17543 17116 17555 17119
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17543 17088 17877 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 17865 17085 17877 17088
rect 17911 17116 17923 17119
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17911 17088 18153 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 18141 17085 18153 17088
rect 18187 17116 18199 17119
rect 18322 17116 18328 17128
rect 18187 17088 18328 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 13954 17051 14012 17057
rect 13954 17017 13966 17051
rect 14000 17017 14012 17051
rect 15470 17048 15476 17060
rect 15431 17020 15476 17048
rect 13954 17011 14012 17017
rect 8812 16952 12480 16980
rect 12621 16983 12679 16989
rect 8812 16940 8818 16952
rect 12621 16949 12633 16983
rect 12667 16980 12679 16983
rect 12710 16980 12716 16992
rect 12667 16952 12716 16980
rect 12667 16949 12679 16952
rect 12621 16943 12679 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 13446 16980 13452 16992
rect 13407 16952 13452 16980
rect 13446 16940 13452 16952
rect 13504 16980 13510 16992
rect 13969 16980 13997 17011
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 15565 17051 15623 17057
rect 15565 17017 15577 17051
rect 15611 17048 15623 17051
rect 17218 17048 17224 17060
rect 15611 17020 17224 17048
rect 15611 17017 15623 17020
rect 15565 17011 15623 17017
rect 13504 16952 13997 16980
rect 15289 16983 15347 16989
rect 13504 16940 13510 16952
rect 15289 16949 15301 16983
rect 15335 16980 15347 16983
rect 15580 16980 15608 17011
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 22094 17048 22100 17060
rect 17328 17020 22100 17048
rect 16390 16980 16396 16992
rect 15335 16952 15608 16980
rect 16351 16952 16396 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 17083 16983 17141 16989
rect 17083 16949 17095 16983
rect 17129 16980 17141 16983
rect 17328 16980 17356 17020
rect 22094 17008 22100 17020
rect 22152 17008 22158 17060
rect 17129 16952 17356 16980
rect 17129 16949 17141 16952
rect 17083 16943 17141 16949
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19705 16983 19763 16989
rect 19705 16980 19717 16983
rect 19484 16952 19717 16980
rect 19484 16940 19490 16952
rect 19705 16949 19717 16952
rect 19751 16949 19763 16983
rect 19705 16943 19763 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 3694 16776 3700 16788
rect 3099 16748 3700 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 6178 16776 6184 16788
rect 6139 16748 6184 16776
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 6730 16776 6736 16788
rect 6691 16748 6736 16776
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 6840 16748 7665 16776
rect 2133 16711 2191 16717
rect 2133 16677 2145 16711
rect 2179 16708 2191 16711
rect 2774 16708 2780 16720
rect 2179 16680 2780 16708
rect 2179 16677 2191 16680
rect 2133 16671 2191 16677
rect 2774 16668 2780 16680
rect 2832 16668 2838 16720
rect 3602 16668 3608 16720
rect 3660 16708 3666 16720
rect 4985 16711 5043 16717
rect 4985 16708 4997 16711
rect 3660 16680 4997 16708
rect 3660 16668 3666 16680
rect 4985 16677 4997 16680
rect 5031 16677 5043 16711
rect 4985 16671 5043 16677
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 4212 16612 4261 16640
rect 4212 16600 4218 16612
rect 4249 16609 4261 16612
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16640 5871 16643
rect 6270 16640 6276 16652
rect 5859 16612 6276 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 6270 16600 6276 16612
rect 6328 16640 6334 16652
rect 6840 16640 6868 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 7800 16748 10333 16776
rect 7800 16736 7806 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 11149 16779 11207 16785
rect 10321 16739 10379 16745
rect 10428 16748 11008 16776
rect 7101 16711 7159 16717
rect 7101 16677 7113 16711
rect 7147 16708 7159 16711
rect 7190 16708 7196 16720
rect 7147 16680 7196 16708
rect 7147 16677 7159 16680
rect 7101 16671 7159 16677
rect 7190 16668 7196 16680
rect 7248 16708 7254 16720
rect 7248 16680 7604 16708
rect 7248 16668 7254 16680
rect 7576 16649 7604 16680
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 9030 16708 9036 16720
rect 8352 16680 9036 16708
rect 8352 16668 8358 16680
rect 9030 16668 9036 16680
rect 9088 16708 9094 16720
rect 9125 16711 9183 16717
rect 9125 16708 9137 16711
rect 9088 16680 9137 16708
rect 9088 16668 9094 16680
rect 9125 16677 9137 16680
rect 9171 16677 9183 16711
rect 9125 16671 9183 16677
rect 9398 16668 9404 16720
rect 9456 16708 9462 16720
rect 10428 16708 10456 16748
rect 10778 16708 10784 16720
rect 9456 16680 10456 16708
rect 10739 16680 10784 16708
rect 9456 16668 9462 16680
rect 10778 16668 10784 16680
rect 10836 16668 10842 16720
rect 10980 16708 11008 16748
rect 11149 16745 11161 16779
rect 11195 16776 11207 16779
rect 11238 16776 11244 16788
rect 11195 16748 11244 16776
rect 11195 16745 11207 16748
rect 11149 16739 11207 16745
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 12989 16779 13047 16785
rect 12989 16776 13001 16779
rect 12584 16748 13001 16776
rect 12584 16736 12590 16748
rect 12989 16745 13001 16748
rect 13035 16745 13047 16779
rect 13538 16776 13544 16788
rect 13499 16748 13544 16776
rect 12989 16739 13047 16745
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 13630 16736 13636 16788
rect 13688 16776 13694 16788
rect 14642 16776 14648 16788
rect 13688 16748 13768 16776
rect 14603 16748 14648 16776
rect 13688 16736 13694 16748
rect 12710 16708 12716 16720
rect 10980 16680 12716 16708
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 13740 16717 13768 16748
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 13725 16711 13783 16717
rect 13725 16677 13737 16711
rect 13771 16677 13783 16711
rect 13725 16671 13783 16677
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 16761 16711 16819 16717
rect 13872 16680 13917 16708
rect 13872 16668 13878 16680
rect 16761 16677 16773 16711
rect 16807 16708 16819 16711
rect 17034 16708 17040 16720
rect 16807 16680 17040 16708
rect 16807 16677 16819 16680
rect 16761 16671 16819 16677
rect 17034 16668 17040 16680
rect 17092 16708 17098 16720
rect 18141 16711 18199 16717
rect 18141 16708 18153 16711
rect 17092 16680 18153 16708
rect 17092 16668 17098 16680
rect 18141 16677 18153 16680
rect 18187 16677 18199 16711
rect 18141 16671 18199 16677
rect 6328 16612 6868 16640
rect 7561 16643 7619 16649
rect 6328 16600 6334 16612
rect 7561 16609 7573 16643
rect 7607 16609 7619 16643
rect 8018 16640 8024 16652
rect 7979 16612 8024 16640
rect 7561 16603 7619 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 8812 16612 9689 16640
rect 8812 16600 8818 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11756 16612 11989 16640
rect 11756 16600 11762 16612
rect 11977 16609 11989 16612
rect 12023 16609 12035 16643
rect 12434 16640 12440 16652
rect 12395 16612 12440 16640
rect 11977 16603 12035 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15470 16600 15476 16652
rect 15528 16600 15534 16652
rect 18782 16640 18788 16652
rect 18743 16612 18788 16640
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16541 2099 16575
rect 2498 16572 2504 16584
rect 2459 16544 2504 16572
rect 2041 16535 2099 16541
rect 2056 16504 2084 16535
rect 2498 16532 2504 16544
rect 2556 16572 2562 16584
rect 3697 16575 3755 16581
rect 3697 16572 3709 16575
rect 2556 16544 3709 16572
rect 2556 16532 2562 16544
rect 3697 16541 3709 16544
rect 3743 16541 3755 16575
rect 3697 16535 3755 16541
rect 4396 16575 4454 16581
rect 4396 16541 4408 16575
rect 4442 16572 4454 16575
rect 4522 16572 4528 16584
rect 4442 16544 4528 16572
rect 4442 16541 4454 16544
rect 4396 16535 4454 16541
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 4614 16532 4620 16584
rect 4672 16572 4678 16584
rect 9306 16572 9312 16584
rect 4672 16544 9312 16572
rect 4672 16532 4678 16544
rect 9306 16532 9312 16544
rect 9364 16572 9370 16584
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 9364 16544 10057 16572
rect 9364 16532 9370 16544
rect 10045 16541 10057 16544
rect 10091 16572 10103 16575
rect 10502 16572 10508 16584
rect 10091 16544 10508 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 12710 16572 12716 16584
rect 12671 16544 12716 16572
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 14366 16572 14372 16584
rect 14327 16544 14372 16572
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 15488 16572 15516 16600
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 14516 16544 15761 16572
rect 14516 16532 14522 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 16666 16572 16672 16584
rect 16627 16544 16672 16572
rect 15749 16535 15807 16541
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16942 16572 16948 16584
rect 16903 16544 16948 16572
rect 16942 16532 16948 16544
rect 17000 16572 17006 16584
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 17000 16544 17601 16572
rect 17000 16532 17006 16544
rect 17589 16541 17601 16544
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 2314 16504 2320 16516
rect 2056 16476 2320 16504
rect 2314 16464 2320 16476
rect 2372 16464 2378 16516
rect 3326 16464 3332 16516
rect 3384 16504 3390 16516
rect 3602 16504 3608 16516
rect 3384 16476 3608 16504
rect 3384 16464 3390 16476
rect 3602 16464 3608 16476
rect 3660 16464 3666 16516
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9088 16476 10732 16504
rect 9088 16464 9094 16476
rect 1762 16436 1768 16448
rect 1723 16408 1768 16436
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 3418 16436 3424 16448
rect 3379 16408 3424 16436
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 4798 16436 4804 16448
rect 4571 16408 4804 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 5353 16439 5411 16445
rect 5353 16405 5365 16439
rect 5399 16436 5411 16439
rect 5442 16436 5448 16448
rect 5399 16408 5448 16436
rect 5399 16405 5411 16408
rect 5353 16399 5411 16405
rect 5442 16396 5448 16408
rect 5500 16436 5506 16448
rect 5629 16439 5687 16445
rect 5629 16436 5641 16439
rect 5500 16408 5641 16436
rect 5500 16396 5506 16408
rect 5629 16405 5641 16408
rect 5675 16405 5687 16439
rect 5629 16399 5687 16405
rect 7469 16439 7527 16445
rect 7469 16405 7481 16439
rect 7515 16436 7527 16439
rect 8202 16436 8208 16448
rect 7515 16408 8208 16436
rect 7515 16405 7527 16408
rect 7469 16399 7527 16405
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 8754 16436 8760 16448
rect 8715 16408 8760 16436
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9815 16439 9873 16445
rect 9815 16436 9827 16439
rect 9456 16408 9827 16436
rect 9456 16396 9462 16408
rect 9815 16405 9827 16408
rect 9861 16405 9873 16439
rect 9950 16436 9956 16448
rect 9911 16408 9956 16436
rect 9815 16399 9873 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10704 16436 10732 16476
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 11793 16507 11851 16513
rect 11793 16504 11805 16507
rect 10836 16476 11805 16504
rect 10836 16464 10842 16476
rect 11793 16473 11805 16476
rect 11839 16504 11851 16507
rect 11974 16504 11980 16516
rect 11839 16476 11980 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 11974 16464 11980 16476
rect 12032 16464 12038 16516
rect 11517 16439 11575 16445
rect 11517 16436 11529 16439
rect 10704 16408 11529 16436
rect 11517 16405 11529 16408
rect 11563 16436 11575 16439
rect 11606 16436 11612 16448
rect 11563 16408 11612 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 11606 16396 11612 16408
rect 11664 16436 11670 16448
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 11664 16408 15485 16436
rect 11664 16396 11670 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 15473 16399 15531 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4341 16235 4399 16241
rect 4341 16232 4353 16235
rect 4212 16204 4353 16232
rect 4212 16192 4218 16204
rect 4341 16201 4353 16204
rect 4387 16232 4399 16235
rect 7650 16232 7656 16244
rect 4387 16204 7656 16232
rect 4387 16201 4399 16204
rect 4341 16195 4399 16201
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 8294 16232 8300 16244
rect 8255 16204 8300 16232
rect 8294 16192 8300 16204
rect 8352 16232 8358 16244
rect 10502 16232 10508 16244
rect 8352 16204 9168 16232
rect 10463 16204 10508 16232
rect 8352 16192 8358 16204
rect 2866 16124 2872 16176
rect 2924 16164 2930 16176
rect 6178 16164 6184 16176
rect 2924 16136 3740 16164
rect 6139 16136 6184 16164
rect 2924 16124 2930 16136
rect 3418 16096 3424 16108
rect 3379 16068 3424 16096
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 3712 16105 3740 16136
rect 6178 16124 6184 16136
rect 6236 16124 6242 16176
rect 7190 16124 7196 16176
rect 7248 16164 7254 16176
rect 7837 16167 7895 16173
rect 7837 16164 7849 16167
rect 7248 16136 7849 16164
rect 7248 16124 7254 16136
rect 7837 16133 7849 16136
rect 7883 16133 7895 16167
rect 9030 16164 9036 16176
rect 8991 16136 9036 16164
rect 7837 16127 7895 16133
rect 9030 16124 9036 16136
rect 9088 16124 9094 16176
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 4798 16096 4804 16108
rect 4711 16068 4804 16096
rect 3697 16059 3755 16065
rect 4798 16056 4804 16068
rect 4856 16096 4862 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 4856 16068 8401 16096
rect 4856 16056 4862 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 8901 16056 8907 16108
rect 8959 16096 8965 16108
rect 9140 16105 9168 16204
rect 10502 16192 10508 16204
rect 10560 16232 10566 16244
rect 15286 16232 15292 16244
rect 10560 16204 15292 16232
rect 10560 16192 10566 16204
rect 15286 16192 15292 16204
rect 15344 16232 15350 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15344 16204 15945 16232
rect 15344 16192 15350 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 15933 16195 15991 16201
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 18230 16232 18236 16244
rect 18191 16204 18236 16232
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 18877 16235 18935 16241
rect 18877 16232 18889 16235
rect 18840 16204 18889 16232
rect 18840 16192 18846 16204
rect 18877 16201 18889 16204
rect 18923 16201 18935 16235
rect 18877 16195 18935 16201
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 13909 16167 13967 16173
rect 13909 16164 13921 16167
rect 13872 16136 13921 16164
rect 13872 16124 13878 16136
rect 13909 16133 13921 16136
rect 13955 16133 13967 16167
rect 13909 16127 13967 16133
rect 15657 16167 15715 16173
rect 15657 16133 15669 16167
rect 15703 16164 15715 16167
rect 16114 16164 16120 16176
rect 15703 16136 16120 16164
rect 15703 16133 15715 16136
rect 15657 16127 15715 16133
rect 9125 16099 9183 16105
rect 8959 16068 9004 16096
rect 8959 16056 8965 16068
rect 9125 16065 9137 16099
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 5442 16028 5448 16040
rect 5403 16000 5448 16028
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 5994 16028 6000 16040
rect 5767 16000 6000 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 5994 15988 6000 16000
rect 6052 16028 6058 16040
rect 7101 16031 7159 16037
rect 6052 16000 6684 16028
rect 6052 15988 6058 16000
rect 1670 15960 1676 15972
rect 1631 15932 1676 15960
rect 1670 15920 1676 15932
rect 1728 15920 1734 15972
rect 3513 15963 3571 15969
rect 3513 15929 3525 15963
rect 3559 15929 3571 15963
rect 5902 15960 5908 15972
rect 5863 15932 5908 15960
rect 3513 15923 3571 15929
rect 2774 15892 2780 15904
rect 2735 15864 2780 15892
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 2958 15852 2964 15904
rect 3016 15892 3022 15904
rect 3145 15895 3203 15901
rect 3145 15892 3157 15895
rect 3016 15864 3157 15892
rect 3016 15852 3022 15864
rect 3145 15861 3157 15864
rect 3191 15892 3203 15895
rect 3528 15892 3556 15923
rect 5902 15920 5908 15932
rect 5960 15920 5966 15972
rect 6656 15969 6684 16000
rect 7101 15997 7113 16031
rect 7147 16028 7159 16031
rect 7190 16028 7196 16040
rect 7147 16000 7196 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7377 16031 7435 16037
rect 7377 15997 7389 16031
rect 7423 16028 7435 16031
rect 9232 16028 9260 16059
rect 12710 16056 12716 16108
rect 12768 16096 12774 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12768 16068 13001 16096
rect 12768 16056 12774 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 13924 16096 13952 16127
rect 16114 16124 16120 16136
rect 16172 16164 16178 16176
rect 18800 16164 18828 16192
rect 16172 16136 18828 16164
rect 16172 16124 16178 16136
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13924 16068 14289 16096
rect 12989 16059 13047 16065
rect 14277 16065 14289 16068
rect 14323 16096 14335 16099
rect 15286 16096 15292 16108
rect 14323 16068 15292 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16096 16543 16099
rect 16666 16096 16672 16108
rect 16531 16068 16672 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 16666 16056 16672 16068
rect 16724 16096 16730 16108
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 16724 16068 17325 16096
rect 16724 16056 16730 16068
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 10778 16028 10784 16040
rect 7423 16000 9260 16028
rect 10739 16000 10784 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 6641 15963 6699 15969
rect 6641 15929 6653 15963
rect 6687 15960 6699 15963
rect 7392 15960 7420 15991
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 11238 16028 11244 16040
rect 11199 16000 11244 16028
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 16028 11575 16031
rect 14734 16028 14740 16040
rect 11563 16000 14740 16028
rect 11563 15997 11575 16000
rect 11517 15991 11575 15997
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 14981 16000 18061 16028
rect 8570 15960 8576 15972
rect 6687 15932 7420 15960
rect 8531 15932 8576 15960
rect 6687 15929 6699 15932
rect 6641 15923 6699 15929
rect 8570 15920 8576 15932
rect 8628 15920 8634 15972
rect 8754 15960 8760 15972
rect 8715 15932 8760 15960
rect 8754 15920 8760 15932
rect 8812 15960 8818 15972
rect 9674 15960 9680 15972
rect 8812 15932 9680 15960
rect 8812 15920 8818 15932
rect 9674 15920 9680 15932
rect 9732 15960 9738 15972
rect 9769 15963 9827 15969
rect 9769 15960 9781 15963
rect 9732 15932 9781 15960
rect 9732 15920 9738 15932
rect 9769 15929 9781 15932
rect 9815 15929 9827 15963
rect 11256 15960 11284 15988
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 11256 15932 11989 15960
rect 9769 15923 9827 15929
rect 11977 15929 11989 15932
rect 12023 15960 12035 15963
rect 12434 15960 12440 15972
rect 12023 15932 12440 15960
rect 12023 15929 12035 15932
rect 11977 15923 12035 15929
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 13310 15963 13368 15969
rect 13310 15960 13322 15963
rect 13004 15932 13322 15960
rect 13004 15904 13032 15932
rect 13310 15929 13322 15932
rect 13356 15960 13368 15963
rect 13446 15960 13452 15972
rect 13356 15932 13452 15960
rect 13356 15929 13368 15932
rect 13310 15923 13368 15929
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 14981 15960 15009 16000
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18095 16000 18521 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 13596 15932 15009 15960
rect 15058 15963 15116 15969
rect 13596 15920 13602 15932
rect 15058 15929 15070 15963
rect 15104 15960 15116 15963
rect 16390 15960 16396 15972
rect 15104 15932 16396 15960
rect 15104 15929 15116 15932
rect 15058 15923 15116 15929
rect 6914 15892 6920 15904
rect 3191 15864 3556 15892
rect 6875 15864 6920 15892
rect 3191 15861 3203 15864
rect 3145 15855 3203 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 8389 15895 8447 15901
rect 8389 15861 8401 15895
rect 8435 15892 8447 15895
rect 9950 15892 9956 15904
rect 8435 15864 9956 15892
rect 8435 15861 8447 15864
rect 8389 15855 8447 15861
rect 9950 15852 9956 15864
rect 10008 15892 10014 15904
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 10008 15864 10241 15892
rect 10008 15852 10014 15864
rect 10229 15861 10241 15864
rect 10275 15892 10287 15895
rect 12066 15892 12072 15904
rect 10275 15864 12072 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 12986 15892 12992 15904
rect 12943 15864 12992 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 13464 15892 13492 15920
rect 14553 15895 14611 15901
rect 14553 15892 14565 15895
rect 13464 15864 14565 15892
rect 14553 15861 14565 15864
rect 14599 15892 14611 15895
rect 15073 15892 15101 15923
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 14599 15864 15101 15892
rect 14599 15861 14611 15864
rect 14553 15855 14611 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 1486 15688 1492 15700
rect 1443 15660 1492 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 1486 15648 1492 15660
rect 1544 15648 1550 15700
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 4617 15691 4675 15697
rect 4617 15688 4629 15691
rect 4580 15660 4629 15688
rect 4580 15648 4586 15660
rect 4617 15657 4629 15660
rect 4663 15657 4675 15691
rect 4617 15651 4675 15657
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 6457 15691 6515 15697
rect 6457 15688 6469 15691
rect 5960 15660 6469 15688
rect 5960 15648 5966 15660
rect 6457 15657 6469 15660
rect 6503 15688 6515 15691
rect 7929 15691 7987 15697
rect 6503 15660 6684 15688
rect 6503 15657 6515 15660
rect 6457 15651 6515 15657
rect 2590 15620 2596 15632
rect 2551 15592 2596 15620
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 5255 15623 5313 15629
rect 5255 15589 5267 15623
rect 5301 15620 5313 15623
rect 6086 15620 6092 15632
rect 5301 15592 6092 15620
rect 5301 15589 5313 15592
rect 5255 15583 5313 15589
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 6270 15620 6276 15632
rect 6227 15592 6276 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4614 15552 4620 15564
rect 4387 15524 4620 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 6656 15561 6684 15660
rect 7929 15657 7941 15691
rect 7975 15688 7987 15691
rect 8018 15688 8024 15700
rect 7975 15660 8024 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 8202 15688 8208 15700
rect 8163 15660 8208 15688
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8536 15660 8585 15688
rect 8536 15648 8542 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 13081 15691 13139 15697
rect 13081 15688 13093 15691
rect 12768 15660 13093 15688
rect 12768 15648 12774 15660
rect 13081 15657 13093 15660
rect 13127 15657 13139 15691
rect 13081 15651 13139 15657
rect 13541 15691 13599 15697
rect 13541 15657 13553 15691
rect 13587 15688 13599 15691
rect 13630 15688 13636 15700
rect 13587 15660 13636 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 14734 15688 14740 15700
rect 14695 15660 14740 15688
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 6822 15580 6828 15632
rect 6880 15620 6886 15632
rect 6962 15623 7020 15629
rect 6962 15620 6974 15623
rect 6880 15592 6974 15620
rect 6880 15580 6886 15592
rect 6962 15589 6974 15592
rect 7008 15589 7020 15623
rect 8220 15620 8248 15648
rect 8938 15620 8944 15632
rect 8220 15592 8944 15620
rect 6962 15583 7020 15589
rect 8938 15580 8944 15592
rect 8996 15620 9002 15632
rect 9214 15620 9220 15632
rect 8996 15592 9220 15620
rect 8996 15580 9002 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 9398 15620 9404 15632
rect 9359 15592 9404 15620
rect 9398 15580 9404 15592
rect 9456 15580 9462 15632
rect 9674 15620 9680 15632
rect 9635 15592 9680 15620
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 12802 15620 12808 15632
rect 12763 15592 12808 15620
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 13814 15620 13820 15632
rect 13775 15592 13820 15620
rect 13814 15580 13820 15592
rect 13872 15580 13878 15632
rect 16114 15620 16120 15632
rect 16075 15592 16120 15620
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 16669 15623 16727 15629
rect 16669 15589 16681 15623
rect 16715 15620 16727 15623
rect 16942 15620 16948 15632
rect 16715 15592 16948 15620
rect 16715 15589 16727 15592
rect 16669 15583 16727 15589
rect 16942 15580 16948 15592
rect 17000 15580 17006 15632
rect 17218 15580 17224 15632
rect 17276 15620 17282 15632
rect 17497 15623 17555 15629
rect 17497 15620 17509 15623
rect 17276 15592 17509 15620
rect 17276 15580 17282 15592
rect 17497 15589 17509 15592
rect 17543 15589 17555 15623
rect 17497 15583 17555 15589
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15521 6699 15555
rect 6641 15515 6699 15521
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 8352 15524 8401 15552
rect 8352 15512 8358 15524
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 8570 15512 8576 15564
rect 8628 15552 8634 15564
rect 9030 15552 9036 15564
rect 8628 15524 9036 15552
rect 8628 15512 8634 15524
rect 9030 15512 9036 15524
rect 9088 15512 9094 15564
rect 10778 15552 10784 15564
rect 9692 15524 10784 15552
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15484 4951 15487
rect 5534 15484 5540 15496
rect 4939 15456 5540 15484
rect 4939 15453 4951 15456
rect 4893 15447 4951 15453
rect 5534 15444 5540 15456
rect 5592 15484 5598 15496
rect 6914 15484 6920 15496
rect 5592 15456 6920 15484
rect 5592 15444 5598 15456
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 9692 15484 9720 15524
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 12069 15555 12127 15561
rect 12069 15552 12081 15555
rect 11756 15524 12081 15552
rect 11756 15512 11762 15524
rect 12069 15521 12081 15524
rect 12115 15521 12127 15555
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12069 15515 12127 15521
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 17586 15552 17592 15564
rect 17547 15524 17592 15552
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 10042 15484 10048 15496
rect 7248 15456 9720 15484
rect 10003 15456 10048 15484
rect 7248 15444 7254 15456
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 12802 15484 12808 15496
rect 10459 15456 12808 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 13722 15484 13728 15496
rect 13683 15456 13728 15484
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14366 15484 14372 15496
rect 14279 15456 14372 15484
rect 14366 15444 14372 15456
rect 14424 15484 14430 15496
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 14424 15456 16037 15484
rect 14424 15444 14430 15456
rect 16025 15453 16037 15456
rect 16071 15484 16083 15487
rect 16390 15484 16396 15496
rect 16071 15456 16396 15484
rect 16071 15453 16083 15456
rect 16025 15447 16083 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 7561 15419 7619 15425
rect 7561 15416 7573 15419
rect 4126 15388 7573 15416
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 2038 15348 2044 15360
rect 1995 15320 2044 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 2038 15308 2044 15320
rect 2096 15308 2102 15360
rect 2314 15348 2320 15360
rect 2275 15320 2320 15348
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 2958 15308 2964 15360
rect 3016 15348 3022 15360
rect 4126 15348 4154 15388
rect 7561 15385 7573 15388
rect 7607 15385 7619 15419
rect 7561 15379 7619 15385
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9272 15388 9858 15416
rect 9272 15376 9278 15388
rect 3016 15320 4154 15348
rect 3016 15308 3022 15320
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 5813 15351 5871 15357
rect 5813 15348 5825 15351
rect 4764 15320 5825 15348
rect 4764 15308 4770 15320
rect 5813 15317 5825 15320
rect 5859 15317 5871 15351
rect 5813 15311 5871 15317
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 7374 15348 7380 15360
rect 6328 15320 7380 15348
rect 6328 15308 6334 15320
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 9830 15357 9858 15388
rect 9815 15351 9873 15357
rect 9815 15317 9827 15351
rect 9861 15317 9873 15351
rect 9815 15311 9873 15317
rect 9953 15351 10011 15357
rect 9953 15317 9965 15351
rect 9999 15348 10011 15351
rect 10134 15348 10140 15360
rect 9999 15320 10140 15348
rect 9999 15317 10011 15320
rect 9953 15311 10011 15317
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 11238 15348 11244 15360
rect 11199 15320 11244 15348
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 11885 15351 11943 15357
rect 11885 15348 11897 15351
rect 11756 15320 11897 15348
rect 11756 15308 11762 15320
rect 11885 15317 11897 15320
rect 11931 15317 11943 15351
rect 11885 15311 11943 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 2498 15104 2504 15156
rect 2556 15104 2562 15156
rect 3418 15104 3424 15156
rect 3476 15144 3482 15156
rect 5629 15147 5687 15153
rect 3476 15116 4476 15144
rect 3476 15104 3482 15116
rect 2133 15079 2191 15085
rect 2133 15045 2145 15079
rect 2179 15076 2191 15079
rect 2516 15076 2544 15104
rect 4338 15076 4344 15088
rect 2179 15048 4344 15076
rect 2179 15045 2191 15048
rect 2133 15039 2191 15045
rect 4338 15036 4344 15048
rect 4396 15036 4402 15088
rect 106 14968 112 15020
rect 164 15008 170 15020
rect 1578 15008 1584 15020
rect 164 14980 1584 15008
rect 164 14968 170 14980
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 15008 2559 15011
rect 2590 15008 2596 15020
rect 2547 14980 2596 15008
rect 2547 14977 2559 14980
rect 2501 14971 2559 14977
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 4448 15008 4476 15116
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 5994 15144 6000 15156
rect 5675 15116 6000 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 6236 15116 6653 15144
rect 6236 15104 6242 15116
rect 6641 15113 6653 15116
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7929 15147 7987 15153
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 8202 15144 8208 15156
rect 7975 15116 8208 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8343 15116 9076 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 5261 15079 5319 15085
rect 5261 15045 5273 15079
rect 5307 15076 5319 15079
rect 6196 15076 6224 15104
rect 5307 15048 6224 15076
rect 8220 15076 8248 15104
rect 9048 15085 9076 15116
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 9456 15116 10517 15144
rect 9456 15104 9462 15116
rect 10505 15113 10517 15116
rect 10551 15144 10563 15147
rect 12434 15144 12440 15156
rect 10551 15116 12440 15144
rect 10551 15113 10563 15116
rect 10505 15107 10563 15113
rect 12434 15104 12440 15116
rect 12492 15104 12498 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 13969 15116 16313 15144
rect 8895 15079 8953 15085
rect 8895 15076 8907 15079
rect 8220 15048 8907 15076
rect 5307 15045 5319 15048
rect 5261 15039 5319 15045
rect 8895 15045 8907 15048
rect 8941 15045 8953 15079
rect 8895 15039 8953 15045
rect 9033 15079 9091 15085
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 10134 15076 10140 15088
rect 9079 15048 10140 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 10778 15036 10784 15088
rect 10836 15076 10842 15088
rect 12161 15079 12219 15085
rect 12161 15076 12173 15079
rect 10836 15048 12173 15076
rect 10836 15036 10842 15048
rect 12161 15045 12173 15048
rect 12207 15045 12219 15079
rect 12161 15039 12219 15045
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 4448 14980 4537 15008
rect 4525 14977 4537 14980
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 8711 14980 9137 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 9125 14977 9137 14980
rect 9171 15008 9183 15011
rect 11422 15008 11428 15020
rect 9171 14980 9674 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 2038 14940 2044 14952
rect 1443 14912 2044 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 2958 14940 2964 14952
rect 2919 14912 2964 14940
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14940 3755 14943
rect 4062 14940 4068 14952
rect 3743 14912 4068 14940
rect 3743 14909 3755 14912
rect 3697 14903 3755 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6380 14912 6837 14940
rect 4080 14872 4108 14900
rect 4249 14875 4307 14881
rect 4249 14872 4261 14875
rect 4080 14844 4261 14872
rect 4249 14841 4261 14844
rect 4295 14841 4307 14875
rect 4249 14835 4307 14841
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14841 4399 14875
rect 4341 14835 4399 14841
rect 4065 14807 4123 14813
rect 4065 14773 4077 14807
rect 4111 14804 4123 14807
rect 4356 14804 4384 14835
rect 4430 14832 4436 14884
rect 4488 14872 4494 14884
rect 5721 14875 5779 14881
rect 5721 14872 5733 14875
rect 4488 14844 5733 14872
rect 4488 14832 4494 14844
rect 5721 14841 5733 14844
rect 5767 14841 5779 14875
rect 5721 14835 5779 14841
rect 6380 14816 6408 14912
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7190 14940 7196 14952
rect 6871 14912 7196 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7374 14940 7380 14952
rect 7335 14912 7380 14940
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 8662 14832 8668 14884
rect 8720 14872 8726 14884
rect 8757 14875 8815 14881
rect 8757 14872 8769 14875
rect 8720 14844 8769 14872
rect 8720 14832 8726 14844
rect 8757 14841 8769 14844
rect 8803 14841 8815 14875
rect 8757 14835 8815 14841
rect 4706 14804 4712 14816
rect 4111 14776 4712 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 6273 14807 6331 14813
rect 6273 14773 6285 14807
rect 6319 14804 6331 14807
rect 6362 14804 6368 14816
rect 6319 14776 6368 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6914 14804 6920 14816
rect 6875 14776 6920 14804
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 9398 14804 9404 14816
rect 9359 14776 9404 14804
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 9646 14804 9674 14980
rect 10704 14980 11428 15008
rect 10704 14949 10732 14980
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 11330 14940 11336 14952
rect 11195 14912 11336 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 10321 14875 10379 14881
rect 10321 14841 10333 14875
rect 10367 14872 10379 14875
rect 11164 14872 11192 14903
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 12176 14940 12204 15039
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13814 15008 13820 15020
rect 13771 14980 13820 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 13814 14968 13820 14980
rect 13872 15008 13878 15020
rect 13969 15008 13997 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 17586 15144 17592 15156
rect 17547 15116 17592 15144
rect 16301 15107 16359 15113
rect 17586 15104 17592 15116
rect 17644 15104 17650 15156
rect 15565 15079 15623 15085
rect 15565 15045 15577 15079
rect 15611 15076 15623 15079
rect 16114 15076 16120 15088
rect 15611 15048 16120 15076
rect 15611 15045 15623 15048
rect 15565 15039 15623 15045
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 13872 14980 13997 15008
rect 14553 15011 14611 15017
rect 13872 14968 13878 14980
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 14642 15008 14648 15020
rect 14599 14980 14648 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 14826 15008 14832 15020
rect 14787 14980 14832 15008
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12176 14912 12449 14940
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12860 14912 12909 14940
rect 12860 14900 12866 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15933 14943 15991 14949
rect 15933 14940 15945 14943
rect 15344 14912 15945 14940
rect 15344 14900 15350 14912
rect 15933 14909 15945 14912
rect 15979 14940 15991 14943
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 15979 14912 16129 14940
rect 15979 14909 15991 14912
rect 15933 14903 15991 14909
rect 16117 14909 16129 14912
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 13170 14872 13176 14884
rect 10367 14844 11192 14872
rect 13131 14844 13176 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 14645 14875 14703 14881
rect 14645 14841 14657 14875
rect 14691 14841 14703 14875
rect 14645 14835 14703 14841
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9646 14776 9873 14804
rect 9861 14773 9873 14776
rect 9907 14804 9919 14807
rect 10042 14804 10048 14816
rect 9907 14776 10048 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10042 14764 10048 14776
rect 10100 14804 10106 14816
rect 10686 14804 10692 14816
rect 10100 14776 10692 14804
rect 10100 14764 10106 14776
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11422 14804 11428 14816
rect 11383 14776 11428 14804
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 11756 14776 11805 14804
rect 11756 14764 11762 14776
rect 11793 14773 11805 14776
rect 11839 14773 11851 14807
rect 11793 14767 11851 14773
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14277 14807 14335 14813
rect 14277 14804 14289 14807
rect 13872 14776 14289 14804
rect 13872 14764 13878 14776
rect 14277 14773 14289 14776
rect 14323 14804 14335 14807
rect 14660 14804 14688 14835
rect 14323 14776 14688 14804
rect 14323 14773 14335 14776
rect 14277 14767 14335 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 4126 14572 7113 14600
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2041 14535 2099 14541
rect 2041 14532 2053 14535
rect 1820 14504 2053 14532
rect 1820 14492 1826 14504
rect 2041 14501 2053 14504
rect 2087 14532 2099 14535
rect 2590 14532 2596 14544
rect 2087 14504 2596 14532
rect 2087 14501 2099 14504
rect 2041 14495 2099 14501
rect 2590 14492 2596 14504
rect 2648 14532 2654 14544
rect 4126 14532 4154 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 7101 14563 7159 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8720 14572 8953 14600
rect 8720 14560 8726 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9272 14572 9321 14600
rect 9272 14560 9278 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 9309 14563 9367 14569
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 9732 14572 10517 14600
rect 9732 14560 9738 14572
rect 10505 14569 10517 14572
rect 10551 14569 10563 14603
rect 10505 14563 10563 14569
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 11333 14603 11391 14609
rect 11333 14600 11345 14603
rect 10836 14572 11345 14600
rect 10836 14560 10842 14572
rect 11333 14569 11345 14572
rect 11379 14600 11391 14603
rect 11422 14600 11428 14612
rect 11379 14572 11428 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12526 14600 12532 14612
rect 12207 14572 12532 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 12860 14572 12909 14600
rect 12860 14560 12866 14572
rect 12897 14569 12909 14572
rect 12943 14569 12955 14603
rect 14642 14600 14648 14612
rect 14603 14572 14648 14600
rect 12897 14563 12955 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 16390 14600 16396 14612
rect 16351 14572 16396 14600
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 5534 14532 5540 14544
rect 2648 14504 4154 14532
rect 5495 14504 5540 14532
rect 2648 14492 2654 14504
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 6546 14541 6552 14544
rect 6543 14532 6552 14541
rect 6459 14504 6552 14532
rect 6543 14495 6552 14504
rect 6604 14532 6610 14544
rect 6822 14532 6828 14544
rect 6604 14504 6828 14532
rect 6546 14492 6552 14495
rect 6604 14492 6610 14504
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 7469 14535 7527 14541
rect 7469 14532 7481 14535
rect 7432 14504 7481 14532
rect 7432 14492 7438 14504
rect 7469 14501 7481 14504
rect 7515 14532 7527 14535
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 7515 14504 7849 14532
rect 7515 14501 7527 14504
rect 7469 14495 7527 14501
rect 7837 14501 7849 14504
rect 7883 14532 7895 14535
rect 7883 14504 8524 14532
rect 7883 14501 7895 14504
rect 7837 14495 7895 14501
rect 4706 14464 4712 14476
rect 4667 14436 4712 14464
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 6181 14467 6239 14473
rect 6181 14464 6193 14467
rect 6144 14436 6193 14464
rect 6144 14424 6150 14436
rect 6181 14433 6193 14436
rect 6227 14464 6239 14467
rect 6914 14464 6920 14476
rect 6227 14436 6920 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14464 8263 14467
rect 8386 14464 8392 14476
rect 8251 14436 8392 14464
rect 8251 14433 8263 14436
rect 8205 14427 8263 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 8496 14473 8524 14504
rect 12342 14492 12348 14544
rect 12400 14532 12406 14544
rect 12820 14532 12848 14560
rect 12400 14504 12848 14532
rect 12400 14492 12406 14504
rect 12986 14492 12992 14544
rect 13044 14532 13050 14544
rect 13630 14532 13636 14544
rect 13044 14504 13636 14532
rect 13044 14492 13050 14504
rect 13630 14492 13636 14504
rect 13688 14532 13694 14544
rect 13770 14535 13828 14541
rect 13770 14532 13782 14535
rect 13688 14504 13782 14532
rect 13688 14492 13694 14504
rect 13770 14501 13782 14504
rect 13816 14501 13828 14535
rect 13770 14495 13828 14501
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 16114 14532 16120 14544
rect 15611 14504 16120 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9398 14464 9404 14476
rect 8527 14436 9404 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9640 14436 9689 14464
rect 9640 14424 9646 14436
rect 9677 14433 9689 14436
rect 9723 14464 9735 14467
rect 9950 14464 9956 14476
rect 9723 14436 9956 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10134 14424 10140 14476
rect 10192 14464 10198 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 10192 14436 10241 14464
rect 10192 14424 10198 14436
rect 10229 14433 10241 14436
rect 10275 14464 10287 14467
rect 10870 14464 10876 14476
rect 10275 14436 10876 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11514 14464 11520 14476
rect 11475 14436 11520 14464
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 12434 14464 12440 14476
rect 12395 14436 12440 14464
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13446 14464 13452 14476
rect 13228 14436 13452 14464
rect 13228 14424 13234 14436
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 16942 14464 16948 14476
rect 16903 14436 16948 14464
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2406 14396 2412 14408
rect 2367 14368 2412 14396
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 3292 14368 4077 14396
rect 3292 14356 3298 14368
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 8404 14396 8432 14424
rect 11698 14396 11704 14408
rect 8404 14368 11704 14396
rect 4065 14359 4123 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 3786 14288 3792 14340
rect 3844 14328 3850 14340
rect 5534 14328 5540 14340
rect 3844 14300 5540 14328
rect 3844 14288 3850 14300
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 8938 14288 8944 14340
rect 8996 14328 9002 14340
rect 9214 14328 9220 14340
rect 8996 14300 9220 14328
rect 8996 14288 9002 14300
rect 9214 14288 9220 14300
rect 9272 14328 9278 14340
rect 9272 14300 10272 14328
rect 9272 14288 9278 14300
rect 3142 14220 3148 14272
rect 3200 14260 3206 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 3200 14232 3249 14260
rect 3200 14220 3206 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 5258 14260 5264 14272
rect 5219 14232 5264 14260
rect 3237 14223 3295 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5442 14220 5448 14272
rect 5500 14260 5506 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 5500 14232 9873 14260
rect 5500 14220 5506 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 10244 14260 10272 14300
rect 11422 14288 11428 14340
rect 11480 14328 11486 14340
rect 11606 14328 11612 14340
rect 11480 14300 11612 14328
rect 11480 14288 11486 14300
rect 11606 14288 11612 14300
rect 11664 14288 11670 14340
rect 11882 14288 11888 14340
rect 11940 14328 11946 14340
rect 13265 14331 13323 14337
rect 13265 14328 13277 14331
rect 11940 14300 13277 14328
rect 11940 14288 11946 14300
rect 13265 14297 13277 14300
rect 13311 14328 13323 14331
rect 13722 14328 13728 14340
rect 13311 14300 13728 14328
rect 13311 14297 13323 14300
rect 13265 14291 13323 14297
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 17083 14331 17141 14337
rect 17083 14297 17095 14331
rect 17129 14328 17141 14331
rect 21358 14328 21364 14340
rect 17129 14300 21364 14328
rect 17129 14297 17141 14300
rect 17083 14291 17141 14297
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 10594 14260 10600 14272
rect 10244 14232 10600 14260
rect 9861 14223 9919 14229
rect 10594 14220 10600 14232
rect 10652 14260 10658 14272
rect 11974 14260 11980 14272
rect 10652 14232 11980 14260
rect 10652 14220 10658 14232
rect 11974 14220 11980 14232
rect 12032 14260 12038 14272
rect 12621 14263 12679 14269
rect 12621 14260 12633 14263
rect 12032 14232 12633 14260
rect 12032 14220 12038 14232
rect 12621 14229 12633 14232
rect 12667 14229 12679 14263
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 12621 14223 12679 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4706 14056 4712 14068
rect 4203 14028 4712 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 10873 14059 10931 14065
rect 10873 14056 10885 14059
rect 6696 14028 10885 14056
rect 6696 14016 6702 14028
rect 10873 14025 10885 14028
rect 10919 14025 10931 14059
rect 10873 14019 10931 14025
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 11974 14056 11980 14068
rect 11931 14028 11980 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12434 14056 12440 14068
rect 12299 14028 12440 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14553 14059 14611 14065
rect 14553 14056 14565 14059
rect 14424 14028 14565 14056
rect 14424 14016 14430 14028
rect 14553 14025 14565 14028
rect 14599 14056 14611 14059
rect 15378 14056 15384 14068
rect 14599 14028 15384 14056
rect 14599 14025 14611 14028
rect 14553 14019 14611 14025
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 3326 13948 3332 14000
rect 3384 13988 3390 14000
rect 7745 13991 7803 13997
rect 7745 13988 7757 13991
rect 3384 13960 7757 13988
rect 3384 13948 3390 13960
rect 7745 13957 7757 13960
rect 7791 13957 7803 13991
rect 7745 13951 7803 13957
rect 8938 13948 8944 14000
rect 8996 13997 9002 14000
rect 8996 13991 9045 13997
rect 8996 13957 8999 13991
rect 9033 13957 9045 13991
rect 9122 13988 9128 14000
rect 9083 13960 9128 13988
rect 8996 13951 9045 13957
rect 8996 13948 9002 13951
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 9950 13988 9956 14000
rect 9911 13960 9956 13988
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 10594 13997 10600 14000
rect 10578 13991 10600 13997
rect 10578 13957 10590 13991
rect 10578 13951 10600 13957
rect 10594 13948 10600 13951
rect 10652 13948 10658 14000
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 10962 13988 10968 14000
rect 10735 13960 10968 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1452 13892 1593 13920
rect 1452 13880 1458 13892
rect 1581 13889 1593 13892
rect 1627 13920 1639 13923
rect 2501 13923 2559 13929
rect 2501 13920 2513 13923
rect 1627 13892 2513 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 2501 13889 2513 13892
rect 2547 13889 2559 13923
rect 3418 13920 3424 13932
rect 3379 13892 3424 13920
rect 2501 13883 2559 13889
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 7374 13920 7380 13932
rect 5184 13892 7380 13920
rect 5184 13861 5212 13892
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 9214 13920 9220 13932
rect 8803 13892 9220 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9674 13880 9680 13932
rect 9732 13880 9738 13932
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5169 13855 5227 13861
rect 5169 13852 5181 13855
rect 5123 13824 5181 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5169 13821 5181 13824
rect 5215 13821 5227 13855
rect 5169 13815 5227 13821
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5316 13824 5641 13852
rect 5316 13812 5322 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 6822 13852 6828 13864
rect 5675 13824 5764 13852
rect 6783 13824 6828 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 1670 13784 1676 13796
rect 1631 13756 1676 13784
rect 1670 13744 1676 13756
rect 1728 13744 1734 13796
rect 2225 13787 2283 13793
rect 2225 13753 2237 13787
rect 2271 13784 2283 13787
rect 2406 13784 2412 13796
rect 2271 13756 2412 13784
rect 2271 13753 2283 13756
rect 2225 13747 2283 13753
rect 2406 13744 2412 13756
rect 2464 13744 2470 13796
rect 3142 13784 3148 13796
rect 2792 13756 3148 13784
rect 1302 13676 1308 13728
rect 1360 13716 1366 13728
rect 2792 13716 2820 13756
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 3234 13744 3240 13796
rect 3292 13784 3298 13796
rect 5736 13784 5764 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13852 8447 13855
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8435 13824 8861 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8849 13821 8861 13824
rect 8895 13852 8907 13855
rect 9692 13852 9720 13880
rect 8895 13824 9720 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 10100 13824 10425 13852
rect 10100 13812 10106 13824
rect 10413 13821 10425 13824
rect 10459 13821 10471 13855
rect 10413 13815 10471 13821
rect 6638 13784 6644 13796
rect 3292 13756 3337 13784
rect 5736 13756 6644 13784
rect 3292 13744 3298 13756
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 7146 13787 7204 13793
rect 7146 13784 7158 13787
rect 6748 13756 7158 13784
rect 1360 13688 2820 13716
rect 2961 13719 3019 13725
rect 1360 13676 1366 13688
rect 2961 13685 2973 13719
rect 3007 13716 3019 13719
rect 3252 13716 3280 13744
rect 5442 13716 5448 13728
rect 3007 13688 3280 13716
rect 5403 13688 5448 13716
rect 3007 13685 3019 13688
rect 2961 13679 3019 13685
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 6052 13688 6193 13716
rect 6052 13676 6058 13688
rect 6181 13685 6193 13688
rect 6227 13716 6239 13719
rect 6546 13716 6552 13728
rect 6227 13688 6552 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6546 13676 6552 13688
rect 6604 13716 6610 13728
rect 6748 13716 6776 13756
rect 7146 13753 7158 13756
rect 7192 13753 7204 13787
rect 7146 13747 7204 13753
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 10704 13784 10732 13951
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 15746 13988 15752 14000
rect 15707 13960 15752 13988
rect 15746 13948 15752 13960
rect 15804 13988 15810 14000
rect 16942 13988 16948 14000
rect 15804 13960 16948 13988
rect 15804 13948 15810 13960
rect 16942 13948 16948 13960
rect 17000 13988 17006 14000
rect 17129 13991 17187 13997
rect 17129 13988 17141 13991
rect 17000 13960 17141 13988
rect 17000 13948 17006 13960
rect 17129 13957 17141 13960
rect 17175 13957 17187 13991
rect 17129 13951 17187 13957
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15470 13920 15476 13932
rect 15059 13892 15476 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 9180 13756 10732 13784
rect 9180 13744 9186 13756
rect 6604 13688 6776 13716
rect 6604 13676 6610 13688
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7282 13716 7288 13728
rect 6880 13688 7288 13716
rect 6880 13676 6886 13688
rect 7282 13676 7288 13688
rect 7340 13716 7346 13728
rect 8018 13716 8024 13728
rect 7340 13688 8024 13716
rect 7340 13676 7346 13688
rect 8018 13676 8024 13688
rect 8076 13676 8082 13728
rect 9490 13716 9496 13728
rect 9451 13688 9496 13716
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 10321 13719 10379 13725
rect 10321 13685 10333 13719
rect 10367 13716 10379 13719
rect 10796 13716 10824 13883
rect 15470 13880 15476 13892
rect 15528 13920 15534 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15528 13892 16681 13920
rect 15528 13880 15534 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 11606 13784 11612 13796
rect 11256 13756 11612 13784
rect 11256 13716 11284 13756
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 12713 13787 12771 13793
rect 12713 13753 12725 13787
rect 12759 13784 12771 13787
rect 13167 13787 13225 13793
rect 13167 13784 13179 13787
rect 12759 13756 13179 13784
rect 12759 13753 12771 13756
rect 12713 13747 12771 13753
rect 13167 13753 13179 13756
rect 13213 13784 13225 13787
rect 13630 13784 13636 13796
rect 13213 13756 13636 13784
rect 13213 13753 13225 13756
rect 13167 13747 13225 13753
rect 13630 13744 13636 13756
rect 13688 13784 13694 13796
rect 14001 13787 14059 13793
rect 14001 13784 14013 13787
rect 13688 13756 14013 13784
rect 13688 13744 13694 13756
rect 14001 13753 14013 13756
rect 14047 13753 14059 13787
rect 15194 13784 15200 13796
rect 15155 13756 15200 13784
rect 14001 13747 14059 13753
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 15289 13787 15347 13793
rect 15289 13753 15301 13787
rect 15335 13784 15347 13787
rect 15378 13784 15384 13796
rect 15335 13756 15384 13784
rect 15335 13753 15347 13756
rect 15289 13747 15347 13753
rect 15378 13744 15384 13756
rect 15436 13744 15442 13796
rect 16485 13787 16543 13793
rect 16485 13784 16497 13787
rect 15948 13756 16497 13784
rect 11514 13716 11520 13728
rect 10367 13688 11284 13716
rect 11475 13688 11520 13716
rect 10367 13685 10379 13688
rect 10321 13679 10379 13685
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 13725 13719 13783 13725
rect 13725 13685 13737 13719
rect 13771 13716 13783 13719
rect 13814 13716 13820 13728
rect 13771 13688 13820 13716
rect 13771 13685 13783 13688
rect 13725 13679 13783 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 15212 13716 15240 13744
rect 15948 13716 15976 13756
rect 16485 13753 16497 13756
rect 16531 13753 16543 13787
rect 16485 13747 16543 13753
rect 16114 13716 16120 13728
rect 15212 13688 15976 13716
rect 16075 13688 16120 13716
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2590 13512 2596 13524
rect 2551 13484 2596 13512
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6236 13484 6285 13512
rect 6236 13472 6242 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 6273 13475 6331 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 9122 13512 9128 13524
rect 9083 13484 9128 13512
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9858 13512 9864 13524
rect 9272 13484 9864 13512
rect 9272 13472 9278 13484
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10008 13484 10701 13512
rect 10008 13472 10014 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 11020 13484 11161 13512
rect 11020 13472 11026 13484
rect 11149 13481 11161 13484
rect 11195 13481 11207 13515
rect 13446 13512 13452 13524
rect 13407 13484 13452 13512
rect 11149 13475 11207 13481
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13444 1823 13447
rect 3326 13444 3332 13456
rect 1811 13416 3332 13444
rect 1811 13413 1823 13416
rect 1765 13407 1823 13413
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 4430 13444 4436 13456
rect 4391 13416 4436 13444
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 6472 13416 8156 13444
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 6472 13385 6500 13416
rect 8128 13388 8156 13416
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 9456 13416 10425 13444
rect 9456 13404 9462 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 12621 13447 12679 13453
rect 12621 13413 12633 13447
rect 12667 13444 12679 13447
rect 12802 13444 12808 13456
rect 12667 13416 12808 13444
rect 12667 13413 12679 13416
rect 12621 13407 12679 13413
rect 12802 13404 12808 13416
rect 12860 13444 12866 13456
rect 12897 13447 12955 13453
rect 12897 13444 12909 13447
rect 12860 13416 12909 13444
rect 12860 13404 12866 13416
rect 12897 13413 12909 13416
rect 12943 13413 12955 13447
rect 12897 13407 12955 13413
rect 13722 13404 13728 13456
rect 13780 13444 13786 13456
rect 13817 13447 13875 13453
rect 13817 13444 13829 13447
rect 13780 13416 13829 13444
rect 13780 13404 13786 13416
rect 13817 13413 13829 13416
rect 13863 13413 13875 13447
rect 13817 13407 13875 13413
rect 14369 13447 14427 13453
rect 14369 13413 14381 13447
rect 14415 13444 14427 13447
rect 14826 13444 14832 13456
rect 14415 13416 14832 13444
rect 14415 13413 14427 13416
rect 14369 13407 14427 13413
rect 14826 13404 14832 13416
rect 14884 13444 14890 13456
rect 15194 13444 15200 13456
rect 14884 13416 15200 13444
rect 14884 13404 14890 13416
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 16025 13447 16083 13453
rect 16025 13413 16037 13447
rect 16071 13444 16083 13447
rect 16114 13444 16120 13456
rect 16071 13416 16120 13444
rect 16071 13413 16083 13416
rect 16025 13407 16083 13413
rect 16114 13404 16120 13416
rect 16172 13404 16178 13456
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 6420 13348 6469 13376
rect 6420 13336 6426 13348
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6638 13376 6644 13388
rect 6599 13348 6644 13376
rect 6457 13339 6515 13345
rect 6638 13336 6644 13348
rect 6696 13336 6702 13388
rect 8110 13376 8116 13388
rect 8071 13348 8116 13376
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8570 13376 8576 13388
rect 8483 13348 8576 13376
rect 8570 13336 8576 13348
rect 8628 13376 8634 13388
rect 9490 13376 9496 13388
rect 8628 13348 9496 13376
rect 8628 13336 8634 13348
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9950 13376 9956 13388
rect 9911 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 11885 13379 11943 13385
rect 11885 13376 11897 13379
rect 11756 13348 11897 13376
rect 11756 13336 11762 13348
rect 11885 13345 11897 13348
rect 11931 13345 11943 13379
rect 12342 13376 12348 13388
rect 12303 13348 12348 13376
rect 11885 13339 11943 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 15378 13376 15384 13388
rect 15339 13348 15384 13376
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 1946 13308 1952 13320
rect 1907 13280 1952 13308
rect 1946 13268 1952 13280
rect 2004 13308 2010 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2004 13280 2973 13308
rect 2004 13268 2010 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 4338 13308 4344 13320
rect 4299 13280 4344 13308
rect 2961 13271 3019 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4614 13308 4620 13320
rect 4575 13280 4620 13308
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13596 13280 13737 13308
rect 13596 13268 13602 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 8352 13212 8984 13240
rect 8352 13200 8358 13212
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 4246 13172 4252 13184
rect 1820 13144 4252 13172
rect 1820 13132 1826 13144
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7374 13172 7380 13184
rect 6972 13144 7380 13172
rect 6972 13132 6978 13144
rect 7374 13132 7380 13144
rect 7432 13172 7438 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7432 13144 7849 13172
rect 7432 13132 7438 13144
rect 7837 13141 7849 13144
rect 7883 13172 7895 13175
rect 8386 13172 8392 13184
rect 7883 13144 8392 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 8956 13172 8984 13212
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 11054 13240 11060 13252
rect 9088 13212 11060 13240
rect 9088 13200 9094 13212
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 9401 13175 9459 13181
rect 9401 13172 9413 13175
rect 8956 13144 9413 13172
rect 9401 13141 9413 13144
rect 9447 13141 9459 13175
rect 9401 13135 9459 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2590 12968 2596 12980
rect 2503 12940 2596 12968
rect 2590 12928 2596 12940
rect 2648 12968 2654 12980
rect 3326 12968 3332 12980
rect 2648 12940 3332 12968
rect 2648 12928 2654 12940
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 6362 12968 6368 12980
rect 6319 12940 6368 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 10873 12971 10931 12977
rect 10873 12937 10885 12971
rect 10919 12968 10931 12971
rect 10962 12968 10968 12980
rect 10919 12940 10968 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 11238 12968 11244 12980
rect 11199 12940 11244 12968
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11756 12940 11989 12968
rect 11756 12928 11762 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13722 12968 13728 12980
rect 13679 12940 13728 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 1596 12872 3004 12900
rect 1596 12841 1624 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1946 12832 1952 12844
rect 1907 12804 1952 12832
rect 1581 12795 1639 12801
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2976 12841 3004 12872
rect 3050 12860 3056 12912
rect 3108 12900 3114 12912
rect 4430 12900 4436 12912
rect 3108 12872 4436 12900
rect 3108 12860 3114 12872
rect 4430 12860 4436 12872
rect 4488 12900 4494 12912
rect 4525 12903 4583 12909
rect 4525 12900 4537 12903
rect 4488 12872 4537 12900
rect 4488 12860 4494 12872
rect 4525 12869 4537 12872
rect 4571 12900 4583 12903
rect 5905 12903 5963 12909
rect 5905 12900 5917 12903
rect 4571 12872 5917 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 5905 12869 5917 12872
rect 5951 12869 5963 12903
rect 10980 12900 11008 12928
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 10980 12872 12633 12900
rect 5905 12863 5963 12869
rect 12621 12869 12633 12872
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3970 12832 3976 12844
rect 3007 12804 3976 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 4154 12832 4160 12844
rect 4067 12804 4160 12832
rect 4154 12792 4160 12804
rect 4212 12832 4218 12844
rect 4614 12832 4620 12844
rect 4212 12804 4620 12832
rect 4212 12792 4218 12804
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5074 12832 5080 12844
rect 5031 12804 5080 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5074 12792 5080 12804
rect 5132 12832 5138 12844
rect 6178 12832 6184 12844
rect 5132 12804 6184 12832
rect 5132 12792 5138 12804
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 8662 12832 8668 12844
rect 6687 12804 7696 12832
rect 8623 12804 8668 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7668 12773 7696 12804
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12832 11023 12835
rect 11422 12832 11428 12844
rect 11011 12804 11428 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 11422 12792 11428 12804
rect 11480 12832 11486 12844
rect 13740 12841 13768 12928
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 11480 12804 11621 12832
rect 11480 12792 11486 12804
rect 11609 12801 11621 12804
rect 11655 12801 11667 12835
rect 11609 12795 11667 12801
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 6972 12736 7113 12764
rect 6972 12724 6978 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 7742 12764 7748 12776
rect 7699 12736 7748 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7742 12724 7748 12736
rect 7800 12764 7806 12776
rect 8570 12764 8576 12776
rect 7800 12736 8576 12764
rect 7800 12724 7806 12736
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9585 12767 9643 12773
rect 8812 12736 9168 12764
rect 8812 12724 8818 12736
rect 1673 12699 1731 12705
rect 1673 12665 1685 12699
rect 1719 12696 1731 12699
rect 1946 12696 1952 12708
rect 1719 12668 1952 12696
rect 1719 12665 1731 12668
rect 1673 12659 1731 12665
rect 1946 12656 1952 12668
rect 2004 12656 2010 12708
rect 3510 12696 3516 12708
rect 3471 12668 3516 12696
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 3605 12699 3663 12705
rect 3605 12665 3617 12699
rect 3651 12665 3663 12699
rect 7834 12696 7840 12708
rect 7795 12668 7840 12696
rect 3605 12659 3663 12665
rect 3234 12628 3240 12640
rect 3195 12600 3240 12628
rect 3234 12588 3240 12600
rect 3292 12628 3298 12640
rect 3620 12628 3648 12659
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 8986 12699 9044 12705
rect 8986 12696 8998 12699
rect 8496 12668 8998 12696
rect 3292 12600 3648 12628
rect 4893 12631 4951 12637
rect 3292 12588 3298 12600
rect 4893 12597 4905 12631
rect 4939 12628 4951 12631
rect 5350 12628 5356 12640
rect 4939 12600 5356 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8496 12637 8524 12668
rect 8986 12665 8998 12668
rect 9032 12665 9044 12699
rect 9140 12696 9168 12736
rect 9585 12733 9597 12767
rect 9631 12764 9643 12767
rect 9858 12764 9864 12776
rect 9631 12736 9864 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10744 12767 10802 12773
rect 10744 12733 10756 12767
rect 10790 12733 10802 12767
rect 10744 12727 10802 12733
rect 10134 12696 10140 12708
rect 9140 12668 10140 12696
rect 8986 12659 9044 12665
rect 10134 12656 10140 12668
rect 10192 12696 10198 12708
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10192 12668 10609 12696
rect 10192 12656 10198 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 7984 12600 8493 12628
rect 7984 12588 7990 12600
rect 8481 12597 8493 12600
rect 8527 12597 8539 12631
rect 9950 12628 9956 12640
rect 9911 12600 9956 12628
rect 8481 12591 8539 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 10759 12628 10787 12727
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12124 12736 12449 12764
rect 12124 12724 12130 12736
rect 12437 12733 12449 12736
rect 12483 12764 12495 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12483 12736 12909 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 13872 12736 13917 12764
rect 13872 12724 13878 12736
rect 11146 12628 11152 12640
rect 10551 12600 11152 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 11146 12588 11152 12600
rect 11204 12628 11210 12640
rect 13078 12628 13084 12640
rect 11204 12600 13084 12628
rect 11204 12588 11210 12600
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 2225 12427 2283 12433
rect 2225 12424 2237 12427
rect 1728 12396 2237 12424
rect 1728 12384 1734 12396
rect 2225 12393 2237 12396
rect 2271 12393 2283 12427
rect 3510 12424 3516 12436
rect 3471 12396 3516 12424
rect 2225 12387 2283 12393
rect 3510 12384 3516 12396
rect 3568 12424 3574 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3568 12396 4077 12424
rect 3568 12384 3574 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 4065 12387 4123 12393
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 4396 12396 4537 12424
rect 4396 12384 4402 12396
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 5074 12424 5080 12436
rect 5035 12396 5080 12424
rect 4525 12387 4583 12393
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 6638 12424 6644 12436
rect 6599 12396 6644 12424
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 7742 12424 7748 12436
rect 7703 12396 7748 12424
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8720 12396 9045 12424
rect 8720 12384 8726 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9033 12387 9091 12393
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11057 12427 11115 12433
rect 11057 12424 11069 12427
rect 11020 12396 11069 12424
rect 11020 12384 11026 12396
rect 11057 12393 11069 12396
rect 11103 12393 11115 12427
rect 11057 12387 11115 12393
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 11885 12427 11943 12433
rect 11885 12424 11897 12427
rect 11848 12396 11897 12424
rect 11848 12384 11854 12396
rect 11885 12393 11897 12396
rect 11931 12393 11943 12427
rect 12342 12424 12348 12436
rect 12303 12396 12348 12424
rect 11885 12387 11943 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 13078 12424 13084 12436
rect 13039 12396 13084 12424
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 13872 12396 13917 12424
rect 13872 12384 13878 12396
rect 3145 12359 3203 12365
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 3234 12356 3240 12368
rect 3191 12328 3240 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 3234 12316 3240 12328
rect 3292 12316 3298 12368
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 5807 12359 5865 12365
rect 5807 12356 5819 12359
rect 5408 12328 5819 12356
rect 5408 12316 5414 12328
rect 5807 12325 5819 12328
rect 5853 12356 5865 12359
rect 5994 12356 6000 12368
rect 5853 12328 6000 12356
rect 5853 12325 5865 12328
rect 5807 12319 5865 12325
rect 5994 12316 6000 12328
rect 6052 12356 6058 12368
rect 6178 12356 6184 12368
rect 6052 12328 6184 12356
rect 6052 12316 6058 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 8158 12359 8216 12365
rect 8158 12356 8170 12359
rect 7984 12328 8170 12356
rect 7984 12316 7990 12328
rect 8158 12325 8170 12328
rect 8204 12325 8216 12359
rect 8158 12319 8216 12325
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9824 12328 9873 12356
rect 9824 12316 9830 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 10778 12316 10784 12368
rect 10836 12356 10842 12368
rect 11241 12359 11299 12365
rect 11241 12356 11253 12359
rect 10836 12328 11253 12356
rect 10836 12316 10842 12328
rect 11241 12325 11253 12328
rect 11287 12325 11299 12359
rect 11241 12319 11299 12325
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12805 12359 12863 12365
rect 12805 12356 12817 12359
rect 11572 12328 12817 12356
rect 11572 12316 11578 12328
rect 12805 12325 12817 12328
rect 12851 12356 12863 12359
rect 13262 12356 13268 12368
rect 12851 12328 13268 12356
rect 12851 12325 12863 12328
rect 12805 12319 12863 12325
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 3050 12288 3056 12300
rect 3011 12260 3056 12288
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 5442 12288 5448 12300
rect 5403 12260 5448 12288
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 7834 12288 7840 12300
rect 7795 12260 7840 12288
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 12986 12288 12992 12300
rect 12947 12260 12992 12288
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9640 12192 9781 12220
rect 9640 12180 9646 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 10042 12220 10048 12232
rect 10003 12192 10048 12220
rect 9769 12183 9827 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11606 12220 11612 12232
rect 11020 12192 11612 12220
rect 11020 12180 11026 12192
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 8536 12124 9413 12152
rect 8536 12112 8542 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 10980 12152 11008 12180
rect 10008 12124 11008 12152
rect 10008 12112 10014 12124
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 13538 12152 13544 12164
rect 11204 12124 13544 12152
rect 11204 12112 11210 12124
rect 13538 12112 13544 12124
rect 13596 12152 13602 12164
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 13596 12124 14105 12152
rect 13596 12112 13602 12124
rect 14093 12121 14105 12124
rect 14139 12121 14151 12155
rect 14093 12115 14151 12121
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 6362 12084 6368 12096
rect 6323 12056 6368 12084
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 6972 12056 7113 12084
rect 6972 12044 6978 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 8754 12084 8760 12096
rect 8715 12056 8760 12084
rect 7101 12047 7159 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10134 12084 10140 12096
rect 9824 12056 10140 12084
rect 9824 12044 9830 12056
rect 10134 12044 10140 12056
rect 10192 12084 10198 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10192 12056 10701 12084
rect 10192 12044 10198 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 11330 12044 11336 12096
rect 11388 12093 11394 12096
rect 11388 12087 11437 12093
rect 11388 12053 11391 12087
rect 11425 12053 11437 12087
rect 11514 12084 11520 12096
rect 11475 12056 11520 12084
rect 11388 12047 11437 12053
rect 11388 12044 11394 12047
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1946 11880 1952 11892
rect 1907 11852 1952 11880
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 3050 11880 3056 11892
rect 2639 11852 3056 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 6178 11880 6184 11892
rect 6091 11852 6184 11880
rect 6178 11840 6184 11852
rect 6236 11880 6242 11892
rect 7926 11880 7932 11892
rect 6236 11852 7932 11880
rect 6236 11840 6242 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 10778 11880 10784 11892
rect 10739 11852 10784 11880
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 10928 11852 11437 11880
rect 10928 11840 10934 11852
rect 11425 11849 11437 11852
rect 11471 11849 11483 11883
rect 11425 11843 11483 11849
rect 9125 11815 9183 11821
rect 9125 11812 9137 11815
rect 8173 11784 9137 11812
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3476 11716 3617 11744
rect 3476 11704 3482 11716
rect 3605 11713 3617 11716
rect 3651 11713 3663 11747
rect 3605 11707 3663 11713
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4338 11744 4344 11756
rect 4295 11716 4344 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4338 11704 4344 11716
rect 4396 11744 4402 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 4396 11716 5457 11744
rect 4396 11704 4402 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 8173 11744 8201 11784
rect 9125 11781 9137 11784
rect 9171 11812 9183 11815
rect 9582 11812 9588 11824
rect 9171 11784 9588 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 12805 11815 12863 11821
rect 12805 11812 12817 11815
rect 11388 11784 12817 11812
rect 11388 11772 11394 11784
rect 12805 11781 12817 11784
rect 12851 11812 12863 11815
rect 12986 11812 12992 11824
rect 12851 11784 12992 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 12986 11772 12992 11784
rect 13044 11772 13050 11824
rect 8478 11744 8484 11756
rect 7147 11716 8201 11744
rect 8439 11716 8484 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 8478 11704 8484 11716
rect 8536 11744 8542 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 8536 11716 9781 11744
rect 8536 11704 8542 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 10042 11744 10048 11756
rect 10003 11716 10048 11744
rect 9769 11707 9827 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 1670 11636 1676 11688
rect 1728 11676 1734 11688
rect 2133 11679 2191 11685
rect 2133 11676 2145 11679
rect 1728 11648 2145 11676
rect 1728 11636 1734 11648
rect 2133 11645 2145 11648
rect 2179 11676 2191 11679
rect 2590 11676 2596 11688
rect 2179 11648 2596 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 11112 11648 11253 11676
rect 11112 11636 11118 11648
rect 11241 11645 11253 11648
rect 11287 11676 11299 11679
rect 11514 11676 11520 11688
rect 11287 11648 11520 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 11514 11636 11520 11648
rect 11572 11676 11578 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11572 11648 11713 11676
rect 11572 11636 11578 11648
rect 11701 11645 11713 11648
rect 11747 11676 11759 11679
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11747 11648 12081 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 13004 11676 13032 11772
rect 17954 11676 17960 11688
rect 13004 11648 17960 11676
rect 12069 11639 12127 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 3694 11617 3700 11620
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11608 3479 11611
rect 3690 11608 3700 11617
rect 3467 11580 3700 11608
rect 3467 11577 3479 11580
rect 3421 11571 3479 11577
rect 3690 11571 3700 11580
rect 3694 11568 3700 11571
rect 3752 11568 3758 11620
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 4632 11580 5181 11608
rect 4632 11552 4660 11580
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 5169 11571 5227 11577
rect 5261 11611 5319 11617
rect 5261 11577 5273 11611
rect 5307 11608 5319 11611
rect 6362 11608 6368 11620
rect 5307 11580 6368 11608
rect 5307 11577 5319 11580
rect 5261 11571 5319 11577
rect 4614 11540 4620 11552
rect 4575 11512 4620 11540
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4982 11540 4988 11552
rect 4895 11512 4988 11540
rect 4982 11500 4988 11512
rect 5040 11540 5046 11552
rect 5276 11540 5304 11571
rect 6362 11568 6368 11580
rect 6420 11568 6426 11620
rect 8202 11608 8208 11620
rect 8163 11580 8208 11608
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8297 11611 8355 11617
rect 8297 11577 8309 11611
rect 8343 11608 8355 11611
rect 8662 11608 8668 11620
rect 8343 11580 8668 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 9858 11608 9864 11620
rect 9819 11580 9864 11608
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 5040 11512 5304 11540
rect 9585 11543 9643 11549
rect 5040 11500 5046 11512
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 9674 11540 9680 11552
rect 9631 11512 9680 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 11020 11512 11069 11540
rect 11020 11500 11026 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 11057 11503 11115 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 2774 11336 2780 11348
rect 2731 11308 2780 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6914 11336 6920 11348
rect 6875 11308 6920 11336
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 7742 11336 7748 11348
rect 7699 11308 7748 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8754 11336 8760 11348
rect 8715 11308 8760 11336
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9858 11336 9864 11348
rect 9539 11308 9864 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 3694 11228 3700 11280
rect 3752 11268 3758 11280
rect 4341 11271 4399 11277
rect 4341 11268 4353 11271
rect 3752 11240 4353 11268
rect 3752 11228 3758 11240
rect 4341 11237 4353 11240
rect 4387 11237 4399 11271
rect 4341 11231 4399 11237
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 7929 11271 7987 11277
rect 7929 11268 7941 11271
rect 7892 11240 7941 11268
rect 7892 11228 7898 11240
rect 7929 11237 7941 11240
rect 7975 11237 7987 11271
rect 8478 11268 8484 11280
rect 8439 11240 8484 11268
rect 7929 11231 7987 11237
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 9674 11268 9680 11280
rect 9635 11240 9680 11268
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2832 11172 2881 11200
rect 2832 11160 2838 11172
rect 2869 11169 2881 11172
rect 2915 11200 2927 11203
rect 3326 11200 3332 11212
rect 2915 11172 3332 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 4982 11200 4988 11212
rect 4943 11172 4988 11200
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 9784 11209 9812 11308
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 4890 11132 4896 11144
rect 1728 11104 4896 11132
rect 1728 11092 1734 11104
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7708 11104 7849 11132
rect 7708 11092 7714 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 8202 11064 8208 11076
rect 7331 11036 8208 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 3513 10999 3571 11005
rect 3513 10996 3525 10999
rect 3476 10968 3525 10996
rect 3476 10956 3482 10968
rect 3513 10965 3525 10968
rect 3559 10965 3571 10999
rect 3513 10959 3571 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2639 10795 2697 10801
rect 2639 10792 2651 10795
rect 2372 10764 2651 10792
rect 2372 10752 2378 10764
rect 2639 10761 2651 10764
rect 2685 10761 2697 10795
rect 2639 10755 2697 10761
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4154 10792 4160 10804
rect 4111 10764 4160 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 2038 10684 2044 10736
rect 2096 10724 2102 10736
rect 3651 10727 3709 10733
rect 3651 10724 3663 10727
rect 2096 10696 3663 10724
rect 2096 10684 2102 10696
rect 3651 10693 3663 10696
rect 3697 10693 3709 10727
rect 4080 10724 4108 10755
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4982 10792 4988 10804
rect 4479 10764 4988 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5675 10795 5733 10801
rect 5675 10792 5687 10795
rect 5592 10764 5687 10792
rect 5592 10752 5598 10764
rect 5675 10761 5687 10764
rect 5721 10761 5733 10795
rect 5675 10755 5733 10761
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8812 10764 8861 10792
rect 8812 10752 8818 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 9766 10792 9772 10804
rect 9631 10764 9772 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 9916 10764 10241 10792
rect 9916 10752 9922 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 10686 10792 10692 10804
rect 10643 10764 10692 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 3651 10687 3709 10693
rect 3896 10696 4108 10724
rect 4663 10727 4721 10733
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2774 10656 2780 10668
rect 2363 10628 2780 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1946 10588 1952 10600
rect 1443 10560 1952 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2498 10588 2504 10600
rect 2556 10597 2562 10600
rect 2556 10591 2594 10597
rect 2446 10560 2504 10588
rect 2498 10548 2504 10560
rect 2582 10588 2594 10591
rect 2961 10591 3019 10597
rect 2961 10588 2973 10591
rect 2582 10560 2973 10588
rect 2582 10557 2594 10560
rect 2556 10551 2594 10557
rect 2961 10557 2973 10560
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 3580 10591 3638 10597
rect 3580 10557 3592 10591
rect 3626 10588 3638 10591
rect 3896 10588 3924 10696
rect 4663 10693 4675 10727
rect 4709 10724 4721 10727
rect 7650 10724 7656 10736
rect 4709 10696 7656 10724
rect 4709 10693 4721 10696
rect 4663 10687 4721 10693
rect 7650 10684 7656 10696
rect 7708 10684 7714 10736
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 6730 10656 6736 10668
rect 4212 10628 6736 10656
rect 4212 10616 4218 10628
rect 6730 10616 6736 10628
rect 6788 10656 6794 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6788 10628 7021 10656
rect 6788 10616 6794 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10656 7803 10659
rect 7834 10656 7840 10668
rect 7791 10628 7840 10656
rect 7791 10625 7803 10628
rect 7745 10619 7803 10625
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 3626 10560 3924 10588
rect 4249 10591 4307 10597
rect 3626 10557 3638 10560
rect 3580 10551 3638 10557
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4560 10591 4618 10597
rect 4560 10588 4572 10591
rect 4295 10560 4572 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4560 10557 4572 10560
rect 4606 10588 4618 10591
rect 4985 10591 5043 10597
rect 4985 10588 4997 10591
rect 4606 10560 4997 10588
rect 4606 10557 4618 10560
rect 4560 10551 4618 10557
rect 4985 10557 4997 10560
rect 5031 10557 5043 10591
rect 4985 10551 5043 10557
rect 2556 10548 2562 10551
rect 5166 10548 5172 10600
rect 5224 10588 5230 10600
rect 5572 10591 5630 10597
rect 5572 10588 5584 10591
rect 5224 10560 5584 10588
rect 5224 10548 5230 10560
rect 5572 10557 5584 10560
rect 5618 10588 5630 10591
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 5618 10560 6009 10588
rect 5618 10557 5630 10560
rect 5572 10551 5630 10557
rect 5997 10557 6009 10560
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8754 10588 8760 10600
rect 8527 10560 8760 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9398 10588 9404 10600
rect 9359 10560 9404 10588
rect 9398 10548 9404 10560
rect 9456 10588 9462 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9456 10560 9873 10588
rect 9456 10548 9462 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10962 10588 10968 10600
rect 10459 10560 10968 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 106 10412 112 10464
rect 164 10452 170 10464
rect 10980 10461 11008 10548
rect 4157 10455 4215 10461
rect 4157 10452 4169 10455
rect 164 10424 4169 10452
rect 164 10412 170 10424
rect 4157 10421 4169 10424
rect 4203 10421 4215 10455
rect 4157 10415 4215 10421
rect 10965 10455 11023 10461
rect 10965 10421 10977 10455
rect 11011 10452 11023 10455
rect 15378 10452 15384 10464
rect 11011 10424 15384 10452
rect 11011 10421 11023 10424
rect 10965 10415 11023 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2547 10251 2605 10257
rect 2547 10217 2559 10251
rect 2593 10248 2605 10251
rect 2682 10248 2688 10260
rect 2593 10220 2688 10248
rect 2593 10217 2605 10220
rect 2547 10211 2605 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 4203 10251 4261 10257
rect 4203 10248 4215 10251
rect 3568 10220 4215 10248
rect 3568 10208 3574 10220
rect 4203 10217 4215 10220
rect 4249 10217 4261 10251
rect 4203 10211 4261 10217
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 7708 10220 8585 10248
rect 7708 10208 7714 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 1535 10183 1593 10189
rect 1535 10149 1547 10183
rect 1581 10180 1593 10183
rect 3142 10180 3148 10192
rect 1581 10152 3148 10180
rect 1581 10149 1593 10152
rect 1535 10143 1593 10149
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 1448 10115 1506 10121
rect 1448 10081 1460 10115
rect 1494 10081 1506 10115
rect 1448 10075 1506 10081
rect 1463 10044 1491 10075
rect 2314 10072 2320 10124
rect 2372 10112 2378 10124
rect 2476 10115 2534 10121
rect 2476 10112 2488 10115
rect 2372 10084 2488 10112
rect 2372 10072 2378 10084
rect 2476 10081 2488 10084
rect 2522 10112 2534 10115
rect 2958 10112 2964 10124
rect 2522 10084 2964 10112
rect 2522 10081 2534 10084
rect 2476 10075 2534 10081
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4100 10115 4158 10121
rect 4100 10112 4112 10115
rect 3936 10084 4112 10112
rect 3936 10072 3942 10084
rect 4100 10081 4112 10084
rect 4146 10081 4158 10115
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 4100 10075 4158 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 8076 10084 8125 10112
rect 8076 10072 8082 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 2038 10044 2044 10056
rect 1463 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10044 2102 10056
rect 3050 10044 3056 10056
rect 2096 10016 3056 10044
rect 2096 10004 2102 10016
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8386 10044 8392 10056
rect 7975 10016 8392 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 1946 9908 1952 9920
rect 1907 9880 1952 9908
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 8294 9908 8300 9920
rect 2740 9880 8300 9908
rect 2740 9868 2746 9880
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 1535 9707 1593 9713
rect 1535 9704 1547 9707
rect 1360 9676 1547 9704
rect 1360 9664 1366 9676
rect 1535 9673 1547 9676
rect 1581 9673 1593 9707
rect 2314 9704 2320 9716
rect 2275 9676 2320 9704
rect 1535 9667 1593 9673
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2547 9707 2605 9713
rect 2547 9673 2559 9707
rect 2593 9704 2605 9707
rect 3418 9704 3424 9716
rect 2593 9676 3424 9704
rect 2593 9673 2605 9676
rect 2547 9667 2605 9673
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 3602 9704 3608 9716
rect 3563 9676 3608 9704
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 4157 9707 4215 9713
rect 4157 9704 4169 9707
rect 3936 9676 4169 9704
rect 3936 9664 3942 9676
rect 4157 9673 4169 9676
rect 4203 9673 4215 9707
rect 4157 9667 4215 9673
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 3145 9639 3203 9645
rect 3145 9636 3157 9639
rect 2188 9608 3157 9636
rect 2188 9596 2194 9608
rect 3145 9605 3157 9608
rect 3191 9636 3203 9639
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 3191 9608 3249 9636
rect 3191 9605 3203 9608
rect 3145 9599 3203 9605
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 4571 9639 4629 9645
rect 4571 9636 4583 9639
rect 4028 9608 4583 9636
rect 4028 9596 4034 9608
rect 4571 9605 4583 9608
rect 4617 9605 4629 9639
rect 4571 9599 4629 9605
rect 106 9528 112 9580
rect 164 9568 170 9580
rect 164 9540 4154 9568
rect 164 9528 170 9540
rect 1464 9503 1522 9509
rect 1464 9469 1476 9503
rect 1510 9500 1522 9503
rect 1854 9500 1860 9512
rect 1510 9472 1860 9500
rect 1510 9469 1522 9472
rect 1464 9463 1522 9469
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2476 9503 2534 9509
rect 2476 9469 2488 9503
rect 2522 9500 2534 9503
rect 2866 9500 2872 9512
rect 2522 9472 2872 9500
rect 2522 9469 2534 9472
rect 2476 9463 2534 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3456 9503 3514 9509
rect 3456 9500 3468 9503
rect 3191 9472 3468 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3456 9469 3468 9472
rect 3502 9469 3514 9503
rect 4126 9500 4154 9540
rect 4500 9503 4558 9509
rect 4500 9500 4512 9503
rect 4126 9472 4512 9500
rect 3456 9463 3514 9469
rect 4500 9469 4512 9472
rect 4546 9500 4558 9503
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4546 9472 4905 9500
rect 4546 9469 4558 9472
rect 4500 9463 4558 9469
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 4893 9463 4951 9469
rect 7116 9472 7389 9500
rect 7116 9376 7144 9472
rect 7377 9469 7389 9472
rect 7423 9500 7435 9503
rect 7558 9500 7564 9512
rect 7423 9472 7564 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7742 9364 7748 9376
rect 7703 9336 7748 9364
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 8076 9336 8309 9364
rect 8076 9324 8082 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 8297 9327 8355 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1535 9163 1593 9169
rect 1535 9129 1547 9163
rect 1581 9160 1593 9163
rect 1670 9160 1676 9172
rect 1581 9132 1676 9160
rect 1581 9129 1593 9132
rect 1535 9123 1593 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2547 9163 2605 9169
rect 2547 9160 2559 9163
rect 2004 9132 2559 9160
rect 2004 9120 2010 9132
rect 2547 9129 2559 9132
rect 2593 9129 2605 9163
rect 2547 9123 2605 9129
rect 7742 9052 7748 9104
rect 7800 9092 7806 9104
rect 7837 9095 7895 9101
rect 7837 9092 7849 9095
rect 7800 9064 7849 9092
rect 7800 9052 7806 9064
rect 7837 9061 7849 9064
rect 7883 9061 7895 9095
rect 7837 9055 7895 9061
rect 8389 9095 8447 9101
rect 8389 9061 8401 9095
rect 8435 9092 8447 9095
rect 9398 9092 9404 9104
rect 8435 9064 9404 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 106 8984 112 9036
rect 164 9024 170 9036
rect 1432 9027 1490 9033
rect 1432 9024 1444 9027
rect 164 8996 1444 9024
rect 164 8984 170 8996
rect 1432 8993 1444 8996
rect 1478 9024 1490 9027
rect 1854 9024 1860 9036
rect 1478 8996 1860 9024
rect 1478 8993 1490 8996
rect 1432 8987 1490 8993
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2038 9024 2044 9036
rect 1995 8996 2044 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2476 9027 2534 9033
rect 2476 8993 2488 9027
rect 2522 9024 2534 9027
rect 3234 9024 3240 9036
rect 2522 8996 3240 9024
rect 2522 8993 2534 8996
rect 2476 8987 2534 8993
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 7098 8888 7104 8900
rect 2004 8860 7104 8888
rect 2004 8848 2010 8860
rect 7098 8848 7104 8860
rect 7156 8888 7162 8900
rect 7285 8891 7343 8897
rect 7285 8888 7297 8891
rect 7156 8860 7297 8888
rect 7156 8848 7162 8860
rect 7285 8857 7297 8860
rect 7331 8857 7343 8891
rect 7285 8851 7343 8857
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1854 8616 1860 8628
rect 1815 8588 1860 8616
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 2222 8616 2228 8628
rect 2183 8588 2228 8616
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 3234 8576 3240 8588
rect 3292 8616 3298 8628
rect 3292 8588 4154 8616
rect 3292 8576 3298 8588
rect 1673 8551 1731 8557
rect 1673 8517 1685 8551
rect 1719 8548 1731 8551
rect 1762 8548 1768 8560
rect 1719 8520 1768 8548
rect 1719 8517 1731 8520
rect 1673 8511 1731 8517
rect 1762 8508 1768 8520
rect 1820 8508 1826 8560
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 2869 8551 2927 8557
rect 2869 8548 2881 8551
rect 2464 8520 2881 8548
rect 2464 8508 2470 8520
rect 2869 8517 2881 8520
rect 2915 8517 2927 8551
rect 4126 8548 4154 8588
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7800 8588 8217 8616
rect 7800 8576 7806 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 10042 8548 10048 8560
rect 4126 8520 10048 8548
rect 2869 8511 2927 8517
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 1464 8415 1522 8421
rect 1464 8381 1476 8415
rect 1510 8412 1522 8415
rect 2222 8412 2228 8424
rect 1510 8384 2228 8412
rect 1510 8381 1522 8384
rect 1464 8375 1522 8381
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2441 8412 2447 8424
rect 2402 8384 2447 8412
rect 2441 8372 2447 8384
rect 2499 8372 2505 8424
rect 7929 8279 7987 8285
rect 7929 8245 7941 8279
rect 7975 8276 7987 8279
rect 8018 8276 8024 8288
rect 7975 8248 8024 8276
rect 7975 8245 7987 8248
rect 7929 8239 7987 8245
rect 8018 8236 8024 8248
rect 8076 8276 8082 8288
rect 8478 8276 8484 8288
rect 8076 8248 8484 8276
rect 8076 8236 8082 8248
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 1535 7803 1593 7809
rect 1535 7769 1547 7803
rect 1581 7800 1593 7803
rect 1670 7800 1676 7812
rect 1581 7772 1676 7800
rect 1581 7769 1593 7772
rect 1535 7763 1593 7769
rect 1670 7760 1676 7772
rect 1728 7760 1734 7812
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 106 7488 112 7540
rect 164 7528 170 7540
rect 1394 7528 1400 7540
rect 164 7500 1400 7528
rect 164 7488 170 7500
rect 1394 7488 1400 7500
rect 1452 7528 1458 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1452 7500 1593 7528
rect 1452 7488 1458 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 1535 6783 1593 6789
rect 1535 6749 1547 6783
rect 1581 6780 1593 6783
rect 12526 6780 12532 6792
rect 1581 6752 12532 6780
rect 1581 6749 1593 6752
rect 1535 6743 1593 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 106 6400 112 6452
rect 164 6440 170 6452
rect 1394 6440 1400 6452
rect 164 6412 1400 6440
rect 164 6400 170 6412
rect 1394 6400 1400 6412
rect 1452 6440 1458 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1452 6412 1593 6440
rect 1452 6400 1458 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 106 5720 112 5772
rect 164 5760 170 5772
rect 1394 5760 1400 5772
rect 1452 5769 1458 5772
rect 1452 5763 1490 5769
rect 164 5732 1400 5760
rect 164 5720 170 5732
rect 1394 5720 1400 5732
rect 1478 5729 1490 5763
rect 1452 5723 1490 5729
rect 1452 5720 1458 5723
rect 1535 5695 1593 5701
rect 1535 5661 1547 5695
rect 1581 5692 1593 5695
rect 12894 5692 12900 5704
rect 1581 5664 12900 5692
rect 1581 5661 1593 5664
rect 1535 5655 1593 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 106 4632 112 4684
rect 164 4672 170 4684
rect 1394 4672 1400 4684
rect 1452 4681 1458 4684
rect 1452 4675 1490 4681
rect 164 4644 1400 4672
rect 164 4632 170 4644
rect 1394 4632 1400 4644
rect 1478 4641 1490 4675
rect 1452 4635 1490 4641
rect 1452 4632 1458 4635
rect 1535 4607 1593 4613
rect 1535 4573 1547 4607
rect 1581 4604 1593 4607
rect 13170 4604 13176 4616
rect 1581 4576 13176 4604
rect 1581 4573 1593 4576
rect 1535 4567 1593 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1452 4236 1593 4264
rect 1452 4224 1458 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1581 4227 1639 4233
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 106 3544 112 3596
rect 164 3584 170 3596
rect 1432 3587 1490 3593
rect 1432 3584 1444 3587
rect 164 3556 1444 3584
rect 164 3544 170 3556
rect 1432 3553 1444 3556
rect 1478 3584 1490 3587
rect 2222 3584 2228 3596
rect 1478 3556 2228 3584
rect 1478 3553 1490 3556
rect 1432 3547 1490 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1432 2975 1490 2981
rect 1432 2972 1444 2975
rect 1360 2944 1444 2972
rect 1360 2932 1366 2944
rect 1432 2941 1444 2944
rect 1478 2972 1490 2975
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1478 2944 1869 2972
rect 1478 2941 1490 2944
rect 1432 2935 1490 2941
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1535 2839 1593 2845
rect 1535 2836 1547 2839
rect 1452 2808 1547 2836
rect 1452 2796 1458 2808
rect 1535 2805 1547 2808
rect 1581 2805 1593 2839
rect 1535 2799 1593 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2547 2635 2605 2641
rect 2547 2601 2559 2635
rect 2593 2632 2605 2635
rect 6270 2632 6276 2644
rect 2593 2604 6276 2632
rect 2593 2601 2605 2604
rect 2547 2595 2605 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 1432 2499 1490 2505
rect 1432 2496 1444 2499
rect 1268 2468 1444 2496
rect 1268 2456 1274 2468
rect 1432 2465 1444 2468
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1432 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 2130 2456 2136 2508
rect 2188 2496 2194 2508
rect 2444 2499 2502 2505
rect 2444 2496 2456 2499
rect 2188 2468 2456 2496
rect 2188 2456 2194 2468
rect 2444 2465 2456 2468
rect 2490 2496 2502 2499
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 2490 2468 2881 2496
rect 2490 2465 2502 2468
rect 2444 2459 2502 2465
rect 2869 2465 2881 2468
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 1535 2431 1593 2437
rect 1535 2397 1547 2431
rect 1581 2428 1593 2431
rect 11146 2428 11152 2440
rect 1581 2400 11152 2428
rect 1581 2397 1593 2400
rect 1535 2391 1593 2397
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 4154 76 4160 128
rect 4212 116 4218 128
rect 5258 116 5264 128
rect 4212 88 5264 116
rect 4212 76 4218 88
rect 5258 76 5264 88
rect 5316 76 5322 128
rect 11054 76 11060 128
rect 11112 116 11118 128
rect 12250 116 12256 128
rect 11112 88 12256 116
rect 11112 76 11118 88
rect 12250 76 12256 88
rect 12308 76 12314 128
rect 17954 76 17960 128
rect 18012 116 18018 128
rect 19242 116 19248 128
rect 18012 88 19248 116
rect 18012 76 18018 88
rect 19242 76 19248 88
rect 19300 76 19306 128
<< via1 >>
rect 2504 26188 2556 26240
rect 18236 26188 18288 26240
rect 1492 26120 1544 26172
rect 16580 26120 16632 26172
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 112 25440 164 25492
rect 15660 25440 15712 25492
rect 17040 25440 17092 25492
rect 2872 25372 2924 25424
rect 2504 25347 2556 25356
rect 2504 25313 2513 25347
rect 2513 25313 2547 25347
rect 2547 25313 2556 25347
rect 2504 25304 2556 25313
rect 6092 25304 6144 25356
rect 8300 25347 8352 25356
rect 8300 25313 8309 25347
rect 8309 25313 8343 25347
rect 8343 25313 8352 25347
rect 8300 25304 8352 25313
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 11796 25304 11848 25356
rect 12900 25347 12952 25356
rect 12900 25313 12909 25347
rect 12909 25313 12943 25347
rect 12943 25313 12952 25347
rect 12900 25304 12952 25313
rect 13912 25347 13964 25356
rect 13912 25313 13921 25347
rect 13921 25313 13955 25347
rect 13955 25313 13964 25347
rect 13912 25304 13964 25313
rect 16580 25347 16632 25356
rect 16580 25313 16589 25347
rect 16589 25313 16623 25347
rect 16623 25313 16632 25347
rect 16580 25304 16632 25313
rect 18236 25347 18288 25356
rect 18236 25313 18245 25347
rect 18245 25313 18279 25347
rect 18279 25313 18288 25347
rect 18236 25304 18288 25313
rect 19340 25347 19392 25356
rect 19340 25313 19349 25347
rect 19349 25313 19383 25347
rect 19383 25313 19392 25347
rect 19340 25304 19392 25313
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 2412 25279 2464 25288
rect 2412 25245 2421 25279
rect 2421 25245 2455 25279
rect 2455 25245 2464 25279
rect 2412 25236 2464 25245
rect 5172 25279 5224 25288
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 5172 25236 5224 25245
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7748 25236 7800 25245
rect 15476 25236 15528 25288
rect 3056 25100 3108 25152
rect 10048 25143 10100 25152
rect 10048 25109 10057 25143
rect 10057 25109 10091 25143
rect 10091 25109 10100 25143
rect 10048 25100 10100 25109
rect 11888 25100 11940 25152
rect 13728 25100 13780 25152
rect 13820 25100 13872 25152
rect 15844 25100 15896 25152
rect 18604 25100 18656 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 5172 24896 5224 24948
rect 9864 24939 9916 24948
rect 9864 24905 9873 24939
rect 9873 24905 9907 24939
rect 9907 24905 9916 24939
rect 9864 24896 9916 24905
rect 11796 24939 11848 24948
rect 11796 24905 11805 24939
rect 11805 24905 11839 24939
rect 11839 24905 11848 24939
rect 11796 24896 11848 24905
rect 12900 24896 12952 24948
rect 13912 24896 13964 24948
rect 14832 24939 14884 24948
rect 14832 24905 14841 24939
rect 14841 24905 14875 24939
rect 14875 24905 14884 24939
rect 14832 24896 14884 24905
rect 15660 24939 15712 24948
rect 15660 24905 15669 24939
rect 15669 24905 15703 24939
rect 15703 24905 15712 24939
rect 15660 24896 15712 24905
rect 16580 24939 16632 24948
rect 16580 24905 16589 24939
rect 16589 24905 16623 24939
rect 16623 24905 16632 24939
rect 16580 24896 16632 24905
rect 18236 24896 18288 24948
rect 5356 24828 5408 24880
rect 18604 24828 18656 24880
rect 1400 24760 1452 24812
rect 1952 24803 2004 24812
rect 1952 24769 1961 24803
rect 1961 24769 1995 24803
rect 1995 24769 2004 24803
rect 1952 24760 2004 24769
rect 6092 24760 6144 24812
rect 9772 24760 9824 24812
rect 4252 24735 4304 24744
rect 4252 24701 4261 24735
rect 4261 24701 4295 24735
rect 4295 24701 4304 24735
rect 4252 24692 4304 24701
rect 6552 24692 6604 24744
rect 8484 24735 8536 24744
rect 8484 24701 8493 24735
rect 8493 24701 8527 24735
rect 8527 24701 8536 24735
rect 8484 24692 8536 24701
rect 10876 24735 10928 24744
rect 10876 24701 10885 24735
rect 10885 24701 10919 24735
rect 10919 24701 10928 24735
rect 10876 24692 10928 24701
rect 12256 24735 12308 24744
rect 12256 24701 12265 24735
rect 12265 24701 12299 24735
rect 12299 24701 12308 24735
rect 12256 24692 12308 24701
rect 14832 24692 14884 24744
rect 2228 24624 2280 24676
rect 2596 24667 2648 24676
rect 2596 24633 2605 24667
rect 2605 24633 2639 24667
rect 2639 24633 2648 24667
rect 2596 24624 2648 24633
rect 5264 24667 5316 24676
rect 5264 24633 5273 24667
rect 5273 24633 5307 24667
rect 5307 24633 5316 24667
rect 5264 24624 5316 24633
rect 2504 24556 2556 24608
rect 3884 24599 3936 24608
rect 3884 24565 3893 24599
rect 3893 24565 3927 24599
rect 3927 24565 3936 24599
rect 3884 24556 3936 24565
rect 5172 24556 5224 24608
rect 6460 24624 6512 24676
rect 6828 24667 6880 24676
rect 6828 24633 6837 24667
rect 6837 24633 6871 24667
rect 6871 24633 6880 24667
rect 6828 24624 6880 24633
rect 10784 24667 10836 24676
rect 10784 24633 10793 24667
rect 10793 24633 10827 24667
rect 10827 24633 10836 24667
rect 10784 24624 10836 24633
rect 12440 24667 12492 24676
rect 12440 24633 12449 24667
rect 12449 24633 12483 24667
rect 12483 24633 12492 24667
rect 12440 24624 12492 24633
rect 14556 24624 14608 24676
rect 15476 24760 15528 24812
rect 15936 24692 15988 24744
rect 17960 24692 18012 24744
rect 18972 24692 19024 24744
rect 17132 24624 17184 24676
rect 18696 24624 18748 24676
rect 19340 24624 19392 24676
rect 8300 24556 8352 24608
rect 8852 24599 8904 24608
rect 8852 24565 8861 24599
rect 8861 24565 8895 24599
rect 8895 24565 8904 24599
rect 8852 24556 8904 24565
rect 16488 24556 16540 24608
rect 16948 24599 17000 24608
rect 16948 24565 16957 24599
rect 16957 24565 16991 24599
rect 16991 24565 17000 24599
rect 16948 24556 17000 24565
rect 17040 24556 17092 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1952 24395 2004 24404
rect 1952 24361 1961 24395
rect 1961 24361 1995 24395
rect 1995 24361 2004 24395
rect 1952 24352 2004 24361
rect 4344 24352 4396 24404
rect 6828 24352 6880 24404
rect 11888 24395 11940 24404
rect 11888 24361 11897 24395
rect 11897 24361 11931 24395
rect 11931 24361 11940 24395
rect 11888 24352 11940 24361
rect 2320 24327 2372 24336
rect 2320 24293 2329 24327
rect 2329 24293 2363 24327
rect 2363 24293 2372 24327
rect 2320 24284 2372 24293
rect 4252 24327 4304 24336
rect 4252 24293 4261 24327
rect 4261 24293 4295 24327
rect 4295 24293 4304 24327
rect 4252 24284 4304 24293
rect 4988 24284 5040 24336
rect 6092 24284 6144 24336
rect 6460 24284 6512 24336
rect 8300 24284 8352 24336
rect 9864 24284 9916 24336
rect 21180 24352 21232 24404
rect 12256 24327 12308 24336
rect 12256 24293 12265 24327
rect 12265 24293 12299 24327
rect 12299 24293 12308 24327
rect 12256 24284 12308 24293
rect 14096 24259 14148 24268
rect 14096 24225 14105 24259
rect 14105 24225 14139 24259
rect 14139 24225 14148 24259
rect 14096 24216 14148 24225
rect 15752 24284 15804 24336
rect 18052 24284 18104 24336
rect 19064 24216 19116 24268
rect 19499 24259 19551 24268
rect 19499 24225 19508 24259
rect 19508 24225 19542 24259
rect 19542 24225 19551 24259
rect 19499 24216 19551 24225
rect 2596 24191 2648 24200
rect 2136 24080 2188 24132
rect 2596 24157 2605 24191
rect 2605 24157 2639 24191
rect 2639 24157 2648 24191
rect 2596 24148 2648 24157
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4620 24148 4672 24200
rect 6368 24148 6420 24200
rect 8392 24191 8444 24200
rect 8392 24157 8401 24191
rect 8401 24157 8435 24191
rect 8435 24157 8444 24191
rect 8392 24148 8444 24157
rect 9772 24148 9824 24200
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10692 24148 10744 24157
rect 13176 24148 13228 24200
rect 14372 24191 14424 24200
rect 14372 24157 14381 24191
rect 14381 24157 14415 24191
rect 14415 24157 14424 24191
rect 14372 24148 14424 24157
rect 8576 24080 8628 24132
rect 17868 24080 17920 24132
rect 5264 24055 5316 24064
rect 5264 24021 5273 24055
rect 5273 24021 5307 24055
rect 5307 24021 5316 24055
rect 5264 24012 5316 24021
rect 6828 24012 6880 24064
rect 14648 24012 14700 24064
rect 15936 24055 15988 24064
rect 15936 24021 15945 24055
rect 15945 24021 15979 24055
rect 15979 24021 15988 24055
rect 15936 24012 15988 24021
rect 16396 24012 16448 24064
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2320 23808 2372 23860
rect 2596 23851 2648 23860
rect 2596 23817 2605 23851
rect 2605 23817 2639 23851
rect 2639 23817 2648 23851
rect 2596 23808 2648 23817
rect 3884 23808 3936 23860
rect 5540 23808 5592 23860
rect 6368 23851 6420 23860
rect 6368 23817 6377 23851
rect 6377 23817 6411 23851
rect 6411 23817 6420 23851
rect 6368 23808 6420 23817
rect 8852 23808 8904 23860
rect 9864 23851 9916 23860
rect 9864 23817 9873 23851
rect 9873 23817 9907 23851
rect 9907 23817 9916 23851
rect 9864 23808 9916 23817
rect 10784 23808 10836 23860
rect 12256 23808 12308 23860
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 14372 23808 14424 23860
rect 15752 23851 15804 23860
rect 15752 23817 15761 23851
rect 15761 23817 15795 23851
rect 15795 23817 15804 23851
rect 15752 23808 15804 23817
rect 18788 23808 18840 23860
rect 19064 23851 19116 23860
rect 19064 23817 19073 23851
rect 19073 23817 19107 23851
rect 19107 23817 19116 23851
rect 19064 23808 19116 23817
rect 22192 23808 22244 23860
rect 27344 23808 27396 23860
rect 1860 23672 1912 23724
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 2320 23672 2372 23724
rect 4160 23672 4212 23724
rect 4620 23715 4672 23724
rect 4620 23681 4629 23715
rect 4629 23681 4663 23715
rect 4663 23681 4672 23715
rect 4620 23672 4672 23681
rect 8116 23672 8168 23724
rect 8392 23672 8444 23724
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 1768 23579 1820 23588
rect 1768 23545 1777 23579
rect 1777 23545 1811 23579
rect 1811 23545 1820 23579
rect 2964 23579 3016 23588
rect 1768 23536 1820 23545
rect 2964 23545 2973 23579
rect 2973 23545 3007 23579
rect 3007 23545 3016 23579
rect 2964 23536 3016 23545
rect 3884 23468 3936 23520
rect 4988 23511 5040 23520
rect 4988 23477 4997 23511
rect 4997 23477 5031 23511
rect 5031 23477 5040 23511
rect 4988 23468 5040 23477
rect 7380 23579 7432 23588
rect 7380 23545 7389 23579
rect 7389 23545 7423 23579
rect 7423 23545 7432 23579
rect 7380 23536 7432 23545
rect 5540 23468 5592 23520
rect 6092 23511 6144 23520
rect 6092 23477 6101 23511
rect 6101 23477 6135 23511
rect 6135 23477 6144 23511
rect 6092 23468 6144 23477
rect 7748 23536 7800 23588
rect 11336 23672 11388 23724
rect 12716 23672 12768 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 14464 23672 14516 23724
rect 20076 23740 20128 23792
rect 25044 23740 25096 23792
rect 16396 23672 16448 23724
rect 19524 23672 19576 23724
rect 16488 23604 16540 23656
rect 18144 23647 18196 23656
rect 18144 23613 18153 23647
rect 18153 23613 18187 23647
rect 18187 23613 18196 23647
rect 18144 23604 18196 23613
rect 19248 23647 19300 23656
rect 19248 23613 19257 23647
rect 19257 23613 19291 23647
rect 19291 23613 19300 23647
rect 19248 23604 19300 23613
rect 11520 23579 11572 23588
rect 7932 23468 7984 23520
rect 8852 23468 8904 23520
rect 10784 23468 10836 23520
rect 11520 23545 11529 23579
rect 11529 23545 11563 23579
rect 11563 23545 11572 23579
rect 11520 23536 11572 23545
rect 14372 23536 14424 23588
rect 14924 23536 14976 23588
rect 21732 23604 21784 23656
rect 22100 23604 22152 23656
rect 20076 23536 20128 23588
rect 23480 23536 23532 23588
rect 14096 23468 14148 23520
rect 19984 23468 20036 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2228 23307 2280 23316
rect 2228 23273 2237 23307
rect 2237 23273 2271 23307
rect 2271 23273 2280 23307
rect 2228 23264 2280 23273
rect 3148 23264 3200 23316
rect 14464 23264 14516 23316
rect 16948 23264 17000 23316
rect 18144 23264 18196 23316
rect 19248 23264 19300 23316
rect 6276 23196 6328 23248
rect 8208 23239 8260 23248
rect 8208 23205 8217 23239
rect 8217 23205 8251 23239
rect 8251 23205 8260 23239
rect 8208 23196 8260 23205
rect 8484 23196 8536 23248
rect 9220 23196 9272 23248
rect 10876 23196 10928 23248
rect 11520 23196 11572 23248
rect 12440 23196 12492 23248
rect 12716 23239 12768 23248
rect 12716 23205 12725 23239
rect 12725 23205 12759 23239
rect 12759 23205 12768 23239
rect 12716 23196 12768 23205
rect 14188 23196 14240 23248
rect 2596 23171 2648 23180
rect 2596 23137 2605 23171
rect 2605 23137 2639 23171
rect 2639 23137 2648 23171
rect 2596 23128 2648 23137
rect 4528 23128 4580 23180
rect 3608 23060 3660 23112
rect 6000 23060 6052 23112
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 8116 23060 8168 23069
rect 9588 23060 9640 23112
rect 10692 23060 10744 23112
rect 11888 23060 11940 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14924 23128 14976 23180
rect 15660 23171 15712 23180
rect 15660 23137 15669 23171
rect 15669 23137 15703 23171
rect 15703 23137 15712 23171
rect 15660 23128 15712 23137
rect 17224 23171 17276 23180
rect 17224 23137 17233 23171
rect 17233 23137 17267 23171
rect 17267 23137 17276 23171
rect 17224 23128 17276 23137
rect 7196 22992 7248 23044
rect 8944 22992 8996 23044
rect 14832 23060 14884 23112
rect 16672 23060 16724 23112
rect 19892 23128 19944 23180
rect 18880 23060 18932 23112
rect 14280 23035 14332 23044
rect 14280 23001 14289 23035
rect 14289 23001 14323 23035
rect 14323 23001 14332 23035
rect 14280 22992 14332 23001
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 1860 22924 1912 22976
rect 3332 22924 3384 22976
rect 5080 22967 5132 22976
rect 5080 22933 5089 22967
rect 5089 22933 5123 22967
rect 5123 22933 5132 22967
rect 5080 22924 5132 22933
rect 5264 22924 5316 22976
rect 7380 22967 7432 22976
rect 7380 22933 7389 22967
rect 7389 22933 7423 22967
rect 7423 22933 7432 22967
rect 7380 22924 7432 22933
rect 8300 22924 8352 22976
rect 8760 22924 8812 22976
rect 9772 22924 9824 22976
rect 12992 22967 13044 22976
rect 12992 22933 13001 22967
rect 13001 22933 13035 22967
rect 13035 22933 13044 22967
rect 12992 22924 13044 22933
rect 16396 22967 16448 22976
rect 16396 22933 16405 22967
rect 16405 22933 16439 22967
rect 16439 22933 16448 22967
rect 16396 22924 16448 22933
rect 18052 22924 18104 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2596 22720 2648 22772
rect 5264 22720 5316 22772
rect 6092 22720 6144 22772
rect 8208 22720 8260 22772
rect 9588 22763 9640 22772
rect 9588 22729 9597 22763
rect 9597 22729 9631 22763
rect 9631 22729 9640 22763
rect 9588 22720 9640 22729
rect 10048 22763 10100 22772
rect 10048 22729 10057 22763
rect 10057 22729 10091 22763
rect 10091 22729 10100 22763
rect 10048 22720 10100 22729
rect 12440 22720 12492 22772
rect 14096 22720 14148 22772
rect 14188 22763 14240 22772
rect 14188 22729 14197 22763
rect 14197 22729 14231 22763
rect 14231 22729 14240 22763
rect 15660 22763 15712 22772
rect 14188 22720 14240 22729
rect 15660 22729 15669 22763
rect 15669 22729 15703 22763
rect 15703 22729 15712 22763
rect 15660 22720 15712 22729
rect 2872 22652 2924 22704
rect 4896 22652 4948 22704
rect 2320 22627 2372 22636
rect 2320 22593 2329 22627
rect 2329 22593 2363 22627
rect 2363 22593 2372 22627
rect 2320 22584 2372 22593
rect 11612 22652 11664 22704
rect 17224 22720 17276 22772
rect 18880 22763 18932 22772
rect 18880 22729 18889 22763
rect 18889 22729 18923 22763
rect 18923 22729 18932 22763
rect 18880 22720 18932 22729
rect 19064 22720 19116 22772
rect 19892 22763 19944 22772
rect 19892 22729 19901 22763
rect 19901 22729 19935 22763
rect 19935 22729 19944 22763
rect 19892 22720 19944 22729
rect 16488 22652 16540 22704
rect 3700 22559 3752 22568
rect 3700 22525 3709 22559
rect 3709 22525 3743 22559
rect 3743 22525 3752 22559
rect 3700 22516 3752 22525
rect 2320 22448 2372 22500
rect 3608 22448 3660 22500
rect 4804 22516 4856 22568
rect 5080 22516 5132 22568
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 14280 22584 14332 22636
rect 15476 22584 15528 22636
rect 16672 22627 16724 22636
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 4528 22423 4580 22432
rect 4528 22389 4537 22423
rect 4537 22389 4571 22423
rect 4571 22389 4580 22423
rect 4528 22380 4580 22389
rect 5080 22380 5132 22432
rect 5448 22448 5500 22500
rect 6276 22423 6328 22432
rect 6276 22389 6285 22423
rect 6285 22389 6319 22423
rect 6319 22389 6328 22423
rect 6276 22380 6328 22389
rect 7196 22516 7248 22568
rect 9036 22516 9088 22568
rect 12256 22516 12308 22568
rect 12992 22516 13044 22568
rect 18512 22559 18564 22568
rect 18512 22525 18521 22559
rect 18521 22525 18555 22559
rect 18555 22525 18564 22559
rect 18512 22516 18564 22525
rect 19524 22516 19576 22568
rect 8852 22448 8904 22500
rect 14740 22491 14792 22500
rect 10048 22380 10100 22432
rect 14740 22457 14749 22491
rect 14749 22457 14783 22491
rect 14783 22457 14792 22491
rect 14740 22448 14792 22457
rect 14832 22491 14884 22500
rect 14832 22457 14841 22491
rect 14841 22457 14875 22491
rect 14875 22457 14884 22491
rect 16396 22491 16448 22500
rect 14832 22448 14884 22457
rect 16396 22457 16405 22491
rect 16405 22457 16439 22491
rect 16439 22457 16448 22491
rect 16396 22448 16448 22457
rect 16488 22491 16540 22500
rect 16488 22457 16497 22491
rect 16497 22457 16531 22491
rect 16531 22457 16540 22491
rect 16488 22448 16540 22457
rect 10876 22380 10928 22432
rect 11244 22423 11296 22432
rect 11244 22389 11253 22423
rect 11253 22389 11287 22423
rect 11287 22389 11296 22423
rect 11244 22380 11296 22389
rect 12808 22423 12860 22432
rect 12808 22389 12817 22423
rect 12817 22389 12851 22423
rect 12851 22389 12860 22423
rect 12808 22380 12860 22389
rect 16580 22380 16632 22432
rect 19524 22423 19576 22432
rect 19524 22389 19533 22423
rect 19533 22389 19567 22423
rect 19567 22389 19576 22423
rect 19524 22380 19576 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2872 22176 2924 22228
rect 4988 22176 5040 22228
rect 7932 22176 7984 22228
rect 8760 22219 8812 22228
rect 8760 22185 8769 22219
rect 8769 22185 8803 22219
rect 8803 22185 8812 22219
rect 8760 22176 8812 22185
rect 11244 22219 11296 22228
rect 11244 22185 11253 22219
rect 11253 22185 11287 22219
rect 11287 22185 11296 22219
rect 11244 22176 11296 22185
rect 12164 22176 12216 22228
rect 13728 22219 13780 22228
rect 13728 22185 13737 22219
rect 13737 22185 13771 22219
rect 13771 22185 13780 22219
rect 13728 22176 13780 22185
rect 14740 22219 14792 22228
rect 14740 22185 14749 22219
rect 14749 22185 14783 22219
rect 14783 22185 14792 22219
rect 14740 22176 14792 22185
rect 15476 22219 15528 22228
rect 15476 22185 15485 22219
rect 15485 22185 15519 22219
rect 15519 22185 15528 22219
rect 15476 22176 15528 22185
rect 24216 22176 24268 22228
rect 1676 22151 1728 22160
rect 1676 22117 1685 22151
rect 1685 22117 1719 22151
rect 1719 22117 1728 22151
rect 1676 22108 1728 22117
rect 5166 22151 5218 22160
rect 5166 22117 5175 22151
rect 5175 22117 5209 22151
rect 5209 22117 5218 22151
rect 5166 22108 5218 22117
rect 6276 22108 6328 22160
rect 6460 22108 6512 22160
rect 8024 22108 8076 22160
rect 8852 22108 8904 22160
rect 10416 22108 10468 22160
rect 12808 22108 12860 22160
rect 15936 22108 15988 22160
rect 16672 22108 16724 22160
rect 2320 22083 2372 22092
rect 2320 22049 2329 22083
rect 2329 22049 2363 22083
rect 2363 22049 2372 22083
rect 2320 22040 2372 22049
rect 9956 22040 10008 22092
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 14096 22040 14148 22092
rect 15568 22040 15620 22092
rect 17132 22040 17184 22092
rect 18420 22040 18472 22092
rect 19524 22040 19576 22092
rect 21364 22083 21416 22092
rect 21364 22049 21373 22083
rect 21373 22049 21407 22083
rect 21407 22049 21416 22083
rect 21364 22040 21416 22049
rect 22468 22083 22520 22092
rect 22468 22049 22477 22083
rect 22477 22049 22511 22083
rect 22511 22049 22520 22083
rect 22468 22040 22520 22049
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 7932 21972 7984 22024
rect 1860 21904 1912 21956
rect 5356 21904 5408 21956
rect 12164 21972 12216 22024
rect 12624 21972 12676 22024
rect 14740 21972 14792 22024
rect 12900 21904 12952 21956
rect 23204 21904 23256 21956
rect 3608 21836 3660 21888
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 10140 21879 10192 21888
rect 10140 21845 10149 21879
rect 10149 21845 10183 21879
rect 10183 21845 10192 21879
rect 10140 21836 10192 21845
rect 13636 21836 13688 21888
rect 15568 21836 15620 21888
rect 17500 21836 17552 21888
rect 18512 21836 18564 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2688 21632 2740 21684
rect 4804 21632 4856 21684
rect 8024 21632 8076 21684
rect 9772 21632 9824 21684
rect 10416 21675 10468 21684
rect 10416 21641 10425 21675
rect 10425 21641 10459 21675
rect 10459 21641 10468 21675
rect 10416 21632 10468 21641
rect 10692 21632 10744 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 14188 21632 14240 21684
rect 16488 21632 16540 21684
rect 17132 21632 17184 21684
rect 1768 21564 1820 21616
rect 2320 21564 2372 21616
rect 6644 21496 6696 21548
rect 6828 21539 6880 21548
rect 6828 21505 6837 21539
rect 6837 21505 6871 21539
rect 6871 21505 6880 21539
rect 6828 21496 6880 21505
rect 5632 21428 5684 21480
rect 8484 21428 8536 21480
rect 2228 21403 2280 21412
rect 2228 21369 2237 21403
rect 2237 21369 2271 21403
rect 2271 21369 2280 21403
rect 2228 21360 2280 21369
rect 2320 21403 2372 21412
rect 2320 21369 2329 21403
rect 2329 21369 2363 21403
rect 2363 21369 2372 21403
rect 2872 21403 2924 21412
rect 2320 21360 2372 21369
rect 2872 21369 2881 21403
rect 2881 21369 2915 21403
rect 2915 21369 2924 21403
rect 2872 21360 2924 21369
rect 5080 21360 5132 21412
rect 10968 21564 11020 21616
rect 14096 21607 14148 21616
rect 14096 21573 14105 21607
rect 14105 21573 14139 21607
rect 14139 21573 14148 21607
rect 14096 21564 14148 21573
rect 22468 21607 22520 21616
rect 22468 21573 22477 21607
rect 22477 21573 22511 21607
rect 22511 21573 22520 21607
rect 22468 21564 22520 21573
rect 21364 21539 21416 21548
rect 21364 21505 21373 21539
rect 21373 21505 21407 21539
rect 21407 21505 21416 21539
rect 21364 21496 21416 21505
rect 10876 21471 10928 21480
rect 10876 21437 10885 21471
rect 10885 21437 10919 21471
rect 10919 21437 10928 21471
rect 10876 21428 10928 21437
rect 10968 21428 11020 21480
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 14648 21471 14700 21480
rect 14648 21437 14657 21471
rect 14657 21437 14691 21471
rect 14691 21437 14700 21471
rect 14648 21428 14700 21437
rect 15936 21471 15988 21480
rect 15936 21437 15945 21471
rect 15945 21437 15979 21471
rect 15979 21437 15988 21471
rect 15936 21428 15988 21437
rect 12164 21360 12216 21412
rect 12808 21360 12860 21412
rect 15292 21360 15344 21412
rect 18788 21428 18840 21480
rect 18328 21360 18380 21412
rect 7932 21292 7984 21344
rect 18512 21335 18564 21344
rect 18512 21301 18521 21335
rect 18521 21301 18555 21335
rect 18555 21301 18564 21335
rect 18512 21292 18564 21301
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1768 21131 1820 21140
rect 1768 21097 1777 21131
rect 1777 21097 1811 21131
rect 1811 21097 1820 21131
rect 1768 21088 1820 21097
rect 2320 21088 2372 21140
rect 4252 21131 4304 21140
rect 4252 21097 4261 21131
rect 4261 21097 4295 21131
rect 4295 21097 4304 21131
rect 4252 21088 4304 21097
rect 5632 21131 5684 21140
rect 5632 21097 5641 21131
rect 5641 21097 5675 21131
rect 5675 21097 5684 21131
rect 5632 21088 5684 21097
rect 7932 21131 7984 21140
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 9864 21088 9916 21140
rect 10876 21088 10928 21140
rect 3700 21020 3752 21072
rect 5080 21020 5132 21072
rect 3240 20952 3292 21004
rect 3792 20884 3844 20936
rect 5172 20952 5224 21004
rect 6276 21020 6328 21072
rect 9036 21020 9088 21072
rect 10692 21020 10744 21072
rect 12256 21063 12308 21072
rect 12256 21029 12265 21063
rect 12265 21029 12299 21063
rect 12299 21029 12308 21063
rect 12256 21020 12308 21029
rect 12900 21088 12952 21140
rect 17316 21063 17368 21072
rect 6092 20995 6144 21004
rect 6092 20961 6101 20995
rect 6101 20961 6135 20995
rect 6135 20961 6144 20995
rect 6092 20952 6144 20961
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 8300 20952 8352 20961
rect 8484 20995 8536 21004
rect 8484 20961 8493 20995
rect 8493 20961 8527 20995
rect 8527 20961 8536 20995
rect 8484 20952 8536 20961
rect 11796 20995 11848 21004
rect 11796 20961 11805 20995
rect 11805 20961 11839 20995
rect 11839 20961 11848 20995
rect 11796 20952 11848 20961
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 12164 20952 12216 21004
rect 17316 21029 17325 21063
rect 17325 21029 17359 21063
rect 17359 21029 17368 21063
rect 17316 21020 17368 21029
rect 13452 20952 13504 21004
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 19064 20995 19116 21004
rect 19064 20961 19073 20995
rect 19073 20961 19107 20995
rect 19107 20961 19116 20995
rect 19064 20952 19116 20961
rect 5448 20748 5500 20800
rect 6920 20791 6972 20800
rect 6920 20757 6929 20791
rect 6929 20757 6963 20791
rect 6963 20757 6972 20791
rect 6920 20748 6972 20757
rect 9496 20791 9548 20800
rect 9496 20757 9505 20791
rect 9505 20757 9539 20791
rect 9539 20757 9548 20791
rect 9496 20748 9548 20757
rect 10968 20748 11020 20800
rect 14464 20884 14516 20936
rect 17224 20927 17276 20936
rect 17224 20893 17233 20927
rect 17233 20893 17267 20927
rect 17267 20893 17276 20927
rect 17224 20884 17276 20893
rect 18236 20884 18288 20936
rect 18788 20816 18840 20868
rect 12900 20748 12952 20800
rect 13176 20748 13228 20800
rect 14648 20791 14700 20800
rect 14648 20757 14657 20791
rect 14657 20757 14691 20791
rect 14691 20757 14700 20791
rect 14648 20748 14700 20757
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16488 20748 16540 20757
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 3884 20587 3936 20596
rect 3884 20553 3893 20587
rect 3893 20553 3927 20587
rect 3927 20553 3936 20587
rect 3884 20544 3936 20553
rect 6000 20544 6052 20596
rect 6276 20587 6328 20596
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 6276 20544 6328 20553
rect 9404 20544 9456 20596
rect 10692 20544 10744 20596
rect 14648 20544 14700 20596
rect 15476 20587 15528 20596
rect 15476 20553 15485 20587
rect 15485 20553 15519 20587
rect 15519 20553 15528 20587
rect 15476 20544 15528 20553
rect 3148 20476 3200 20528
rect 2872 20451 2924 20460
rect 2872 20417 2881 20451
rect 2881 20417 2915 20451
rect 2915 20417 2924 20451
rect 2872 20408 2924 20417
rect 3240 20408 3292 20460
rect 6460 20408 6512 20460
rect 2872 20272 2924 20324
rect 5172 20340 5224 20392
rect 5448 20340 5500 20392
rect 5908 20340 5960 20392
rect 6920 20340 6972 20392
rect 8300 20340 8352 20392
rect 11796 20476 11848 20528
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 11336 20451 11388 20460
rect 11336 20417 11345 20451
rect 11345 20417 11379 20451
rect 11379 20417 11388 20451
rect 11336 20408 11388 20417
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 14832 20451 14884 20460
rect 14832 20417 14841 20451
rect 14841 20417 14875 20451
rect 14875 20417 14884 20451
rect 14832 20408 14884 20417
rect 16488 20544 16540 20596
rect 17316 20544 17368 20596
rect 19064 20587 19116 20596
rect 19064 20553 19073 20587
rect 19073 20553 19107 20587
rect 19107 20553 19116 20587
rect 19064 20544 19116 20553
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 9496 20340 9548 20392
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 6644 20272 6696 20324
rect 9680 20272 9732 20324
rect 3148 20247 3200 20256
rect 3148 20213 3157 20247
rect 3157 20213 3191 20247
rect 3191 20213 3200 20247
rect 3148 20204 3200 20213
rect 8484 20247 8536 20256
rect 8484 20213 8493 20247
rect 8493 20213 8527 20247
rect 8527 20213 8536 20247
rect 8484 20204 8536 20213
rect 10968 20204 11020 20256
rect 11796 20247 11848 20256
rect 11796 20213 11805 20247
rect 11805 20213 11839 20247
rect 11839 20213 11848 20247
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 14648 20315 14700 20324
rect 14648 20281 14657 20315
rect 14657 20281 14691 20315
rect 14691 20281 14700 20315
rect 14648 20272 14700 20281
rect 16856 20272 16908 20324
rect 18144 20272 18196 20324
rect 18236 20315 18288 20324
rect 18236 20281 18245 20315
rect 18245 20281 18279 20315
rect 18279 20281 18288 20315
rect 18788 20315 18840 20324
rect 18236 20272 18288 20281
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 11796 20204 11848 20213
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2228 20000 2280 20052
rect 6000 20000 6052 20052
rect 9680 20000 9732 20052
rect 14556 20000 14608 20052
rect 17316 20000 17368 20052
rect 26332 20000 26384 20052
rect 1676 19932 1728 19984
rect 3056 19932 3108 19984
rect 4344 19932 4396 19984
rect 4804 19975 4856 19984
rect 4804 19941 4813 19975
rect 4813 19941 4847 19975
rect 4847 19941 4856 19975
rect 4804 19932 4856 19941
rect 5080 19932 5132 19984
rect 6368 19932 6420 19984
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 7104 19864 7156 19916
rect 8300 19907 8352 19916
rect 8300 19873 8309 19907
rect 8309 19873 8343 19907
rect 8343 19873 8352 19907
rect 8300 19864 8352 19873
rect 8760 19864 8812 19916
rect 10876 19932 10928 19984
rect 14188 19932 14240 19984
rect 15292 19932 15344 19984
rect 17960 19975 18012 19984
rect 17960 19941 17969 19975
rect 17969 19941 18003 19975
rect 18003 19941 18012 19975
rect 17960 19932 18012 19941
rect 9864 19864 9916 19916
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 12164 19907 12216 19916
rect 12164 19873 12173 19907
rect 12173 19873 12207 19907
rect 12207 19873 12216 19907
rect 12164 19864 12216 19873
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 24216 19864 24268 19916
rect 2136 19839 2188 19848
rect 2136 19805 2145 19839
rect 2145 19805 2179 19839
rect 2179 19805 2188 19839
rect 2136 19796 2188 19805
rect 4528 19796 4580 19848
rect 5908 19796 5960 19848
rect 8668 19839 8720 19848
rect 3240 19728 3292 19780
rect 3792 19771 3844 19780
rect 3792 19737 3801 19771
rect 3801 19737 3835 19771
rect 3835 19737 3844 19771
rect 3792 19728 3844 19737
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 13084 19796 13136 19848
rect 13820 19796 13872 19848
rect 15660 19796 15712 19848
rect 16028 19839 16080 19848
rect 16028 19805 16037 19839
rect 16037 19805 16071 19839
rect 16071 19805 16080 19839
rect 16028 19796 16080 19805
rect 18328 19839 18380 19848
rect 18328 19805 18337 19839
rect 18337 19805 18371 19839
rect 18371 19805 18380 19839
rect 18328 19796 18380 19805
rect 7932 19660 7984 19712
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 14832 19660 14884 19712
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 19524 19703 19576 19712
rect 19524 19669 19533 19703
rect 19533 19669 19567 19703
rect 19567 19669 19576 19703
rect 19524 19660 19576 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 4344 19456 4396 19508
rect 8300 19499 8352 19508
rect 8300 19465 8309 19499
rect 8309 19465 8343 19499
rect 8343 19465 8352 19499
rect 8300 19456 8352 19465
rect 9404 19456 9456 19508
rect 9864 19456 9916 19508
rect 12164 19499 12216 19508
rect 12164 19465 12173 19499
rect 12173 19465 12207 19499
rect 12207 19465 12216 19499
rect 12164 19456 12216 19465
rect 12808 19499 12860 19508
rect 12808 19465 12817 19499
rect 12817 19465 12851 19499
rect 12851 19465 12860 19499
rect 12808 19456 12860 19465
rect 14648 19456 14700 19508
rect 15292 19456 15344 19508
rect 17960 19456 18012 19508
rect 19340 19499 19392 19508
rect 19340 19465 19349 19499
rect 19349 19465 19383 19499
rect 19383 19465 19392 19499
rect 19340 19456 19392 19465
rect 2044 19388 2096 19440
rect 3516 19388 3568 19440
rect 4804 19388 4856 19440
rect 9588 19431 9640 19440
rect 9588 19397 9597 19431
rect 9597 19397 9631 19431
rect 9631 19397 9640 19431
rect 9588 19388 9640 19397
rect 10876 19388 10928 19440
rect 11796 19431 11848 19440
rect 11796 19397 11805 19431
rect 11805 19397 11839 19431
rect 11839 19397 11848 19431
rect 11796 19388 11848 19397
rect 19524 19388 19576 19440
rect 1676 19320 1728 19372
rect 3424 19320 3476 19372
rect 4528 19363 4580 19372
rect 4528 19329 4537 19363
rect 4537 19329 4571 19363
rect 4571 19329 4580 19363
rect 4528 19320 4580 19329
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 5172 19252 5224 19304
rect 2044 19184 2096 19236
rect 2228 19227 2280 19236
rect 2228 19193 2237 19227
rect 2237 19193 2271 19227
rect 2271 19193 2280 19227
rect 2228 19184 2280 19193
rect 6092 19252 6144 19304
rect 7656 19295 7708 19304
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 7932 19252 7984 19304
rect 9864 19320 9916 19372
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 16028 19320 16080 19372
rect 16856 19320 16908 19372
rect 24216 19320 24268 19372
rect 13084 19252 13136 19304
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 18696 19252 18748 19304
rect 4804 19116 4856 19168
rect 5172 19159 5224 19168
rect 5172 19125 5181 19159
rect 5181 19125 5215 19159
rect 5215 19125 5224 19159
rect 5172 19116 5224 19125
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 8024 19184 8076 19236
rect 9312 19227 9364 19236
rect 9312 19193 9321 19227
rect 9321 19193 9355 19227
rect 9355 19193 9364 19227
rect 9312 19184 9364 19193
rect 16396 19227 16448 19236
rect 16396 19193 16405 19227
rect 16405 19193 16439 19227
rect 16439 19193 16448 19227
rect 16396 19184 16448 19193
rect 7288 19116 7340 19168
rect 9864 19116 9916 19168
rect 10140 19116 10192 19168
rect 13360 19159 13412 19168
rect 13360 19125 13369 19159
rect 13369 19125 13403 19159
rect 13403 19125 13412 19159
rect 13360 19116 13412 19125
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 19064 19184 19116 19236
rect 14280 19116 14332 19125
rect 16856 19116 16908 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2044 18955 2096 18964
rect 2044 18921 2053 18955
rect 2053 18921 2087 18955
rect 2087 18921 2096 18955
rect 2044 18912 2096 18921
rect 2136 18912 2188 18964
rect 5080 18955 5132 18964
rect 2412 18844 2464 18896
rect 3424 18844 3476 18896
rect 5080 18921 5089 18955
rect 5089 18921 5123 18955
rect 5123 18921 5132 18955
rect 5080 18912 5132 18921
rect 8484 18912 8536 18964
rect 12992 18912 13044 18964
rect 4252 18887 4304 18896
rect 4252 18853 4261 18887
rect 4261 18853 4295 18887
rect 4295 18853 4304 18887
rect 4252 18844 4304 18853
rect 6184 18887 6236 18896
rect 6184 18853 6187 18887
rect 6187 18853 6221 18887
rect 6221 18853 6236 18887
rect 6184 18844 6236 18853
rect 6644 18844 6696 18896
rect 8024 18887 8076 18896
rect 8024 18853 8033 18887
rect 8033 18853 8067 18887
rect 8067 18853 8076 18887
rect 8024 18844 8076 18853
rect 6000 18776 6052 18828
rect 9404 18844 9456 18896
rect 13360 18844 13412 18896
rect 15476 18887 15528 18896
rect 15476 18853 15485 18887
rect 15485 18853 15519 18887
rect 15519 18853 15528 18887
rect 15476 18844 15528 18853
rect 3792 18708 3844 18760
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 2228 18640 2280 18692
rect 3148 18640 3200 18692
rect 8760 18819 8812 18828
rect 8760 18785 8769 18819
rect 8769 18785 8803 18819
rect 8803 18785 8812 18819
rect 8760 18776 8812 18785
rect 9496 18776 9548 18828
rect 11796 18776 11848 18828
rect 14280 18776 14332 18828
rect 16856 18819 16908 18828
rect 16856 18785 16865 18819
rect 16865 18785 16899 18819
rect 16899 18785 16908 18819
rect 16856 18776 16908 18785
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 19064 18819 19116 18828
rect 19064 18785 19073 18819
rect 19073 18785 19107 18819
rect 19107 18785 19116 18819
rect 19064 18776 19116 18785
rect 9036 18708 9088 18760
rect 10140 18708 10192 18760
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 1492 18572 1544 18624
rect 3516 18572 3568 18624
rect 7932 18640 7984 18692
rect 11612 18640 11664 18692
rect 12808 18640 12860 18692
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 7656 18572 7708 18624
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 9404 18572 9456 18624
rect 9680 18572 9732 18624
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 10784 18615 10836 18624
rect 10784 18581 10793 18615
rect 10793 18581 10827 18615
rect 10827 18581 10836 18615
rect 10784 18572 10836 18581
rect 11796 18615 11848 18624
rect 11796 18581 11805 18615
rect 11805 18581 11839 18615
rect 11839 18581 11848 18615
rect 11796 18572 11848 18581
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 18144 18615 18196 18624
rect 18144 18581 18153 18615
rect 18153 18581 18187 18615
rect 18187 18581 18196 18615
rect 18144 18572 18196 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2412 18411 2464 18420
rect 2412 18377 2421 18411
rect 2421 18377 2455 18411
rect 2455 18377 2464 18411
rect 2412 18368 2464 18377
rect 2504 18368 2556 18420
rect 1492 18139 1544 18148
rect 1492 18105 1501 18139
rect 1501 18105 1535 18139
rect 1535 18105 1544 18139
rect 1492 18096 1544 18105
rect 1676 18096 1728 18148
rect 2688 18096 2740 18148
rect 4252 18368 4304 18420
rect 4804 18368 4856 18420
rect 6552 18368 6604 18420
rect 9680 18368 9732 18420
rect 10784 18368 10836 18420
rect 10968 18411 11020 18420
rect 10968 18377 10977 18411
rect 10977 18377 11011 18411
rect 11011 18377 11020 18411
rect 10968 18368 11020 18377
rect 12164 18368 12216 18420
rect 13452 18368 13504 18420
rect 15476 18368 15528 18420
rect 16856 18411 16908 18420
rect 5264 18300 5316 18352
rect 6184 18343 6236 18352
rect 6184 18309 6193 18343
rect 6193 18309 6227 18343
rect 6227 18309 6236 18343
rect 6184 18300 6236 18309
rect 9496 18300 9548 18352
rect 10324 18300 10376 18352
rect 12532 18300 12584 18352
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 3148 18232 3200 18241
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 6552 18232 6604 18284
rect 4712 18164 4764 18216
rect 7012 18232 7064 18284
rect 8300 18232 8352 18284
rect 9588 18232 9640 18284
rect 9956 18232 10008 18284
rect 10140 18232 10192 18284
rect 10968 18232 11020 18284
rect 13544 18300 13596 18352
rect 16856 18377 16865 18411
rect 16865 18377 16899 18411
rect 16899 18377 16908 18411
rect 16856 18368 16908 18377
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 15844 18300 15896 18352
rect 18696 18343 18748 18352
rect 4988 18096 5040 18148
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 5448 18028 5500 18080
rect 6552 18071 6604 18080
rect 6552 18037 6561 18071
rect 6561 18037 6595 18071
rect 6595 18037 6604 18071
rect 6552 18028 6604 18037
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 9864 18164 9916 18216
rect 8576 18071 8628 18080
rect 8576 18037 8585 18071
rect 8585 18037 8619 18071
rect 8619 18037 8628 18071
rect 8576 18028 8628 18037
rect 10048 18028 10100 18080
rect 10232 18164 10284 18216
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 14372 18275 14424 18284
rect 12808 18232 12860 18241
rect 10324 18139 10376 18148
rect 10324 18105 10333 18139
rect 10333 18105 10367 18139
rect 10367 18105 10376 18139
rect 10324 18096 10376 18105
rect 10784 18096 10836 18148
rect 12532 18164 12584 18216
rect 12440 18139 12492 18148
rect 12440 18105 12449 18139
rect 12449 18105 12483 18139
rect 12483 18105 12492 18139
rect 12440 18096 12492 18105
rect 13268 18096 13320 18148
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 18696 18309 18705 18343
rect 18705 18309 18739 18343
rect 18739 18309 18748 18343
rect 18696 18300 18748 18309
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 14464 18139 14516 18148
rect 14464 18105 14473 18139
rect 14473 18105 14507 18139
rect 14507 18105 14516 18139
rect 14464 18096 14516 18105
rect 16580 18139 16632 18148
rect 13360 18028 13412 18080
rect 15568 18028 15620 18080
rect 15752 18071 15804 18080
rect 15752 18037 15761 18071
rect 15761 18037 15795 18071
rect 15795 18037 15804 18071
rect 16580 18105 16589 18139
rect 16589 18105 16623 18139
rect 16623 18105 16632 18139
rect 16580 18096 16632 18105
rect 18236 18139 18288 18148
rect 18236 18105 18245 18139
rect 18245 18105 18279 18139
rect 18279 18105 18288 18139
rect 18236 18096 18288 18105
rect 15752 18028 15804 18037
rect 17592 18028 17644 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 4712 17867 4764 17876
rect 4712 17833 4721 17867
rect 4721 17833 4755 17867
rect 4755 17833 4764 17867
rect 4712 17824 4764 17833
rect 4988 17824 5040 17876
rect 6000 17867 6052 17876
rect 6000 17833 6009 17867
rect 6009 17833 6043 17867
rect 6043 17833 6052 17867
rect 6000 17824 6052 17833
rect 9404 17824 9456 17876
rect 12440 17824 12492 17876
rect 13452 17867 13504 17876
rect 13452 17833 13461 17867
rect 13461 17833 13495 17867
rect 13495 17833 13504 17867
rect 13452 17824 13504 17833
rect 13728 17867 13780 17876
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 13820 17824 13872 17876
rect 15384 17824 15436 17876
rect 15844 17867 15896 17876
rect 15844 17833 15853 17867
rect 15853 17833 15887 17867
rect 15887 17833 15896 17867
rect 15844 17824 15896 17833
rect 16396 17824 16448 17876
rect 2136 17799 2188 17808
rect 2136 17765 2145 17799
rect 2145 17765 2179 17799
rect 2179 17765 2188 17799
rect 2136 17756 2188 17765
rect 5264 17756 5316 17808
rect 9312 17756 9364 17808
rect 10600 17756 10652 17808
rect 12900 17756 12952 17808
rect 19340 17824 19392 17876
rect 18328 17799 18380 17808
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 8760 17688 8812 17740
rect 10324 17688 10376 17740
rect 10784 17688 10836 17740
rect 11980 17688 12032 17740
rect 12532 17731 12584 17740
rect 2504 17620 2556 17672
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 3056 17620 3108 17672
rect 4160 17620 4212 17672
rect 5172 17620 5224 17672
rect 7288 17552 7340 17604
rect 7748 17552 7800 17604
rect 10048 17620 10100 17672
rect 12532 17697 12541 17731
rect 12541 17697 12575 17731
rect 12575 17697 12584 17731
rect 12532 17688 12584 17697
rect 13544 17688 13596 17740
rect 18328 17765 18337 17799
rect 18337 17765 18371 17799
rect 18371 17765 18380 17799
rect 18328 17756 18380 17765
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 19432 17688 19484 17740
rect 16764 17620 16816 17672
rect 18420 17620 18472 17672
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 9588 17552 9640 17604
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 3516 17527 3568 17536
rect 3516 17493 3525 17527
rect 3525 17493 3559 17527
rect 3559 17493 3568 17527
rect 3516 17484 3568 17493
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 8668 17484 8720 17536
rect 9496 17527 9548 17536
rect 9496 17493 9505 17527
rect 9505 17493 9539 17527
rect 9539 17493 9548 17527
rect 9496 17484 9548 17493
rect 9956 17527 10008 17536
rect 9956 17493 9965 17527
rect 9965 17493 9999 17527
rect 9999 17493 10008 17527
rect 9956 17484 10008 17493
rect 10140 17484 10192 17536
rect 10968 17552 11020 17604
rect 12900 17552 12952 17604
rect 13820 17552 13872 17604
rect 12072 17484 12124 17536
rect 15568 17552 15620 17604
rect 17316 17527 17368 17536
rect 17316 17493 17325 17527
rect 17325 17493 17359 17527
rect 17359 17493 17368 17527
rect 17316 17484 17368 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 2136 17280 2188 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 5264 17280 5316 17332
rect 6184 17280 6236 17332
rect 7012 17280 7064 17332
rect 8576 17280 8628 17332
rect 10324 17280 10376 17332
rect 10968 17280 11020 17332
rect 12532 17280 12584 17332
rect 13176 17280 13228 17332
rect 15752 17280 15804 17332
rect 16764 17323 16816 17332
rect 16764 17289 16773 17323
rect 16773 17289 16807 17323
rect 16807 17289 16816 17323
rect 16764 17280 16816 17289
rect 18236 17280 18288 17332
rect 18420 17280 18472 17332
rect 2596 17212 2648 17264
rect 3700 17212 3752 17264
rect 8208 17212 8260 17264
rect 3516 17144 3568 17196
rect 5448 17119 5500 17128
rect 5448 17085 5457 17119
rect 5457 17085 5491 17119
rect 5491 17085 5500 17119
rect 5448 17076 5500 17085
rect 8024 17144 8076 17196
rect 12072 17212 12124 17264
rect 15292 17212 15344 17264
rect 16580 17212 16632 17264
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 7656 17076 7708 17128
rect 8668 17119 8720 17128
rect 8668 17085 8677 17119
rect 8677 17085 8711 17119
rect 8711 17085 8720 17119
rect 8668 17076 8720 17085
rect 10784 17119 10836 17128
rect 10784 17085 10790 17119
rect 10790 17085 10836 17119
rect 10784 17076 10836 17085
rect 11244 17144 11296 17196
rect 18236 17144 18288 17196
rect 11612 17076 11664 17128
rect 3516 16940 3568 16992
rect 6736 17008 6788 17060
rect 7012 17008 7064 17060
rect 8576 17051 8628 17060
rect 8576 17017 8585 17051
rect 8585 17017 8619 17051
rect 8619 17017 8628 17051
rect 8576 17008 8628 17017
rect 10048 17008 10100 17060
rect 10600 17051 10652 17060
rect 10600 17017 10609 17051
rect 10609 17017 10643 17051
rect 10643 17017 10652 17051
rect 10600 17008 10652 17017
rect 11244 17008 11296 17060
rect 6828 16940 6880 16992
rect 7472 16940 7524 16992
rect 8760 16940 8812 16992
rect 12808 17076 12860 17128
rect 14648 17076 14700 17128
rect 16948 17119 17000 17128
rect 16948 17085 16957 17119
rect 16957 17085 16991 17119
rect 16991 17085 17000 17119
rect 16948 17076 17000 17085
rect 17316 17076 17368 17128
rect 18328 17076 18380 17128
rect 15476 17051 15528 17060
rect 12716 16940 12768 16992
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 15476 17017 15485 17051
rect 15485 17017 15519 17051
rect 15519 17017 15528 17051
rect 15476 17008 15528 17017
rect 13452 16940 13504 16949
rect 17224 17008 17276 17060
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 22100 17008 22152 17060
rect 19432 16940 19484 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3700 16736 3752 16788
rect 6184 16779 6236 16788
rect 6184 16745 6193 16779
rect 6193 16745 6227 16779
rect 6227 16745 6236 16779
rect 6184 16736 6236 16745
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 2780 16668 2832 16720
rect 3608 16668 3660 16720
rect 4160 16600 4212 16652
rect 6276 16600 6328 16652
rect 7748 16736 7800 16788
rect 7196 16668 7248 16720
rect 8300 16668 8352 16720
rect 9036 16668 9088 16720
rect 9404 16668 9456 16720
rect 10784 16711 10836 16720
rect 10784 16677 10793 16711
rect 10793 16677 10827 16711
rect 10827 16677 10836 16711
rect 10784 16668 10836 16677
rect 11244 16736 11296 16788
rect 12532 16736 12584 16788
rect 13544 16779 13596 16788
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 13636 16736 13688 16788
rect 14648 16779 14700 16788
rect 12716 16668 12768 16720
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 13820 16711 13872 16720
rect 13820 16677 13829 16711
rect 13829 16677 13863 16711
rect 13863 16677 13872 16711
rect 13820 16668 13872 16677
rect 17040 16668 17092 16720
rect 8024 16643 8076 16652
rect 8024 16609 8033 16643
rect 8033 16609 8067 16643
rect 8067 16609 8076 16643
rect 8024 16600 8076 16609
rect 8760 16600 8812 16652
rect 11704 16600 11756 16652
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15476 16600 15528 16652
rect 18788 16643 18840 16652
rect 18788 16609 18797 16643
rect 18797 16609 18831 16643
rect 18831 16609 18840 16643
rect 18788 16600 18840 16609
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 4528 16532 4580 16584
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 9312 16532 9364 16584
rect 10508 16532 10560 16584
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 14464 16532 14516 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 2320 16464 2372 16516
rect 3332 16464 3384 16516
rect 3608 16464 3660 16516
rect 9036 16464 9088 16516
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 4804 16396 4856 16448
rect 5448 16396 5500 16448
rect 8208 16396 8260 16448
rect 8760 16439 8812 16448
rect 8760 16405 8769 16439
rect 8769 16405 8803 16439
rect 8803 16405 8812 16439
rect 8760 16396 8812 16405
rect 9404 16396 9456 16448
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10784 16464 10836 16516
rect 11980 16464 12032 16516
rect 11612 16396 11664 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 4160 16192 4212 16244
rect 7656 16192 7708 16244
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 10508 16235 10560 16244
rect 8300 16192 8352 16201
rect 2872 16124 2924 16176
rect 6184 16167 6236 16176
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 6184 16133 6193 16167
rect 6193 16133 6227 16167
rect 6227 16133 6236 16167
rect 6184 16124 6236 16133
rect 7196 16124 7248 16176
rect 9036 16167 9088 16176
rect 9036 16133 9045 16167
rect 9045 16133 9079 16167
rect 9079 16133 9088 16167
rect 9036 16124 9088 16133
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 4804 16056 4856 16065
rect 8907 16099 8959 16108
rect 8907 16065 8916 16099
rect 8916 16065 8950 16099
rect 8950 16065 8959 16099
rect 10508 16201 10517 16235
rect 10517 16201 10551 16235
rect 10551 16201 10560 16235
rect 10508 16192 10560 16201
rect 15292 16192 15344 16244
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 18236 16235 18288 16244
rect 18236 16201 18245 16235
rect 18245 16201 18279 16235
rect 18279 16201 18288 16235
rect 18236 16192 18288 16201
rect 18788 16192 18840 16244
rect 13820 16124 13872 16176
rect 8907 16056 8959 16065
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 6000 15988 6052 16040
rect 1676 15963 1728 15972
rect 1676 15929 1685 15963
rect 1685 15929 1719 15963
rect 1719 15929 1728 15963
rect 1676 15920 1728 15929
rect 5908 15963 5960 15972
rect 2780 15895 2832 15904
rect 2780 15861 2789 15895
rect 2789 15861 2823 15895
rect 2823 15861 2832 15895
rect 2780 15852 2832 15861
rect 2964 15852 3016 15904
rect 5908 15929 5917 15963
rect 5917 15929 5951 15963
rect 5951 15929 5960 15963
rect 5908 15920 5960 15929
rect 7196 15988 7248 16040
rect 12716 16056 12768 16108
rect 16120 16124 16172 16176
rect 15292 16056 15344 16108
rect 16672 16056 16724 16108
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 8576 15963 8628 15972
rect 8576 15929 8585 15963
rect 8585 15929 8619 15963
rect 8619 15929 8628 15963
rect 8576 15920 8628 15929
rect 8760 15963 8812 15972
rect 8760 15929 8769 15963
rect 8769 15929 8803 15963
rect 8803 15929 8812 15963
rect 8760 15920 8812 15929
rect 9680 15920 9732 15972
rect 12440 15920 12492 15972
rect 13452 15920 13504 15972
rect 13544 15920 13596 15972
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 9956 15852 10008 15904
rect 12072 15852 12124 15904
rect 12992 15852 13044 15904
rect 16396 15920 16448 15972
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1492 15648 1544 15700
rect 4528 15648 4580 15700
rect 5908 15648 5960 15700
rect 2596 15623 2648 15632
rect 2596 15589 2605 15623
rect 2605 15589 2639 15623
rect 2639 15589 2648 15623
rect 2596 15580 2648 15589
rect 6092 15580 6144 15632
rect 6276 15580 6328 15632
rect 4620 15512 4672 15564
rect 8024 15648 8076 15700
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 8484 15648 8536 15700
rect 12716 15648 12768 15700
rect 13636 15648 13688 15700
rect 14740 15691 14792 15700
rect 14740 15657 14749 15691
rect 14749 15657 14783 15691
rect 14783 15657 14792 15691
rect 14740 15648 14792 15657
rect 6828 15580 6880 15632
rect 8944 15623 8996 15632
rect 8944 15589 8953 15623
rect 8953 15589 8987 15623
rect 8987 15589 8996 15623
rect 8944 15580 8996 15589
rect 9220 15580 9272 15632
rect 9404 15623 9456 15632
rect 9404 15589 9413 15623
rect 9413 15589 9447 15623
rect 9447 15589 9456 15623
rect 9404 15580 9456 15589
rect 9680 15623 9732 15632
rect 9680 15589 9689 15623
rect 9689 15589 9723 15623
rect 9723 15589 9732 15623
rect 9680 15580 9732 15589
rect 12808 15623 12860 15632
rect 12808 15589 12817 15623
rect 12817 15589 12851 15623
rect 12851 15589 12860 15623
rect 12808 15580 12860 15589
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 13820 15580 13872 15589
rect 16120 15623 16172 15632
rect 16120 15589 16129 15623
rect 16129 15589 16163 15623
rect 16163 15589 16172 15623
rect 16120 15580 16172 15589
rect 16948 15580 17000 15632
rect 17224 15580 17276 15632
rect 8300 15512 8352 15564
rect 8576 15512 8628 15564
rect 9036 15512 9088 15564
rect 10784 15555 10836 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 5540 15444 5592 15496
rect 6920 15444 6972 15496
rect 7196 15444 7248 15496
rect 10784 15521 10793 15555
rect 10793 15521 10827 15555
rect 10827 15521 10836 15555
rect 10784 15512 10836 15521
rect 11704 15512 11756 15564
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 17592 15512 17644 15521
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 12808 15444 12860 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 16396 15444 16448 15496
rect 2044 15308 2096 15360
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 2964 15308 3016 15360
rect 9220 15376 9272 15428
rect 4712 15308 4764 15360
rect 6276 15308 6328 15360
rect 7380 15308 7432 15360
rect 10140 15308 10192 15360
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 11704 15308 11756 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2504 15104 2556 15156
rect 3424 15104 3476 15156
rect 4344 15036 4396 15088
rect 112 14968 164 15020
rect 1584 14968 1636 15020
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 6000 15104 6052 15156
rect 6184 15104 6236 15156
rect 6828 15104 6880 15156
rect 8208 15104 8260 15156
rect 9404 15104 9456 15156
rect 12440 15104 12492 15156
rect 10140 15036 10192 15088
rect 10784 15036 10836 15088
rect 2044 14900 2096 14952
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 4068 14900 4120 14952
rect 4436 14832 4488 14884
rect 7196 14900 7248 14952
rect 7380 14943 7432 14952
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 8668 14832 8720 14884
rect 4712 14764 4764 14816
rect 6368 14764 6420 14816
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 6920 14764 6972 14773
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 11428 14968 11480 15020
rect 11336 14900 11388 14952
rect 13820 14968 13872 15020
rect 17592 15147 17644 15156
rect 17592 15113 17601 15147
rect 17601 15113 17635 15147
rect 17635 15113 17644 15147
rect 17592 15104 17644 15113
rect 16120 15036 16172 15088
rect 14648 14968 14700 15020
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 12808 14900 12860 14952
rect 15292 14900 15344 14952
rect 13176 14875 13228 14884
rect 13176 14841 13185 14875
rect 13185 14841 13219 14875
rect 13219 14841 13228 14875
rect 13176 14832 13228 14841
rect 10048 14764 10100 14816
rect 10692 14764 10744 14816
rect 11428 14807 11480 14816
rect 11428 14773 11437 14807
rect 11437 14773 11471 14807
rect 11471 14773 11480 14807
rect 11428 14764 11480 14773
rect 11704 14764 11756 14816
rect 13820 14764 13872 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 1768 14492 1820 14544
rect 2596 14492 2648 14544
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 8668 14560 8720 14612
rect 9220 14560 9272 14612
rect 9680 14560 9732 14612
rect 10784 14560 10836 14612
rect 11428 14560 11480 14612
rect 12532 14560 12584 14612
rect 12808 14560 12860 14612
rect 14648 14603 14700 14612
rect 14648 14569 14657 14603
rect 14657 14569 14691 14603
rect 14691 14569 14700 14603
rect 14648 14560 14700 14569
rect 16396 14603 16448 14612
rect 16396 14569 16405 14603
rect 16405 14569 16439 14603
rect 16439 14569 16448 14603
rect 16396 14560 16448 14569
rect 5540 14535 5592 14544
rect 5540 14501 5549 14535
rect 5549 14501 5583 14535
rect 5583 14501 5592 14535
rect 5540 14492 5592 14501
rect 6552 14535 6604 14544
rect 6552 14501 6555 14535
rect 6555 14501 6589 14535
rect 6589 14501 6604 14535
rect 6552 14492 6604 14501
rect 6828 14492 6880 14544
rect 7380 14492 7432 14544
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 6092 14424 6144 14476
rect 6920 14424 6972 14476
rect 8392 14424 8444 14476
rect 12348 14492 12400 14544
rect 12992 14492 13044 14544
rect 13636 14492 13688 14544
rect 16120 14492 16172 14544
rect 9404 14424 9456 14476
rect 9588 14424 9640 14476
rect 9956 14424 10008 14476
rect 10140 14424 10192 14476
rect 10876 14424 10928 14476
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 13176 14424 13228 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 3240 14356 3292 14408
rect 11704 14356 11756 14408
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 3792 14288 3844 14340
rect 5540 14288 5592 14340
rect 8944 14288 8996 14340
rect 9220 14288 9272 14340
rect 3148 14220 3200 14272
rect 5264 14263 5316 14272
rect 5264 14229 5273 14263
rect 5273 14229 5307 14263
rect 5307 14229 5316 14263
rect 5264 14220 5316 14229
rect 5448 14220 5500 14272
rect 11428 14288 11480 14340
rect 11612 14288 11664 14340
rect 11888 14288 11940 14340
rect 13728 14288 13780 14340
rect 21364 14288 21416 14340
rect 10600 14220 10652 14272
rect 11980 14220 12032 14272
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4712 14016 4764 14068
rect 6644 14016 6696 14068
rect 11980 14016 12032 14068
rect 12440 14016 12492 14068
rect 14372 14016 14424 14068
rect 15384 14016 15436 14068
rect 3332 13948 3384 14000
rect 8944 13948 8996 14000
rect 9128 13991 9180 14000
rect 9128 13957 9137 13991
rect 9137 13957 9171 13991
rect 9171 13957 9180 13991
rect 9128 13948 9180 13957
rect 9956 13991 10008 14000
rect 9956 13957 9965 13991
rect 9965 13957 9999 13991
rect 9999 13957 10008 13991
rect 9956 13948 10008 13957
rect 10600 13991 10652 14000
rect 10600 13957 10624 13991
rect 10624 13957 10652 13991
rect 10600 13948 10652 13957
rect 1400 13880 1452 13932
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 7380 13880 7432 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9680 13880 9732 13932
rect 5264 13812 5316 13864
rect 6828 13855 6880 13864
rect 1676 13787 1728 13796
rect 1676 13753 1685 13787
rect 1685 13753 1719 13787
rect 1719 13753 1728 13787
rect 1676 13744 1728 13753
rect 2412 13744 2464 13796
rect 3148 13787 3200 13796
rect 1308 13676 1360 13728
rect 3148 13753 3157 13787
rect 3157 13753 3191 13787
rect 3191 13753 3200 13787
rect 3148 13744 3200 13753
rect 3240 13787 3292 13796
rect 3240 13753 3249 13787
rect 3249 13753 3283 13787
rect 3283 13753 3292 13787
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 10048 13812 10100 13864
rect 3240 13744 3292 13753
rect 6644 13744 6696 13796
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 6000 13676 6052 13728
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 9128 13744 9180 13796
rect 10968 13948 11020 14000
rect 15752 13991 15804 14000
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 15752 13948 15804 13957
rect 16948 13948 17000 14000
rect 6552 13676 6604 13685
rect 6828 13676 6880 13728
rect 7288 13676 7340 13728
rect 8024 13676 8076 13728
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 15476 13880 15528 13932
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 11612 13744 11664 13796
rect 13636 13744 13688 13796
rect 15200 13787 15252 13796
rect 15200 13753 15209 13787
rect 15209 13753 15243 13787
rect 15243 13753 15252 13787
rect 15200 13744 15252 13753
rect 15384 13744 15436 13796
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 13820 13676 13872 13728
rect 16120 13719 16172 13728
rect 16120 13685 16129 13719
rect 16129 13685 16163 13719
rect 16163 13685 16172 13719
rect 16120 13676 16172 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2596 13515 2648 13524
rect 2596 13481 2605 13515
rect 2605 13481 2639 13515
rect 2639 13481 2648 13515
rect 2596 13472 2648 13481
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 6184 13472 6236 13524
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 9220 13472 9272 13524
rect 9864 13472 9916 13524
rect 9956 13472 10008 13524
rect 10968 13472 11020 13524
rect 13452 13515 13504 13524
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 3332 13404 3384 13456
rect 4436 13447 4488 13456
rect 4436 13413 4445 13447
rect 4445 13413 4479 13447
rect 4479 13413 4488 13447
rect 4436 13404 4488 13413
rect 6368 13336 6420 13388
rect 9404 13404 9456 13456
rect 12808 13404 12860 13456
rect 13728 13404 13780 13456
rect 14832 13404 14884 13456
rect 15200 13404 15252 13456
rect 16120 13404 16172 13456
rect 6644 13379 6696 13388
rect 6644 13345 6653 13379
rect 6653 13345 6687 13379
rect 6687 13345 6696 13379
rect 6644 13336 6696 13345
rect 8116 13379 8168 13388
rect 8116 13345 8125 13379
rect 8125 13345 8159 13379
rect 8159 13345 8168 13379
rect 8116 13336 8168 13345
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 9496 13336 9548 13388
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 11704 13336 11756 13388
rect 12348 13379 12400 13388
rect 12348 13345 12357 13379
rect 12357 13345 12391 13379
rect 12391 13345 12400 13379
rect 12348 13336 12400 13345
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 1952 13311 2004 13320
rect 1952 13277 1961 13311
rect 1961 13277 1995 13311
rect 1995 13277 2004 13311
rect 1952 13268 2004 13277
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 4344 13268 4396 13277
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 13544 13268 13596 13320
rect 8300 13200 8352 13252
rect 1768 13132 1820 13184
rect 4252 13132 4304 13184
rect 6920 13132 6972 13184
rect 7380 13132 7432 13184
rect 8392 13132 8444 13184
rect 9036 13200 9088 13252
rect 11060 13200 11112 13252
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 3332 12928 3384 12980
rect 6368 12928 6420 12980
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 10968 12928 11020 12980
rect 11244 12971 11296 12980
rect 11244 12937 11253 12971
rect 11253 12937 11287 12971
rect 11287 12937 11296 12971
rect 11244 12928 11296 12937
rect 11704 12928 11756 12980
rect 13728 12928 13780 12980
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 3056 12860 3108 12912
rect 4436 12860 4488 12912
rect 3976 12792 4028 12844
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 4620 12792 4672 12844
rect 5080 12792 5132 12844
rect 6184 12792 6236 12844
rect 8668 12835 8720 12844
rect 6920 12724 6972 12776
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 11428 12792 11480 12844
rect 7748 12724 7800 12776
rect 8576 12724 8628 12776
rect 8760 12724 8812 12776
rect 1952 12656 2004 12708
rect 3516 12699 3568 12708
rect 3516 12665 3525 12699
rect 3525 12665 3559 12699
rect 3559 12665 3568 12699
rect 3516 12656 3568 12665
rect 7840 12699 7892 12708
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 7840 12665 7849 12699
rect 7849 12665 7883 12699
rect 7883 12665 7892 12699
rect 7840 12656 7892 12665
rect 3240 12588 3292 12597
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 7932 12588 7984 12640
rect 9864 12724 9916 12776
rect 10140 12656 10192 12708
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 9956 12588 10008 12597
rect 12072 12724 12124 12776
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 11152 12588 11204 12640
rect 13084 12588 13136 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 1676 12384 1728 12436
rect 3516 12427 3568 12436
rect 3516 12393 3525 12427
rect 3525 12393 3559 12427
rect 3559 12393 3568 12427
rect 3516 12384 3568 12393
rect 4344 12384 4396 12436
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 6644 12427 6696 12436
rect 6644 12393 6653 12427
rect 6653 12393 6687 12427
rect 6687 12393 6696 12427
rect 6644 12384 6696 12393
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 8668 12384 8720 12436
rect 10968 12384 11020 12436
rect 11796 12384 11848 12436
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 13820 12427 13872 12436
rect 13820 12393 13829 12427
rect 13829 12393 13863 12427
rect 13863 12393 13872 12427
rect 13820 12384 13872 12393
rect 3240 12316 3292 12368
rect 5356 12316 5408 12368
rect 6000 12316 6052 12368
rect 6184 12316 6236 12368
rect 7932 12316 7984 12368
rect 9772 12316 9824 12368
rect 10784 12316 10836 12368
rect 11520 12316 11572 12368
rect 13268 12316 13320 12368
rect 3056 12291 3108 12300
rect 3056 12257 3065 12291
rect 3065 12257 3099 12291
rect 3099 12257 3108 12291
rect 3056 12248 3108 12257
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 9588 12180 9640 12232
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10968 12180 11020 12232
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 8484 12112 8536 12164
rect 9956 12112 10008 12164
rect 11152 12112 11204 12164
rect 13544 12112 13596 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 6368 12087 6420 12096
rect 6368 12053 6377 12087
rect 6377 12053 6411 12087
rect 6411 12053 6420 12087
rect 6368 12044 6420 12053
rect 6920 12044 6972 12096
rect 8760 12087 8812 12096
rect 8760 12053 8769 12087
rect 8769 12053 8803 12087
rect 8803 12053 8812 12087
rect 8760 12044 8812 12053
rect 9772 12044 9824 12096
rect 10140 12044 10192 12096
rect 11336 12044 11388 12096
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1952 11883 2004 11892
rect 1952 11849 1961 11883
rect 1961 11849 1995 11883
rect 1995 11849 2004 11883
rect 1952 11840 2004 11849
rect 3056 11840 3108 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 7932 11883 7984 11892
rect 6184 11840 6236 11849
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 10876 11840 10928 11892
rect 3424 11704 3476 11756
rect 4344 11704 4396 11756
rect 9588 11772 9640 11824
rect 11336 11772 11388 11824
rect 12992 11772 13044 11824
rect 8484 11747 8536 11756
rect 8484 11713 8493 11747
rect 8493 11713 8527 11747
rect 8527 11713 8536 11747
rect 8484 11704 8536 11713
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 1676 11636 1728 11688
rect 2596 11636 2648 11688
rect 11060 11636 11112 11688
rect 11520 11636 11572 11688
rect 17960 11636 18012 11688
rect 3700 11611 3752 11620
rect 3700 11577 3702 11611
rect 3702 11577 3736 11611
rect 3736 11577 3752 11611
rect 3700 11568 3752 11577
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 4988 11543 5040 11552
rect 4988 11509 4997 11543
rect 4997 11509 5031 11543
rect 5031 11509 5040 11543
rect 6368 11568 6420 11620
rect 8208 11611 8260 11620
rect 8208 11577 8217 11611
rect 8217 11577 8251 11611
rect 8251 11577 8260 11611
rect 8208 11568 8260 11577
rect 8668 11568 8720 11620
rect 9864 11611 9916 11620
rect 9864 11577 9873 11611
rect 9873 11577 9907 11611
rect 9907 11577 9916 11611
rect 9864 11568 9916 11577
rect 4988 11500 5040 11509
rect 9680 11500 9732 11552
rect 10968 11500 11020 11552
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2780 11296 2832 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 7748 11296 7800 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 3700 11228 3752 11280
rect 7840 11228 7892 11280
rect 8484 11271 8536 11280
rect 8484 11237 8493 11271
rect 8493 11237 8527 11271
rect 8527 11237 8536 11271
rect 8484 11228 8536 11237
rect 9680 11271 9732 11280
rect 9680 11237 9689 11271
rect 9689 11237 9723 11271
rect 9723 11237 9732 11271
rect 9680 11228 9732 11237
rect 2780 11160 2832 11212
rect 3332 11160 3384 11212
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 9864 11296 9916 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 1676 11092 1728 11144
rect 4896 11092 4948 11144
rect 7656 11092 7708 11144
rect 8208 11024 8260 11076
rect 3424 10956 3476 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2320 10752 2372 10804
rect 2044 10684 2096 10736
rect 4160 10752 4212 10804
rect 4988 10752 5040 10804
rect 5540 10752 5592 10804
rect 8760 10752 8812 10804
rect 9772 10752 9824 10804
rect 9864 10752 9916 10804
rect 10692 10752 10744 10804
rect 2780 10616 2832 10668
rect 1952 10548 2004 10600
rect 2504 10591 2556 10600
rect 2504 10557 2548 10591
rect 2548 10557 2556 10591
rect 2504 10548 2556 10557
rect 7656 10684 7708 10736
rect 4160 10616 4212 10668
rect 6736 10616 6788 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 5172 10548 5224 10600
rect 8760 10548 8812 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10968 10548 11020 10600
rect 112 10412 164 10464
rect 15384 10412 15436 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2688 10208 2740 10260
rect 3516 10208 3568 10260
rect 7656 10208 7708 10260
rect 3148 10140 3200 10192
rect 2320 10072 2372 10124
rect 2964 10072 3016 10124
rect 3884 10072 3936 10124
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 8024 10072 8076 10124
rect 2044 10004 2096 10056
rect 3056 10004 3108 10056
rect 8392 10004 8444 10056
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 2688 9868 2740 9920
rect 8300 9868 8352 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1308 9664 1360 9716
rect 2320 9707 2372 9716
rect 2320 9673 2329 9707
rect 2329 9673 2363 9707
rect 2363 9673 2372 9707
rect 2320 9664 2372 9673
rect 3424 9664 3476 9716
rect 3608 9707 3660 9716
rect 3608 9673 3617 9707
rect 3617 9673 3651 9707
rect 3651 9673 3660 9707
rect 3608 9664 3660 9673
rect 3884 9664 3936 9716
rect 2136 9596 2188 9648
rect 3976 9596 4028 9648
rect 112 9528 164 9580
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 7564 9460 7616 9512
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 7748 9367 7800 9376
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 8024 9324 8076 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9120 1728 9172
rect 1952 9120 2004 9172
rect 7748 9052 7800 9104
rect 9404 9052 9456 9104
rect 112 8984 164 9036
rect 1860 8984 1912 9036
rect 2044 8984 2096 9036
rect 3240 8984 3292 9036
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 1952 8848 2004 8900
rect 7104 8848 7156 8900
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1860 8619 1912 8628
rect 1860 8585 1869 8619
rect 1869 8585 1903 8619
rect 1903 8585 1912 8619
rect 1860 8576 1912 8585
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 1768 8508 1820 8560
rect 2412 8508 2464 8560
rect 7748 8576 7800 8628
rect 10048 8508 10100 8560
rect 2228 8372 2280 8424
rect 2447 8415 2499 8424
rect 2447 8381 2456 8415
rect 2456 8381 2490 8415
rect 2490 8381 2499 8415
rect 2447 8372 2499 8381
rect 8024 8236 8076 8288
rect 8484 8236 8536 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 1676 7760 1728 7812
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 112 7488 164 7540
rect 1400 7488 1452 7540
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 12532 6740 12584 6792
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 112 6400 164 6452
rect 1400 6400 1452 6452
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 112 5720 164 5772
rect 1400 5763 1452 5772
rect 1400 5729 1444 5763
rect 1444 5729 1452 5763
rect 1400 5720 1452 5729
rect 12900 5652 12952 5704
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1400 5312 1452 5364
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 112 4632 164 4684
rect 1400 4675 1452 4684
rect 1400 4641 1444 4675
rect 1444 4641 1452 4675
rect 1400 4632 1452 4641
rect 13176 4564 13228 4616
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1400 4224 1452 4276
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 112 3544 164 3596
rect 2228 3544 2280 3596
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 1308 2932 1360 2984
rect 1400 2796 1452 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 6276 2592 6328 2644
rect 1216 2456 1268 2508
rect 2136 2456 2188 2508
rect 11152 2388 11204 2440
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 4160 76 4212 128
rect 5264 76 5316 128
rect 11060 76 11112 128
rect 12256 76 12308 128
rect 17960 76 18012 128
rect 19248 76 19300 128
<< metal2 >>
rect 478 27520 534 28000
rect 1490 27520 1546 28000
rect 2502 27520 2558 28000
rect 3514 27520 3570 28000
rect 4618 27568 4674 28000
rect 112 25492 164 25498
rect 112 25434 164 25440
rect 124 25401 152 25434
rect 110 25392 166 25401
rect 110 25327 166 25336
rect 492 22001 520 27520
rect 1504 26178 1532 27520
rect 2516 26246 2544 27520
rect 3146 26888 3202 26897
rect 3146 26823 3202 26832
rect 2504 26240 2556 26246
rect 2504 26182 2556 26188
rect 1492 26172 1544 26178
rect 1492 26114 1544 26120
rect 2872 25424 2924 25430
rect 2872 25366 2924 25372
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 1412 24818 1440 25230
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1952 24812 2004 24818
rect 1952 24754 2004 24760
rect 1964 24410 1992 24754
rect 2228 24676 2280 24682
rect 2228 24618 2280 24624
rect 1952 24404 2004 24410
rect 1952 24346 2004 24352
rect 2136 24132 2188 24138
rect 2136 24074 2188 24080
rect 2148 23730 2176 24074
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 1768 23588 1820 23594
rect 1768 23530 1820 23536
rect 1780 23474 1808 23530
rect 1688 23446 1808 23474
rect 1688 22982 1716 23446
rect 1872 22982 1900 23666
rect 2240 23322 2268 24618
rect 2320 24336 2372 24342
rect 2320 24278 2372 24284
rect 2332 23866 2360 24278
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2320 23724 2372 23730
rect 2320 23666 2372 23672
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1688 22166 1716 22918
rect 2332 22642 2360 23666
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2320 22500 2372 22506
rect 2320 22442 2372 22448
rect 1676 22160 1728 22166
rect 1676 22102 1728 22108
rect 2332 22098 2360 22442
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 478 21992 534 22001
rect 478 21927 534 21936
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1768 21616 1820 21622
rect 1768 21558 1820 21564
rect 1780 21146 1808 21558
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1582 20632 1638 20641
rect 1582 20567 1638 20576
rect 110 20088 166 20097
rect 110 20023 166 20032
rect 124 15026 152 20023
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18154 1532 18566
rect 1492 18148 1544 18154
rect 1492 18090 1544 18096
rect 1504 15706 1532 18090
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1596 15162 1624 20567
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1688 19378 1716 19926
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1688 17542 1716 18090
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17338 1716 17478
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 16046 1808 16390
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 112 15020 164 15026
rect 112 14962 164 14968
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1308 13728 1360 13734
rect 1308 13670 1360 13676
rect 110 10840 166 10849
rect 110 10775 166 10784
rect 124 10470 152 10775
rect 112 10464 164 10470
rect 112 10406 164 10412
rect 110 9752 166 9761
rect 1320 9722 1348 13670
rect 1412 12442 1440 13874
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1596 10810 1624 14962
rect 1688 14618 1716 15914
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1688 13802 1716 14554
rect 1780 14550 1808 15982
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1676 13320 1728 13326
rect 1872 13308 1900 21898
rect 2332 21622 2360 22034
rect 2320 21616 2372 21622
rect 2320 21558 2372 21564
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 2240 20058 2268 21354
rect 2332 21146 2360 21354
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2056 19446 2084 19858
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 2056 19242 2084 19382
rect 2044 19236 2096 19242
rect 2044 19178 2096 19184
rect 2056 18970 2084 19178
rect 2148 18970 2176 19790
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2240 18698 2268 19178
rect 2424 18902 2452 25230
rect 2516 24614 2544 25298
rect 2596 24676 2648 24682
rect 2596 24618 2648 24624
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2412 18896 2464 18902
rect 2412 18838 2464 18844
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2424 18426 2452 18838
rect 2516 18426 2544 24550
rect 2608 24206 2636 24618
rect 2596 24200 2648 24206
rect 2648 24160 2820 24188
rect 2596 24142 2648 24148
rect 2686 23896 2742 23905
rect 2596 23860 2648 23866
rect 2686 23831 2742 23840
rect 2596 23802 2648 23808
rect 2608 23186 2636 23802
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2608 22778 2636 23122
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2700 21690 2728 23831
rect 2792 22545 2820 24160
rect 2884 22710 2912 25366
rect 3056 25152 3108 25158
rect 3056 25094 3108 25100
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 2976 23497 3004 23530
rect 2962 23488 3018 23497
rect 2962 23423 3018 23432
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2778 22536 2834 22545
rect 2778 22471 2834 22480
rect 2884 22234 2912 22646
rect 2872 22228 2924 22234
rect 2872 22170 2924 22176
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2884 20913 2912 21354
rect 2870 20904 2926 20913
rect 2870 20839 2926 20848
rect 2884 20466 2912 20839
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2136 17808 2188 17814
rect 2136 17750 2188 17756
rect 2148 17338 2176 17750
rect 2700 17678 2728 18090
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2226 17504 2282 17513
rect 2226 17439 2282 17448
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2134 16552 2190 16561
rect 2134 16487 2190 16496
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 2056 14958 2084 15302
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 13326 1992 14350
rect 1728 13280 1900 13308
rect 1952 13320 2004 13326
rect 1676 13262 1728 13268
rect 1952 13262 2004 13268
rect 1688 12442 1716 13262
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1688 11354 1716 11630
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 110 9687 166 9696
rect 1308 9716 1360 9722
rect 124 9586 152 9687
rect 1308 9658 1360 9664
rect 112 9580 164 9586
rect 112 9522 164 9528
rect 1688 9178 1716 11086
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 112 9036 164 9042
rect 112 8978 164 8984
rect 124 8809 152 8978
rect 1674 8936 1730 8945
rect 1674 8871 1730 8880
rect 110 8800 166 8809
rect 110 8735 166 8744
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 110 7712 166 7721
rect 110 7647 166 7656
rect 124 7546 152 7647
rect 1412 7546 1440 7890
rect 1688 7818 1716 8871
rect 1780 8566 1808 13126
rect 1964 12850 1992 13262
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1858 12336 1914 12345
rect 1858 12271 1914 12280
rect 1872 9518 1900 12271
rect 1964 12102 1992 12650
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11898 1992 12038
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2056 10742 2084 14894
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9926 1992 10542
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1964 9178 1992 9862
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2056 9042 2084 9998
rect 2148 9654 2176 16487
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1872 8634 1900 8978
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 112 7540 164 7546
rect 112 7482 164 7488
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 110 6624 166 6633
rect 110 6559 166 6568
rect 124 6458 152 6559
rect 1412 6458 1440 6802
rect 112 6452 164 6458
rect 112 6394 164 6400
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 112 5772 164 5778
rect 112 5714 164 5720
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 124 5681 152 5714
rect 110 5672 166 5681
rect 110 5607 166 5616
rect 1412 5370 1440 5714
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 112 4684 164 4690
rect 112 4626 164 4632
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 124 4593 152 4626
rect 110 4584 166 4593
rect 110 4519 166 4528
rect 1412 4282 1440 4626
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1596 3738 1624 6151
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 112 3596 164 3602
rect 112 3538 164 3544
rect 124 3505 152 3538
rect 110 3496 166 3505
rect 110 3431 166 3440
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1398 2952 1454 2961
rect 1320 2825 1348 2926
rect 1398 2887 1454 2896
rect 1412 2854 1440 2887
rect 1400 2848 1452 2854
rect 1306 2816 1362 2825
rect 1400 2790 1452 2796
rect 1306 2751 1362 2760
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1228 2009 1256 2450
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1766 82 1822 480
rect 1964 82 1992 8842
rect 2240 8634 2268 17439
rect 2516 17252 2544 17614
rect 2884 17524 2912 20266
rect 3068 19990 3096 25094
rect 3160 23322 3188 26823
rect 3148 23316 3200 23322
rect 3148 23258 3200 23264
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 3148 20528 3200 20534
rect 3148 20470 3200 20476
rect 3160 20262 3188 20470
rect 3252 20466 3280 20946
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3056 19984 3108 19990
rect 3056 19926 3108 19932
rect 3160 18698 3188 20198
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3160 18193 3188 18226
rect 3146 18184 3202 18193
rect 3146 18119 3202 18128
rect 3160 17882 3188 18119
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3252 17762 3280 19722
rect 3160 17734 3280 17762
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2700 17496 2912 17524
rect 2596 17264 2648 17270
rect 2516 17224 2596 17252
rect 2516 16590 2544 17224
rect 2596 17206 2648 17212
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 15366 2360 16458
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 10810 2360 15302
rect 2516 15162 2544 15438
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2608 15026 2636 15574
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 13802 2452 14350
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2332 9722 2360 10066
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2240 8430 2268 8570
rect 2424 8566 2452 13738
rect 2502 13696 2558 13705
rect 2502 13631 2558 13640
rect 2516 10606 2544 13631
rect 2608 13530 2636 14486
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2608 11694 2636 12922
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2700 10266 2728 17496
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2792 15910 2820 16662
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 11354 2820 15846
rect 2884 15502 2912 16118
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2780 11348 2832 11354
rect 2884 11336 2912 15438
rect 2976 15366 3004 15846
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2976 14958 3004 15302
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2976 14618 3004 14894
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3068 14498 3096 17614
rect 2976 14470 3096 14498
rect 2976 11506 3004 14470
rect 3160 14396 3188 17734
rect 3344 16522 3372 22918
rect 3528 22409 3556 27520
rect 5630 27554 5686 28000
rect 4618 27503 4674 27512
rect 5460 27526 5686 27554
rect 4632 27443 4660 27503
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5184 24954 5212 25230
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 4252 24744 4304 24750
rect 4252 24686 4304 24692
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 23866 3924 24550
rect 4264 24342 4292 24686
rect 5184 24614 5212 24890
rect 5356 24880 5408 24886
rect 5356 24822 5408 24828
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 4344 24404 4396 24410
rect 4344 24346 4396 24352
rect 4252 24336 4304 24342
rect 4252 24278 4304 24284
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3896 23526 3924 23802
rect 4172 23730 4200 24142
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3608 23112 3660 23118
rect 4172 23089 4200 23666
rect 3608 23054 3660 23060
rect 4158 23080 4214 23089
rect 3620 22506 3648 23054
rect 4158 23015 4214 23024
rect 4250 22672 4306 22681
rect 4250 22607 4306 22616
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3608 22500 3660 22506
rect 3608 22442 3660 22448
rect 3514 22400 3570 22409
rect 3514 22335 3570 22344
rect 3620 21894 3648 22442
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 19378 3464 19654
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3436 18902 3464 19314
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3436 18290 3464 18838
rect 3528 18630 3556 19382
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17202 3556 17478
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3528 17105 3556 17138
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16114 3464 16390
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3436 15162 3464 16050
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3068 14368 3188 14396
rect 3240 14408 3292 14414
rect 3068 13002 3096 14368
rect 3240 14350 3292 14356
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3160 13802 3188 14214
rect 3252 13802 3280 14350
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3344 13462 3372 13942
rect 3436 13938 3464 15098
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3528 13814 3556 16934
rect 3620 16726 3648 21830
rect 3712 21078 3740 22510
rect 3882 21720 3938 21729
rect 3882 21655 3938 21664
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3804 19786 3832 20878
rect 3896 20602 3924 21655
rect 4264 21146 4292 22607
rect 4252 21140 4304 21146
rect 4252 21082 4304 21088
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 4356 19990 4384 24346
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4632 23730 4660 24142
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 5000 23526 5028 24278
rect 5276 24070 5304 24618
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 4540 22438 4568 23122
rect 4896 22704 4948 22710
rect 4896 22646 4948 22652
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4540 21049 4568 22374
rect 4816 22030 4844 22510
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4816 21690 4844 21966
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4526 21040 4582 21049
rect 4526 20975 4582 20984
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 3792 19780 3844 19786
rect 3792 19722 3844 19728
rect 4356 19514 4384 19926
rect 4528 19848 4580 19854
rect 4816 19825 4844 19926
rect 4528 19790 4580 19796
rect 4802 19816 4858 19825
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4540 19378 4568 19790
rect 4802 19751 4858 19760
rect 4816 19446 4844 19751
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4252 18896 4304 18902
rect 4066 18864 4122 18873
rect 4252 18838 4304 18844
rect 4066 18799 4122 18808
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3712 16794 3740 17206
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 16720 3660 16726
rect 3608 16662 3660 16668
rect 3608 16516 3660 16522
rect 3608 16458 3660 16464
rect 3436 13786 3556 13814
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3068 12974 3188 13002
rect 3344 12986 3372 13398
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 3068 12306 3096 12854
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 11898 3096 12242
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2976 11478 3096 11506
rect 2884 11308 3004 11336
rect 2780 11290 2832 11296
rect 2870 11248 2926 11257
rect 2780 11212 2832 11218
rect 2870 11183 2926 11192
rect 2780 11154 2832 11160
rect 2792 10674 2820 11154
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 8634 2728 9862
rect 2884 9518 2912 11183
rect 2976 10130 3004 11308
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 3068 10062 3096 11478
rect 3160 10198 3188 12974
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3252 12374 3280 12582
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3436 11880 3464 13786
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3528 12442 3556 12650
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3514 12064 3570 12073
rect 3514 11999 3570 12008
rect 3344 11852 3464 11880
rect 3344 11218 3372 11852
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3436 11014 3464 11698
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3436 9722 3464 10950
rect 3528 10266 3556 11999
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3620 9722 3648 16458
rect 3804 14346 3832 18702
rect 3882 15464 3938 15473
rect 3882 15399 3938 15408
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3712 11286 3740 11562
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3896 10130 3924 15399
rect 4080 14958 4108 18799
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 17762 4200 18702
rect 4264 18426 4292 18838
rect 4816 18426 4844 19110
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4724 17882 4752 18158
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4172 17734 4292 17762
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4172 17338 4200 17614
rect 4264 17542 4292 17734
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16250 4200 16594
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4264 13190 4292 17478
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4540 15745 4568 16526
rect 4526 15736 4582 15745
rect 4526 15671 4528 15680
rect 4580 15671 4582 15680
rect 4528 15642 4580 15648
rect 4540 15611 4568 15642
rect 4632 15570 4660 16526
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 16114 4844 16390
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4356 14872 4384 15030
rect 4436 14884 4488 14890
rect 4356 14844 4436 14872
rect 4436 14826 4488 14832
rect 4724 14822 4752 15302
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 14482 4752 14758
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 14074 4752 14418
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 9722 3924 10066
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 9654 4016 12786
rect 4172 10810 4200 12786
rect 4356 12442 4384 13262
rect 4448 12918 4476 13398
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4632 12850 4660 13262
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4356 11762 4384 12378
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4618 11656 4674 11665
rect 4618 11591 4674 11600
rect 4632 11558 4660 11591
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4908 11150 4936 22646
rect 5000 22234 5028 23462
rect 5080 22976 5132 22982
rect 5080 22918 5132 22924
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 5092 22574 5120 22918
rect 5276 22778 5304 22918
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5092 22148 5120 22374
rect 5166 22160 5218 22166
rect 5092 22120 5166 22148
rect 5092 21418 5120 22120
rect 5166 22102 5218 22108
rect 5368 21962 5396 24822
rect 5460 23769 5488 27526
rect 5630 27520 5686 27526
rect 6642 27520 6698 28000
rect 7654 27520 7710 28000
rect 8758 27520 8814 28000
rect 9770 27520 9826 28000
rect 10782 27520 10838 28000
rect 11794 27520 11850 28000
rect 12898 27520 12954 28000
rect 13910 27520 13966 28000
rect 14922 27554 14978 28000
rect 15934 27554 15990 28000
rect 14844 27526 14978 27554
rect 5538 25800 5594 25809
rect 5538 25735 5594 25744
rect 5552 23866 5580 25735
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6104 24818 6132 25298
rect 6092 24812 6144 24818
rect 6092 24754 6144 24760
rect 6104 24342 6132 24754
rect 6552 24744 6604 24750
rect 6552 24686 6604 24692
rect 6460 24676 6512 24682
rect 6460 24618 6512 24624
rect 6472 24342 6500 24618
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6460 24336 6512 24342
rect 6460 24278 6512 24284
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5446 23760 5502 23769
rect 5446 23695 5502 23704
rect 6104 23526 6132 24278
rect 6368 24200 6420 24206
rect 6472 24177 6500 24278
rect 6368 24142 6420 24148
rect 6458 24168 6514 24177
rect 6380 23866 6408 24142
rect 6458 24103 6514 24112
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 5448 22500 5500 22506
rect 5448 22442 5500 22448
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 5080 21072 5132 21078
rect 5080 21014 5132 21020
rect 5092 19990 5120 21014
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 5184 20398 5212 20946
rect 5460 20806 5488 22442
rect 5552 22137 5580 23462
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5538 22128 5594 22137
rect 5538 22063 5594 22072
rect 6012 21894 6040 23054
rect 6104 22778 6132 23462
rect 6276 23248 6328 23254
rect 6276 23190 6328 23196
rect 6092 22772 6144 22778
rect 6092 22714 6144 22720
rect 6288 22438 6316 23190
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6288 22166 6316 22374
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5644 21146 5672 21422
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5460 20398 5488 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20602 6040 21830
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5908 20392 5960 20398
rect 6104 20380 6132 20946
rect 6288 20602 6316 21014
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 5960 20352 6132 20380
rect 5908 20334 5960 20340
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5092 19310 5120 19926
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19310 5212 19654
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5092 18970 5120 19246
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 5000 17882 5028 18090
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5184 17678 5212 19110
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5276 18086 5304 18294
rect 5460 18086 5488 20334
rect 5920 19854 5948 20334
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 18834 6040 19994
rect 6380 19990 6408 20946
rect 6472 20466 6500 22102
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 19310 6132 19858
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5276 17814 5304 18022
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5276 17338 5304 17750
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5460 17134 5488 18022
rect 6012 17882 6040 18770
rect 6196 18358 6224 18838
rect 6564 18426 6592 24686
rect 6656 22681 6684 27520
rect 7668 24721 7696 27520
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7654 24712 7710 24721
rect 6828 24676 6880 24682
rect 7654 24647 7710 24656
rect 6828 24618 6880 24624
rect 6840 24410 6868 24618
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6642 22672 6698 22681
rect 6642 22607 6698 22616
rect 6840 21554 6868 24006
rect 7760 23594 7788 25230
rect 8312 24614 8340 25298
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8300 24608 8352 24614
rect 8300 24550 8352 24556
rect 8312 24342 8340 24550
rect 8300 24336 8352 24342
rect 8300 24278 8352 24284
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7208 22574 7236 22986
rect 7392 22982 7420 23530
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6656 21457 6684 21490
rect 6642 21448 6698 21457
rect 6642 21383 6698 21392
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20398 6960 20742
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6656 18902 6684 20266
rect 6932 19174 6960 20334
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7116 19334 7144 19858
rect 7116 19306 7236 19334
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 7024 18290 7052 18566
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6564 18086 6592 18226
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5460 16454 5488 17070
rect 6196 16794 6224 17274
rect 7024 17066 7052 17274
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 6748 16794 6776 17002
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 16046 5488 16390
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6196 16182 6224 16730
rect 6840 16674 6868 16934
rect 7208 16833 7236 19306
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7300 18222 7328 19110
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7300 17610 7328 18158
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7194 16824 7250 16833
rect 7194 16759 7250 16768
rect 7208 16726 7236 16759
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6748 16646 6868 16674
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 5170 14376 5226 14385
rect 5170 14311 5226 14320
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5092 12442 5120 12786
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5000 11218 5028 11494
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 5000 10810 5028 11154
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3252 8634 3280 8978
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2424 8430 2452 8502
rect 2228 8424 2280 8430
rect 2424 8424 2499 8430
rect 2424 8384 2447 8424
rect 2228 8366 2280 8372
rect 2447 8366 2499 8372
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2240 3194 2268 3538
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2148 1057 2176 2450
rect 2134 1048 2190 1057
rect 2134 983 2190 992
rect 4172 134 4200 10610
rect 5184 10606 5212 14311
rect 5460 14278 5488 15982
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5920 15706 5948 15914
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 14550 5580 15438
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15162 6040 15982
rect 6092 15632 6144 15638
rect 6196 15620 6224 16118
rect 6288 15638 6316 16594
rect 6144 15592 6224 15620
rect 6092 15574 6144 15580
rect 6196 15162 6224 15592
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5276 13870 5304 14214
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 12374 5396 12582
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5460 12306 5488 13670
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5460 11354 5488 12242
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 10810 5580 14282
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12374 6040 13670
rect 6104 13530 6132 14418
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6196 12850 6224 13466
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6196 11898 6224 12310
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6288 2650 6316 15302
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 13394 6408 14758
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6564 13734 6592 14486
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6656 13802 6684 14010
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6656 13394 6684 13738
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6380 12986 6408 13330
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6656 12442 6684 13330
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 11626 6408 12038
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6748 11218 6776 16646
rect 7208 16182 7236 16662
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7208 16046 7236 16118
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6840 15162 6868 15574
rect 6932 15502 6960 15846
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6840 14550 6868 15098
rect 7208 14958 7236 15438
rect 7392 15366 7420 22918
rect 7944 22234 7972 23462
rect 8128 23118 8156 23666
rect 8208 23248 8260 23254
rect 8208 23190 8260 23196
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8220 22778 8248 23190
rect 8312 22982 8340 24278
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8404 23730 8432 24142
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8496 23254 8524 24686
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8484 23248 8536 23254
rect 8484 23190 8536 23196
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7944 21350 7972 21966
rect 8036 21690 8064 22102
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 8588 21593 8616 24074
rect 8772 23225 8800 27520
rect 9784 24818 9812 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10796 25514 10824 27520
rect 10796 25486 11008 25514
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9876 24954 9904 25298
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8864 23866 8892 24550
rect 9876 24342 9904 24890
rect 9864 24336 9916 24342
rect 9864 24278 9916 24284
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8864 23526 8892 23802
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9232 23633 9260 23666
rect 9218 23624 9274 23633
rect 9218 23559 9274 23568
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 9232 23254 9260 23559
rect 9220 23248 9272 23254
rect 8758 23216 8814 23225
rect 9220 23190 9272 23196
rect 8758 23151 8814 23160
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 8944 23044 8996 23050
rect 8944 22986 8996 22992
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8772 22234 8800 22918
rect 8956 22545 8984 22986
rect 9600 22778 9628 23054
rect 9784 22982 9812 24142
rect 9876 23866 9904 24278
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9036 22568 9088 22574
rect 8942 22536 8998 22545
rect 8852 22500 8904 22506
rect 9036 22510 9088 22516
rect 8942 22471 8998 22480
rect 8852 22442 8904 22448
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8864 22166 8892 22442
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 9048 21894 9076 22510
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8574 21584 8630 21593
rect 8574 21519 8630 21528
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7944 21146 7972 21286
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 8496 21010 8524 21422
rect 9048 21078 9076 21830
rect 9784 21690 9812 22918
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9876 21146 9904 23802
rect 10060 22778 10088 25094
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 23118 10732 24142
rect 10796 23866 10824 24618
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10796 23526 10824 23802
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10888 23254 10916 24686
rect 10876 23248 10928 23254
rect 10876 23190 10928 23196
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10060 22438 10088 22714
rect 10704 22642 10732 23054
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10888 22438 10916 23190
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9036 21072 9088 21078
rect 9968 21026 9996 22034
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 9036 21014 9088 21020
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 9784 20998 9996 21026
rect 8312 20398 8340 20946
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8312 19922 8340 20334
rect 8496 20262 8524 20946
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 9416 20210 9444 20538
rect 9508 20398 9536 20742
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9692 20330 9720 20878
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7944 19310 7972 19654
rect 8312 19514 8340 19858
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7668 18630 7696 19246
rect 7944 18698 7972 19246
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 8036 18902 8064 19178
rect 8496 18970 8524 20198
rect 9416 20182 9536 20210
rect 8666 19952 8722 19961
rect 8666 19887 8722 19896
rect 8760 19916 8812 19922
rect 8680 19854 8708 19887
rect 8760 19858 8812 19864
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 8772 18834 8800 19858
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9416 19514 9444 19654
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8772 18737 8800 18770
rect 9036 18760 9088 18766
rect 8482 18728 8538 18737
rect 7932 18692 7984 18698
rect 8482 18663 8538 18672
rect 8758 18728 8814 18737
rect 9036 18702 9088 18708
rect 8758 18663 8814 18672
rect 7932 18634 7984 18640
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18290 8340 18566
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7484 16998 7512 17682
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7668 16250 7696 17070
rect 7760 16794 7788 17546
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 8036 16658 8064 17138
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 8036 15706 8064 16594
rect 8220 16454 8248 17206
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 15706 8248 16390
rect 8312 16250 8340 16662
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8496 15706 8524 18663
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17338 8616 18022
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8588 17066 8616 17274
rect 8680 17134 8708 17478
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 15978 8616 17002
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 8220 15162 8248 15642
rect 8588 15570 8616 15914
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6932 14482 6960 14758
rect 7392 14550 7420 14894
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13734 6868 13806
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7300 13530 7328 13670
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7392 13190 7420 13874
rect 8036 13734 8064 14554
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 6932 12782 6960 13126
rect 8128 12986 8156 13330
rect 8206 13288 8262 13297
rect 8312 13258 8340 15506
rect 8680 14890 8708 17070
rect 8772 16998 8800 17682
rect 9048 17202 9076 18702
rect 9324 17814 9352 19178
rect 9416 18902 9444 19450
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9416 18630 9444 18838
rect 9508 18834 9536 20182
rect 9692 20058 9720 20266
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 17882 9444 18566
rect 9508 18358 9536 18770
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9312 17808 9364 17814
rect 9312 17750 9364 17756
rect 9508 17542 9536 18294
rect 9600 18290 9628 19382
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 18426 9720 18566
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 9048 16726 9076 17138
rect 9402 16824 9458 16833
rect 9402 16759 9458 16768
rect 9416 16726 9444 16759
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8772 16454 8800 16594
rect 9048 16522 9076 16662
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8772 15978 8800 16390
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8907 16108 8959 16114
rect 8959 16056 8984 16096
rect 8907 16050 8984 16056
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8956 15638 8984 16050
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 9048 15570 9076 16118
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8680 14618 8708 14826
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8206 13223 8262 13232
rect 8300 13252 8352 13258
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 6932 12102 6960 12718
rect 7760 12442 7788 12718
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7852 12306 7880 12650
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 12374 7972 12582
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 12300 7892 12306
rect 7760 12260 7840 12288
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11354 6960 12038
rect 7760 11354 7788 12260
rect 7840 12242 7892 12248
rect 7944 11898 7972 12310
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8220 11626 8248 13223
rect 8300 13194 8352 13200
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10674 6776 11154
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7668 10742 7696 11086
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 7668 10266 7696 10678
rect 7852 10674 7880 11222
rect 8220 11082 8248 11562
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7576 9518 7604 10066
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 8036 9382 8064 10066
rect 8312 9926 8340 13194
rect 8404 13190 8432 14418
rect 8680 14113 8708 14554
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8758 14240 8814 14249
rect 8758 14175 8814 14184
rect 8666 14104 8722 14113
rect 8666 14039 8722 14048
rect 8680 13814 8708 14039
rect 8496 13786 8708 13814
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8496 13002 8524 13786
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8404 12974 8524 13002
rect 8404 10062 8432 12974
rect 8588 12782 8616 13330
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12850 8708 13262
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8680 12442 8708 12786
rect 8772 12782 8800 14175
rect 8956 14006 8984 14282
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 9048 13258 9076 15506
rect 9232 15434 9260 15574
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 14618 9260 15370
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9232 14346 9260 14554
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9140 13802 9168 13942
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13530 9168 13738
rect 9232 13530 9260 13874
rect 9324 13814 9352 16526
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 15745 9444 16390
rect 9402 15736 9458 15745
rect 9402 15671 9458 15680
rect 9416 15638 9444 15671
rect 9404 15632 9456 15638
rect 9404 15574 9456 15580
rect 9416 15162 9444 15574
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14482 9444 14758
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9508 14249 9536 17478
rect 9600 14482 9628 17546
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9692 15638 9720 15914
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 9692 14618 9720 15574
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9494 14240 9550 14249
rect 9494 14175 9550 14184
rect 9692 13938 9720 14554
rect 9680 13932 9732 13938
rect 9600 13892 9680 13920
rect 9324 13786 9444 13814
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9416 13462 9444 13786
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9508 13394 9536 13670
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9600 13274 9628 13892
rect 9680 13874 9732 13880
rect 9784 13814 9812 20998
rect 10152 20466 10180 21830
rect 10428 21690 10456 22102
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21078 10732 21626
rect 10980 21622 11008 25486
rect 11808 25362 11836 27520
rect 12912 25362 12940 27520
rect 13924 25362 13952 27520
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 13912 25356 13964 25362
rect 13912 25298 13964 25304
rect 11808 24954 11836 25298
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11900 24410 11928 25094
rect 12912 24954 12940 25298
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 12900 24948 12952 24954
rect 12900 24890 12952 24896
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 12268 24342 12296 24686
rect 12440 24676 12492 24682
rect 12440 24618 12492 24624
rect 12256 24336 12308 24342
rect 12256 24278 12308 24284
rect 12268 23866 12296 24278
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11256 22234 11284 22374
rect 11244 22228 11296 22234
rect 11244 22170 11296 22176
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10888 21146 10916 21422
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10704 20602 10732 21014
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9876 19922 9904 20334
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10888 19990 10916 21082
rect 10980 20806 11008 21422
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20262 11008 20742
rect 11348 20466 11376 23666
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11532 23254 11560 23530
rect 12268 23474 12296 23802
rect 12176 23446 12296 23474
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 11532 22692 11560 23190
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11612 22704 11664 22710
rect 11532 22664 11612 22692
rect 11612 22646 11664 22652
rect 11900 22098 11928 23054
rect 12176 22234 12204 23446
rect 12452 23254 12480 24618
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 13188 23730 13216 24142
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 12728 23254 12756 23666
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12452 22778 12480 23190
rect 13740 23118 13768 25094
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 13004 22574 13032 22918
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12176 21418 12204 21966
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 12176 21010 12204 21354
rect 12268 21078 12296 22510
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12820 22166 12848 22374
rect 13740 22234 13768 23054
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 11808 20534 11836 20946
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11808 20262 11836 20470
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 19514 9904 19858
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 10888 19446 10916 19926
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9876 19174 9904 19314
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18766 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18290 9996 18566
rect 10152 18290 10180 18702
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18426 10824 18566
rect 10980 18426 11008 20198
rect 11808 19922 11836 20198
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11808 19446 11836 19858
rect 12176 19514 12204 19858
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9876 16436 9904 18158
rect 9968 17542 9996 18226
rect 10232 18216 10284 18222
rect 10152 18164 10232 18170
rect 10152 18158 10284 18164
rect 10152 18142 10272 18158
rect 10336 18154 10364 18294
rect 10796 18154 10824 18362
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10324 18148 10376 18154
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17678 10088 18022
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 10060 17066 10088 17614
rect 10152 17542 10180 18142
rect 10324 18090 10376 18096
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 9956 16448 10008 16454
rect 9876 16408 9956 16436
rect 9956 16390 10008 16396
rect 9968 15910 9996 16390
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 10060 15502 10088 17002
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 14822 10088 15438
rect 10152 15366 10180 17478
rect 10336 17338 10364 17682
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10612 17066 10640 17750
rect 10796 17746 10824 18090
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10980 17610 11008 18226
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10980 17338 11008 17546
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10796 16833 10824 17070
rect 10782 16824 10838 16833
rect 10782 16759 10838 16768
rect 10796 16726 10824 16759
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10520 16250 10548 16526
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10796 16046 10824 16458
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15570 10824 15982
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10152 15094 10180 15302
rect 10796 15094 10824 15506
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10152 14482 10180 15030
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9968 14006 9996 14418
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10060 13870 10088 14039
rect 10612 14006 10640 14214
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10048 13864 10100 13870
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9416 13246 9628 13274
rect 9692 13786 9812 13814
rect 9968 13812 10048 13814
rect 9968 13806 10100 13812
rect 9968 13786 10088 13806
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11762 8524 12106
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8496 11286 8524 11698
rect 8668 11620 8720 11626
rect 8772 11608 8800 12038
rect 8720 11580 8800 11608
rect 8668 11562 8720 11568
rect 8772 11354 8800 11580
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8772 10810 8800 11290
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8772 10606 8800 10746
rect 9416 10606 9444 13246
rect 9692 12424 9720 13786
rect 9968 13530 9996 13786
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9876 13376 9904 13466
rect 9956 13388 10008 13394
rect 9876 13348 9956 13376
rect 9956 13330 10008 13336
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9508 12396 9720 12424
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7116 8906 7144 9318
rect 7760 9110 7788 9318
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7760 8634 7788 9046
rect 8036 9042 8064 9318
rect 9416 9110 9444 10542
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 8036 8294 8064 8978
rect 9508 8945 9536 12396
rect 9772 12368 9824 12374
rect 9692 12328 9772 12356
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 11830 9628 12174
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9692 11558 9720 12328
rect 9772 12310 9824 12316
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11286 9720 11494
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9784 10810 9812 12038
rect 9876 11626 9904 12718
rect 9968 12646 9996 13330
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12170 9996 12582
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10060 11762 10088 12174
rect 10152 12102 10180 12650
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9876 11354 9904 11562
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9876 10810 9904 11290
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9494 8936 9550 8945
rect 9494 8871 9550 8880
rect 10060 8566 10088 11698
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 10810 10732 14758
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10796 12374 10824 14554
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 11898 10824 12310
rect 10888 11898 10916 14418
rect 10980 14006 11008 17274
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11256 17066 11284 17138
rect 11624 17134 11652 18634
rect 11808 18630 11836 18770
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11150 16824 11206 16833
rect 11256 16794 11284 17002
rect 11150 16759 11206 16768
rect 11244 16788 11296 16794
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10980 13530 11008 13942
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10980 12986 11008 13466
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10980 12442 11008 12922
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10980 11558 11008 12174
rect 11072 11694 11100 13194
rect 11164 12646 11192 16759
rect 11244 16730 11296 16736
rect 11624 16454 11652 17070
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11256 15366 11284 15982
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11256 12986 11284 15302
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10980 10606 11008 11494
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 1766 54 1992 82
rect 4160 128 4212 134
rect 4160 70 4212 76
rect 5262 128 5318 480
rect 5262 76 5264 128
rect 5316 76 5318 128
rect 1766 0 1822 54
rect 5262 0 5318 76
rect 8496 82 8524 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 8758 82 8814 480
rect 11072 134 11100 11630
rect 11164 2446 11192 12106
rect 11348 12102 11376 14894
rect 11440 14822 11468 14962
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14618 11468 14758
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11440 12850 11468 14282
rect 11532 13734 11560 14418
rect 11624 14346 11652 16390
rect 11716 15570 11744 16594
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 15366 11744 15506
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 14822 11744 15302
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11716 14414 11744 14758
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11532 12374 11560 13670
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11624 12238 11652 13738
rect 11716 13394 11744 14350
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 12986 11744 13330
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11808 12442 11836 18566
rect 12176 18426 12204 19450
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12544 18222 12572 18294
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12452 17882 12480 18090
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 11992 16522 12020 17682
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12084 17270 12112 17478
rect 12544 17338 12572 17682
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12544 16794 12572 17274
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 12452 15978 12480 16594
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11348 11830 11376 12038
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11348 11354 11376 11766
rect 11532 11694 11560 12038
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11900 6225 11928 14282
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 14074 12020 14214
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12084 12782 12112 15846
rect 12544 15570 12572 16730
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12360 13394 12388 14486
rect 12452 14482 12480 15098
rect 12544 14618 12572 15506
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12452 14074 12480 14418
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12360 12442 12388 13330
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12636 9674 12664 21966
rect 12820 21690 12848 22102
rect 12900 21956 12952 21962
rect 12900 21898 12952 21904
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12820 21418 12848 21626
rect 12912 21486 12940 21898
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12820 19514 12848 21354
rect 12912 21146 12940 21422
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 13452 21004 13504 21010
rect 13504 20964 13584 20992
rect 13452 20946 13504 20952
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 12912 20398 12940 20742
rect 13188 20466 13216 20742
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12820 18290 12848 18634
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12912 17814 12940 20334
rect 13556 20262 13584 20964
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13004 19378 13032 19654
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13004 18970 13032 19314
rect 13096 19310 13124 19790
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13360 19168 13412 19174
rect 13174 19136 13230 19145
rect 13360 19110 13412 19116
rect 13174 19071 13230 19080
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16726 12756 16934
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12728 16114 12756 16526
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15706 12756 16050
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12820 15638 12848 17070
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12820 14958 12848 15438
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12820 14618 12848 14894
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13462 12848 13806
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12544 9646 12664 9674
rect 12544 6798 12572 9646
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 11886 6216 11942 6225
rect 11886 6151 11942 6160
rect 12912 5710 12940 17546
rect 13188 17338 13216 19071
rect 13372 18902 13400 19110
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13004 14550 13032 15846
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13188 14482 13216 14826
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13280 13814 13308 18090
rect 13372 18086 13400 18838
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 16980 13400 18022
rect 13464 17882 13492 18362
rect 13556 18358 13584 20198
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13556 17746 13584 18294
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 16992 13504 16998
rect 13372 16952 13452 16980
rect 13452 16934 13504 16940
rect 13464 15978 13492 16934
rect 13556 16794 13584 17682
rect 13648 16794 13676 21830
rect 13832 19854 13860 25094
rect 13924 24954 13952 25298
rect 14844 24954 14872 27526
rect 14922 27520 14978 27526
rect 15580 27526 15990 27554
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14844 24750 14872 24890
rect 15488 24818 15516 25230
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14108 23866 14136 24210
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14384 23866 14412 24142
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 14108 23526 14136 23802
rect 14384 23594 14412 23802
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14372 23588 14424 23594
rect 14372 23530 14424 23536
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14108 22778 14136 23462
rect 14476 23322 14504 23666
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 14200 22778 14228 23190
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 14108 21622 14136 22034
rect 14200 21690 14228 22714
rect 14292 22642 14320 22986
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14188 19984 14240 19990
rect 14240 19944 14320 19972
rect 14188 19926 14240 19932
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 14292 19174 14320 19944
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18834 14320 19110
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13740 17882 13768 18702
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 18290 14412 18566
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14476 18154 14504 20878
rect 14568 20466 14596 24618
rect 14648 24064 14700 24070
rect 14648 24006 14700 24012
rect 14660 21570 14688 24006
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14924 23588 14976 23594
rect 14924 23530 14976 23536
rect 14936 23186 14964 23530
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14844 22506 14872 23054
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 14740 22500 14792 22506
rect 14740 22442 14792 22448
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14752 22234 14780 22442
rect 15488 22234 15516 22578
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 14752 22030 14780 22170
rect 15580 22098 15608 27526
rect 15934 27520 15990 27526
rect 17038 27520 17094 28000
rect 18050 27520 18106 28000
rect 19062 27554 19118 28000
rect 18800 27526 19118 27554
rect 16580 26172 16632 26178
rect 16580 26114 16632 26120
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15672 24954 15700 25434
rect 16592 25362 16620 26114
rect 17052 25498 17080 27520
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15752 24336 15804 24342
rect 15752 24278 15804 24284
rect 15764 23866 15792 24278
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15672 22778 15700 23122
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15580 21593 15608 21830
rect 15566 21584 15622 21593
rect 14660 21542 14780 21570
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14660 20806 14688 21422
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14568 20058 14596 20402
rect 14660 20330 14688 20538
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14660 19514 14688 20266
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14464 18148 14516 18154
rect 14464 18090 14516 18096
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13832 17610 13860 17818
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14660 16794 14688 17070
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13188 13786 13308 13814
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13096 12442 13124 12582
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13004 11830 13032 12242
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 13188 4622 13216 13786
rect 13464 13530 13492 14418
rect 13556 14113 13584 15914
rect 13648 15706 13676 16730
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13832 16182 13860 16662
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13542 14104 13598 14113
rect 13542 14039 13598 14048
rect 13648 13802 13676 14486
rect 13740 14346 13768 15438
rect 13832 15026 13860 15574
rect 14384 15502 14412 16526
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13280 11558 13308 12310
rect 13556 12170 13584 13262
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 5273 13308 11494
rect 13648 7993 13676 13738
rect 13832 13734 13860 14758
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14074 14412 14214
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13740 12986 13768 13398
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13832 12782 13860 13670
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12442 13860 12718
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13634 7984 13690 7993
rect 13634 7919 13690 7928
rect 13266 5264 13322 5273
rect 13266 5199 13322 5208
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 14476 2961 14504 16526
rect 14752 16130 14780 21542
rect 15566 21519 15622 21528
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14844 19718 14872 20402
rect 15304 19990 15332 21354
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15488 20602 15516 20946
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 18290 14872 19654
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 19926
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15396 17882 15424 18702
rect 15488 18426 15516 18838
rect 15672 18766 15700 19790
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15856 18358 15884 25094
rect 16592 24954 16620 25298
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 15948 24070 15976 24686
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 15948 23633 15976 24006
rect 16408 23730 16436 24006
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16500 23662 16528 24550
rect 16488 23656 16540 23662
rect 15934 23624 15990 23633
rect 16488 23598 16540 23604
rect 15934 23559 15990 23568
rect 16960 23322 16988 24550
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22692 16436 22918
rect 16488 22704 16540 22710
rect 16408 22664 16488 22692
rect 16408 22506 16436 22664
rect 16488 22646 16540 22652
rect 16684 22642 16712 23054
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16396 22500 16448 22506
rect 16396 22442 16448 22448
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15948 21486 15976 22102
rect 16500 21690 16528 22442
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16500 20602 16528 20742
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16026 19952 16082 19961
rect 16026 19887 16082 19896
rect 16040 19854 16068 19887
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19378 16068 19790
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17270 15332 17682
rect 15580 17610 15608 18022
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15764 17338 15792 18022
rect 15856 17882 15884 18294
rect 16408 17882 16436 19178
rect 16592 18873 16620 22374
rect 16684 22166 16712 22578
rect 16672 22160 16724 22166
rect 16672 22102 16724 22108
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 19378 16896 20266
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16856 19168 16908 19174
rect 16960 19145 16988 19246
rect 16856 19110 16908 19116
rect 16946 19136 17002 19145
rect 16578 18864 16634 18873
rect 16868 18834 16896 19110
rect 16946 19071 17002 19080
rect 16578 18799 16634 18808
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16868 18426 16896 18770
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16658 15516 17002
rect 16408 16998 16436 17818
rect 16592 17270 16620 18090
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17338 16804 17614
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16948 17128 17000 17134
rect 17052 17105 17080 24550
rect 17144 22098 17172 24618
rect 17868 24132 17920 24138
rect 17868 24074 17920 24080
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 17236 22778 17264 23122
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17144 21690 17172 22034
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17316 21072 17368 21078
rect 17512 21049 17540 21830
rect 17316 21014 17368 21020
rect 17498 21040 17554 21049
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 19718 17264 20878
rect 17328 20602 17356 21014
rect 17498 20975 17554 20984
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17328 20058 17356 20538
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17328 18737 17356 18770
rect 17314 18728 17370 18737
rect 17314 18663 17370 18672
rect 17328 18426 17356 18663
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17328 17134 17356 17478
rect 17316 17128 17368 17134
rect 16948 17070 17000 17076
rect 17038 17096 17094 17105
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16594
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14660 16102 14780 16130
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 15292 16108 15344 16114
rect 14660 15026 14688 16102
rect 15292 16050 15344 16056
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15706 14780 15982
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14660 14618 14688 14962
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14844 13462 14872 14962
rect 15304 14958 15332 16050
rect 16132 15638 16160 16118
rect 16408 15978 16436 16934
rect 16960 16590 16988 17070
rect 17316 17070 17368 17076
rect 17038 17031 17094 17040
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16684 16114 16712 16526
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16960 15638 16988 16526
rect 17052 16250 17080 16662
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17236 15638 17264 17002
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 16132 15094 16160 15574
rect 17604 15570 17632 18022
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 16408 14618 16436 15438
rect 17604 15162 17632 15506
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15396 13802 15424 14010
rect 15488 13938 15516 14350
rect 15764 14006 15792 14350
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15212 13462 15240 13738
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15396 13394 15424 13738
rect 16132 13734 16160 14486
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16960 14006 16988 14418
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16132 13462 16160 13670
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12986 15424 13330
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 17880 11665 17908 24074
rect 17972 23769 18000 24686
rect 18064 24342 18092 27520
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18248 25362 18276 26182
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18248 24954 18276 25298
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 18616 24886 18644 25094
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 18052 24336 18104 24342
rect 18052 24278 18104 24284
rect 17958 23760 18014 23769
rect 17958 23695 18014 23704
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18156 23322 18184 23598
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17972 19514 18000 19926
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 18064 13297 18092 22918
rect 18510 22672 18566 22681
rect 18510 22607 18566 22616
rect 18524 22574 18552 22607
rect 18512 22568 18564 22574
rect 18512 22510 18564 22516
rect 18708 22137 18736 24618
rect 18800 23866 18828 27526
rect 19062 27520 19118 27526
rect 20074 27520 20130 28000
rect 21178 27520 21234 28000
rect 22190 27520 22246 28000
rect 23202 27520 23258 28000
rect 24214 27520 24270 28000
rect 25318 27554 25374 28000
rect 25056 27526 25374 27554
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18984 24177 19012 24686
rect 19352 24682 19380 25298
rect 19522 24712 19578 24721
rect 19340 24676 19392 24682
rect 19522 24647 19578 24656
rect 19340 24618 19392 24624
rect 19536 24274 19564 24647
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19499 24268 19564 24274
rect 19551 24216 19564 24268
rect 19499 24210 19564 24216
rect 18970 24168 19026 24177
rect 18970 24103 19026 24112
rect 19076 23866 19104 24210
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 19260 23662 19288 24006
rect 19536 23730 19564 24210
rect 20088 23798 20116 27520
rect 21192 24410 21220 27520
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 22204 23866 22232 27520
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 19260 23322 19288 23598
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 19890 23216 19946 23225
rect 19890 23151 19892 23160
rect 19944 23151 19946 23160
rect 19892 23122 19944 23128
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 19062 23080 19118 23089
rect 18892 22778 18920 23054
rect 19062 23015 19118 23024
rect 19076 22778 19104 23015
rect 19904 22778 19932 23122
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19524 22568 19576 22574
rect 19522 22536 19524 22545
rect 19576 22536 19578 22545
rect 19522 22471 19578 22480
rect 19536 22438 19564 22471
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19996 22137 20024 23462
rect 18694 22128 18750 22137
rect 18420 22092 18472 22098
rect 19982 22128 20038 22137
rect 18694 22063 18750 22072
rect 19524 22092 19576 22098
rect 18420 22034 18472 22040
rect 19982 22063 20038 22072
rect 19524 22034 19576 22040
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18156 20466 18184 20742
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18248 20330 18276 20878
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18156 20210 18184 20266
rect 18340 20210 18368 21354
rect 18432 21332 18460 22034
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18524 21457 18552 21830
rect 18788 21480 18840 21486
rect 18510 21448 18566 21457
rect 18788 21422 18840 21428
rect 18510 21383 18566 21392
rect 18512 21344 18564 21350
rect 18432 21304 18512 21332
rect 18512 21286 18564 21292
rect 18524 20913 18552 21286
rect 18510 20904 18566 20913
rect 18800 20874 18828 21422
rect 19536 21350 19564 22034
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18510 20839 18566 20848
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18800 20330 18828 20810
rect 19076 20602 19104 20946
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18156 20182 18368 20210
rect 18340 19854 18368 20182
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 19352 19514 19380 19858
rect 19536 19825 19564 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19522 19816 19578 19825
rect 19522 19751 19578 19760
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18156 18290 18184 18566
rect 18708 18358 18736 19246
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19076 18834 19104 19178
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19076 18426 19104 18770
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18248 17338 18276 18090
rect 18328 17808 18380 17814
rect 18328 17750 18380 17756
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18248 16250 18276 17138
rect 18340 17134 18368 17750
rect 18708 17678 18736 18294
rect 19352 17882 19380 19450
rect 19536 19446 19564 19654
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20088 18193 20116 23530
rect 21744 22817 21772 23598
rect 21730 22808 21786 22817
rect 21730 22743 21786 22752
rect 21364 22092 21416 22098
rect 21364 22034 21416 22040
rect 21376 21554 21404 22034
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 20074 18184 20130 18193
rect 20074 18119 20130 18128
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18432 17338 18460 17614
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 19444 16998 19472 17682
rect 22112 17066 22140 23598
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 22480 21622 22508 22034
rect 23216 21962 23244 27520
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19444 16833 19472 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19430 16824 19486 16833
rect 19622 16816 19918 16836
rect 19430 16759 19486 16768
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18800 16250 18828 16594
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 23492 14385 23520 23530
rect 24228 22234 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 25056 23798 25084 27526
rect 25318 27520 25374 27526
rect 26330 27520 26386 28000
rect 27342 27520 27398 28000
rect 25044 23792 25096 23798
rect 25044 23734 25096 23740
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 26344 20058 26372 27520
rect 27356 23866 27384 27520
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 24216 19916 24268 19922
rect 24216 19858 24268 19864
rect 24228 19378 24256 19858
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 21454 14376 21510 14385
rect 21376 14346 21454 14362
rect 21364 14340 21454 14346
rect 21416 14334 21454 14340
rect 21454 14311 21510 14320
rect 23478 14376 23534 14385
rect 23478 14311 23534 14320
rect 21364 14282 21416 14288
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 18050 13288 18106 13297
rect 18050 13223 18106 13232
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 17960 11688 18012 11694
rect 17866 11656 17922 11665
rect 17960 11630 18012 11636
rect 17866 11591 17922 11600
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14462 2952 14518 2961
rect 14462 2887 14518 2896
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 8496 54 8814 82
rect 11060 128 11112 134
rect 11060 70 11112 76
rect 12254 128 12310 480
rect 12254 76 12256 128
rect 12308 76 12310 128
rect 8758 0 8814 54
rect 12254 0 12310 76
rect 15396 82 15424 10406
rect 15750 82 15806 480
rect 17972 134 18000 11630
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 25962 7984 26018 7993
rect 25962 7919 26018 7928
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 22466 5264 22522 5273
rect 22466 5199 22522 5208
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 15396 54 15806 82
rect 17960 128 18012 134
rect 17960 70 18012 76
rect 19246 128 19302 480
rect 19246 76 19248 128
rect 19300 76 19302 128
rect 15750 0 15806 54
rect 19246 0 19302 76
rect 22480 82 22508 5199
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 22742 82 22798 480
rect 22480 54 22798 82
rect 25976 82 26004 7919
rect 26238 82 26294 480
rect 25976 54 26294 82
rect 22742 0 22798 54
rect 26238 0 26294 54
<< via2 >>
rect 110 25336 166 25392
rect 3146 26832 3202 26888
rect 478 21936 534 21992
rect 1582 20576 1638 20632
rect 110 20032 166 20088
rect 110 10784 166 10840
rect 110 9696 166 9752
rect 2686 23840 2742 23896
rect 2962 23432 3018 23488
rect 2778 22480 2834 22536
rect 2870 20848 2926 20904
rect 2226 17448 2282 17504
rect 2134 16496 2190 16552
rect 1674 8880 1730 8936
rect 110 8744 166 8800
rect 110 7656 166 7712
rect 1858 12280 1914 12336
rect 110 6568 166 6624
rect 1582 6160 1638 6216
rect 110 5616 166 5672
rect 110 4528 166 4584
rect 110 3440 166 3496
rect 1398 2896 1454 2952
rect 1306 2760 1362 2816
rect 1214 1944 1270 2000
rect 3146 18128 3202 18184
rect 2502 13640 2558 13696
rect 4618 27512 4674 27568
rect 4158 23024 4214 23080
rect 4250 22616 4306 22672
rect 3514 22344 3570 22400
rect 3514 17040 3570 17096
rect 3882 21664 3938 21720
rect 4526 20984 4582 21040
rect 4802 19760 4858 19816
rect 4066 18808 4122 18864
rect 2870 11192 2926 11248
rect 3514 12008 3570 12064
rect 3882 15408 3938 15464
rect 4526 15700 4582 15736
rect 4526 15680 4528 15700
rect 4528 15680 4580 15700
rect 4580 15680 4582 15700
rect 4618 11600 4674 11656
rect 5538 25744 5594 25800
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5446 23704 5502 23760
rect 6458 24112 6514 24168
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5538 22072 5594 22128
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 7654 24656 7710 24712
rect 6642 22616 6698 22672
rect 6642 21392 6698 21448
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 7194 16768 7250 16824
rect 5170 14320 5226 14376
rect 2134 992 2190 1048
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9218 23568 9274 23624
rect 8758 23160 8814 23216
rect 8942 22480 8998 22536
rect 8574 21528 8630 21584
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 8666 19896 8722 19952
rect 8482 18672 8538 18728
rect 8758 18672 8814 18728
rect 8206 13232 8262 13288
rect 9402 16768 9458 16824
rect 8758 14184 8814 14240
rect 8666 14048 8722 14104
rect 9402 15680 9458 15736
rect 9494 14184 9550 14240
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10782 16768 10838 16824
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10046 14048 10102 14104
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 9494 8880 9550 8936
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11150 16768 11206 16824
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 13174 19080 13230 19136
rect 11886 6160 11942 6216
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 13542 14048 13598 14104
rect 13634 7928 13690 7984
rect 13266 5208 13322 5264
rect 15566 21528 15622 21584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15934 23568 15990 23624
rect 16026 19896 16082 19952
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 16578 18808 16634 18864
rect 16946 19080 17002 19136
rect 17498 20984 17554 21040
rect 17314 18672 17370 18728
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 17038 17040 17094 17096
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 17958 23704 18014 23760
rect 18510 22616 18566 22672
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19522 24656 19578 24712
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 18970 24112 19026 24168
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19890 23180 19946 23216
rect 19890 23160 19892 23180
rect 19892 23160 19944 23180
rect 19944 23160 19946 23180
rect 19062 23024 19118 23080
rect 19522 22516 19524 22536
rect 19524 22516 19576 22536
rect 19576 22516 19578 22536
rect 19522 22480 19578 22516
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 18694 22072 18750 22128
rect 19982 22072 20038 22128
rect 18510 21392 18566 21448
rect 18510 20848 18566 20904
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19522 19760 19578 19816
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 21730 22752 21786 22808
rect 20074 18128 20130 18184
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19430 16768 19486 16824
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 21454 14320 21510 14376
rect 23478 14320 23534 14376
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18050 13232 18106 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 17866 11600 17922 11656
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14462 2896 14518 2952
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 25962 7928 26018 7984
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 22466 5208 22522 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 4613 27570 4679 27573
rect 6678 27570 6684 27572
rect 4613 27568 6684 27570
rect 4613 27512 4618 27568
rect 4674 27512 6684 27568
rect 4613 27510 6684 27512
rect 4613 27507 4679 27510
rect 6678 27508 6684 27510
rect 6748 27508 6754 27572
rect 0 27344 480 27464
rect 62 26890 122 27344
rect 3141 26890 3207 26893
rect 62 26888 3207 26890
rect 62 26832 3146 26888
rect 3202 26832 3207 26888
rect 62 26830 3207 26832
rect 3141 26827 3207 26830
rect 0 26256 480 26376
rect 62 25802 122 26256
rect 5533 25802 5599 25805
rect 62 25800 5599 25802
rect 62 25744 5538 25800
rect 5594 25744 5599 25800
rect 62 25742 5599 25744
rect 5533 25739 5599 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25392 480 25424
rect 0 25336 110 25392
rect 166 25336 480 25392
rect 0 25304 480 25336
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 7649 24714 7715 24717
rect 19517 24714 19583 24717
rect 7649 24712 19583 24714
rect 7649 24656 7654 24712
rect 7710 24656 19522 24712
rect 19578 24656 19583 24712
rect 7649 24654 19583 24656
rect 7649 24651 7715 24654
rect 19517 24651 19583 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24216 480 24336
rect 62 23898 122 24216
rect 6453 24170 6519 24173
rect 18965 24170 19031 24173
rect 6453 24168 19031 24170
rect 6453 24112 6458 24168
rect 6514 24112 18970 24168
rect 19026 24112 19031 24168
rect 6453 24110 19031 24112
rect 6453 24107 6519 24110
rect 18965 24107 19031 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2681 23898 2747 23901
rect 62 23896 2747 23898
rect 62 23840 2686 23896
rect 2742 23840 2747 23896
rect 62 23838 2747 23840
rect 2681 23835 2747 23838
rect 5441 23762 5507 23765
rect 17953 23762 18019 23765
rect 5441 23760 18019 23762
rect 5441 23704 5446 23760
rect 5502 23704 17958 23760
rect 18014 23704 18019 23760
rect 5441 23702 18019 23704
rect 5441 23699 5507 23702
rect 17953 23699 18019 23702
rect 9213 23626 9279 23629
rect 15929 23626 15995 23629
rect 9213 23624 15995 23626
rect 9213 23568 9218 23624
rect 9274 23568 15934 23624
rect 15990 23568 15995 23624
rect 9213 23566 15995 23568
rect 9213 23563 9279 23566
rect 15929 23563 15995 23566
rect 2814 23428 2820 23492
rect 2884 23490 2890 23492
rect 2957 23490 3023 23493
rect 2884 23488 3023 23490
rect 2884 23432 2962 23488
rect 3018 23432 3023 23488
rect 2884 23430 3023 23432
rect 2884 23428 2890 23430
rect 2957 23427 3023 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 8753 23218 8819 23221
rect 19885 23218 19951 23221
rect 8753 23216 19951 23218
rect 8753 23160 8758 23216
rect 8814 23160 19890 23216
rect 19946 23160 19951 23216
rect 8753 23158 19951 23160
rect 8753 23155 8819 23158
rect 19885 23155 19951 23158
rect 62 22674 122 23128
rect 4153 23082 4219 23085
rect 19057 23082 19123 23085
rect 4153 23080 19123 23082
rect 4153 23024 4158 23080
rect 4214 23024 19062 23080
rect 19118 23024 19123 23080
rect 4153 23022 19123 23024
rect 4153 23019 4219 23022
rect 19057 23019 19123 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 17718 22748 17724 22812
rect 17788 22810 17794 22812
rect 21725 22810 21791 22813
rect 17788 22808 21791 22810
rect 17788 22752 21730 22808
rect 21786 22752 21791 22808
rect 17788 22750 21791 22752
rect 17788 22748 17794 22750
rect 21725 22747 21791 22750
rect 4245 22674 4311 22677
rect 62 22672 4311 22674
rect 62 22616 4250 22672
rect 4306 22616 4311 22672
rect 62 22614 4311 22616
rect 4245 22611 4311 22614
rect 6637 22674 6703 22677
rect 18505 22674 18571 22677
rect 6637 22672 18571 22674
rect 6637 22616 6642 22672
rect 6698 22616 18510 22672
rect 18566 22616 18571 22672
rect 6637 22614 18571 22616
rect 6637 22611 6703 22614
rect 18505 22611 18571 22614
rect 2773 22538 2839 22541
rect 8937 22538 9003 22541
rect 19517 22538 19583 22541
rect 2773 22536 9003 22538
rect 2773 22480 2778 22536
rect 2834 22480 8942 22536
rect 8998 22480 9003 22536
rect 2773 22478 9003 22480
rect 2773 22475 2839 22478
rect 8937 22475 9003 22478
rect 9078 22536 19583 22538
rect 9078 22480 19522 22536
rect 19578 22480 19583 22536
rect 9078 22478 19583 22480
rect 3509 22402 3575 22405
rect 9078 22402 9138 22478
rect 19517 22475 19583 22478
rect 3509 22400 9138 22402
rect 3509 22344 3514 22400
rect 3570 22344 9138 22400
rect 3509 22342 9138 22344
rect 3509 22339 3575 22342
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 62 21722 122 22176
rect 5533 22130 5599 22133
rect 6126 22130 6132 22132
rect 5533 22128 6132 22130
rect 5533 22072 5538 22128
rect 5594 22072 6132 22128
rect 5533 22070 6132 22072
rect 5533 22067 5599 22070
rect 6126 22068 6132 22070
rect 6196 22068 6202 22132
rect 18689 22130 18755 22133
rect 9630 22128 18755 22130
rect 9630 22072 18694 22128
rect 18750 22072 18755 22128
rect 9630 22070 18755 22072
rect 473 21994 539 21997
rect 9630 21994 9690 22070
rect 18689 22067 18755 22070
rect 18822 22068 18828 22132
rect 18892 22130 18898 22132
rect 19977 22130 20043 22133
rect 18892 22128 20043 22130
rect 18892 22072 19982 22128
rect 20038 22072 20043 22128
rect 18892 22070 20043 22072
rect 18892 22068 18898 22070
rect 19977 22067 20043 22070
rect 473 21992 9690 21994
rect 473 21936 478 21992
rect 534 21936 9690 21992
rect 473 21934 9690 21936
rect 473 21931 539 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 3877 21722 3943 21725
rect 62 21720 3943 21722
rect 62 21664 3882 21720
rect 3938 21664 3943 21720
rect 62 21662 3943 21664
rect 3877 21659 3943 21662
rect 8569 21586 8635 21589
rect 15561 21586 15627 21589
rect 8569 21584 15627 21586
rect 8569 21528 8574 21584
rect 8630 21528 15566 21584
rect 15622 21528 15627 21584
rect 8569 21526 15627 21528
rect 8569 21523 8635 21526
rect 15561 21523 15627 21526
rect 6637 21450 6703 21453
rect 18505 21450 18571 21453
rect 6637 21448 18571 21450
rect 6637 21392 6642 21448
rect 6698 21392 18510 21448
rect 18566 21392 18571 21448
rect 6637 21390 18571 21392
rect 6637 21387 6703 21390
rect 18505 21387 18571 21390
rect 10277 21248 10597 21249
rect 0 21088 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 62 20634 122 21088
rect 4521 21042 4587 21045
rect 17493 21042 17559 21045
rect 4521 21040 17559 21042
rect 4521 20984 4526 21040
rect 4582 20984 17498 21040
rect 17554 20984 17559 21040
rect 4521 20982 17559 20984
rect 4521 20979 4587 20982
rect 17493 20979 17559 20982
rect 2865 20906 2931 20909
rect 18505 20906 18571 20909
rect 2865 20904 18571 20906
rect 2865 20848 2870 20904
rect 2926 20848 18510 20904
rect 18566 20848 18571 20904
rect 2865 20846 18571 20848
rect 2865 20843 2931 20846
rect 18505 20843 18571 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 1577 20634 1643 20637
rect 62 20632 1643 20634
rect 62 20576 1582 20632
rect 1638 20576 1643 20632
rect 62 20574 1643 20576
rect 1577 20571 1643 20574
rect 10277 20160 10597 20161
rect 0 20088 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 20032 110 20088
rect 166 20032 480 20088
rect 0 20000 480 20032
rect 8661 19954 8727 19957
rect 16021 19954 16087 19957
rect 8661 19952 16087 19954
rect 8661 19896 8666 19952
rect 8722 19896 16026 19952
rect 16082 19896 16087 19952
rect 8661 19894 16087 19896
rect 8661 19891 8727 19894
rect 16021 19891 16087 19894
rect 4797 19818 4863 19821
rect 19517 19818 19583 19821
rect 4797 19816 19583 19818
rect 4797 19760 4802 19816
rect 4858 19760 19522 19816
rect 19578 19760 19583 19816
rect 4797 19758 19583 19760
rect 4797 19755 4863 19758
rect 19517 19755 19583 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19048 480 19168
rect 13169 19138 13235 19141
rect 16941 19138 17007 19141
rect 13169 19136 17007 19138
rect 13169 19080 13174 19136
rect 13230 19080 16946 19136
rect 17002 19080 17007 19136
rect 13169 19078 17007 19080
rect 13169 19075 13235 19078
rect 16941 19075 17007 19078
rect 10277 19072 10597 19073
rect 62 18730 122 19048
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 4061 18866 4127 18869
rect 16573 18866 16639 18869
rect 4061 18864 16639 18866
rect 4061 18808 4066 18864
rect 4122 18808 16578 18864
rect 16634 18808 16639 18864
rect 4061 18806 16639 18808
rect 4061 18803 4127 18806
rect 16573 18803 16639 18806
rect 8477 18730 8543 18733
rect 62 18728 8543 18730
rect 62 18672 8482 18728
rect 8538 18672 8543 18728
rect 62 18670 8543 18672
rect 8477 18667 8543 18670
rect 8753 18730 8819 18733
rect 17309 18730 17375 18733
rect 8753 18728 17375 18730
rect 8753 18672 8758 18728
rect 8814 18672 17314 18728
rect 17370 18672 17375 18728
rect 8753 18670 17375 18672
rect 8753 18667 8819 18670
rect 17309 18667 17375 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 3141 18186 3207 18189
rect 20069 18186 20135 18189
rect 3141 18184 20135 18186
rect 3141 18128 3146 18184
rect 3202 18128 20074 18184
rect 20130 18128 20135 18184
rect 3141 18126 20135 18128
rect 3141 18123 3207 18126
rect 20069 18123 20135 18126
rect 0 17960 480 18080
rect 10277 17984 10597 17985
rect 62 17506 122 17960
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 2221 17506 2287 17509
rect 62 17504 2287 17506
rect 62 17448 2226 17504
rect 2282 17448 2287 17504
rect 62 17446 2287 17448
rect 2221 17443 2287 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17008 480 17128
rect 3509 17098 3575 17101
rect 17033 17098 17099 17101
rect 3509 17096 17099 17098
rect 3509 17040 3514 17096
rect 3570 17040 17038 17096
rect 17094 17040 17099 17096
rect 3509 17038 17099 17040
rect 3509 17035 3575 17038
rect 17033 17035 17099 17038
rect 62 16554 122 17008
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 7189 16826 7255 16829
rect 9397 16826 9463 16829
rect 7189 16824 9463 16826
rect 7189 16768 7194 16824
rect 7250 16768 9402 16824
rect 9458 16768 9463 16824
rect 7189 16766 9463 16768
rect 7189 16763 7255 16766
rect 9397 16763 9463 16766
rect 10777 16826 10843 16829
rect 11145 16826 11211 16829
rect 19425 16826 19491 16829
rect 10777 16824 19491 16826
rect 10777 16768 10782 16824
rect 10838 16768 11150 16824
rect 11206 16768 19430 16824
rect 19486 16768 19491 16824
rect 10777 16766 19491 16768
rect 10777 16763 10843 16766
rect 11145 16763 11211 16766
rect 19425 16763 19491 16766
rect 2129 16554 2195 16557
rect 62 16552 2195 16554
rect 62 16496 2134 16552
rect 2190 16496 2195 16552
rect 62 16494 2195 16496
rect 2129 16491 2195 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 15920 480 16040
rect 62 15466 122 15920
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 4521 15738 4587 15741
rect 9397 15738 9463 15741
rect 4521 15736 9463 15738
rect 4521 15680 4526 15736
rect 4582 15680 9402 15736
rect 9458 15680 9463 15736
rect 4521 15678 9463 15680
rect 4521 15675 4587 15678
rect 9397 15675 9463 15678
rect 3877 15466 3943 15469
rect 62 15464 3943 15466
rect 62 15408 3882 15464
rect 3938 15408 3943 15464
rect 62 15406 3943 15408
rect 3877 15403 3943 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14832 480 14952
rect 62 14378 122 14832
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 5165 14378 5231 14381
rect 62 14376 5231 14378
rect 62 14320 5170 14376
rect 5226 14320 5231 14376
rect 62 14318 5231 14320
rect 5165 14315 5231 14318
rect 21449 14378 21515 14381
rect 23473 14378 23539 14381
rect 21449 14376 23539 14378
rect 21449 14320 21454 14376
rect 21510 14320 23478 14376
rect 23534 14320 23539 14376
rect 21449 14318 23539 14320
rect 21449 14315 21515 14318
rect 23473 14315 23539 14318
rect 8753 14242 8819 14245
rect 9489 14242 9555 14245
rect 8753 14240 9555 14242
rect 8753 14184 8758 14240
rect 8814 14184 9494 14240
rect 9550 14184 9555 14240
rect 8753 14182 9555 14184
rect 8753 14179 8819 14182
rect 9489 14179 9555 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8661 14106 8727 14109
rect 10041 14106 10107 14109
rect 13537 14106 13603 14109
rect 8661 14104 13603 14106
rect 8661 14048 8666 14104
rect 8722 14048 10046 14104
rect 10102 14048 13542 14104
rect 13598 14048 13603 14104
rect 8661 14046 13603 14048
rect 8661 14043 8727 14046
rect 10041 14043 10107 14046
rect 13537 14043 13603 14046
rect 0 13880 480 14000
rect 62 13698 122 13880
rect 2497 13698 2563 13701
rect 62 13696 2563 13698
rect 62 13640 2502 13696
rect 2558 13640 2563 13696
rect 62 13638 2563 13640
rect 2497 13635 2563 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8201 13290 8267 13293
rect 18045 13290 18111 13293
rect 8201 13288 18111 13290
rect 8201 13232 8206 13288
rect 8262 13232 18050 13288
rect 18106 13232 18111 13288
rect 8201 13230 18111 13232
rect 8201 13227 8267 13230
rect 18045 13227 18111 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12792 480 12912
rect 62 12338 122 12792
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1853 12338 1919 12341
rect 62 12336 1919 12338
rect 62 12280 1858 12336
rect 1914 12280 1919 12336
rect 62 12278 1919 12280
rect 1853 12275 1919 12278
rect 2814 12004 2820 12068
rect 2884 12066 2890 12068
rect 3509 12066 3575 12069
rect 2884 12064 3575 12066
rect 2884 12008 3514 12064
rect 3570 12008 3575 12064
rect 2884 12006 3575 12008
rect 2884 12004 2890 12006
rect 3509 12003 3575 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11704 480 11824
rect 62 11250 122 11704
rect 4613 11658 4679 11661
rect 17861 11658 17927 11661
rect 4613 11656 17927 11658
rect 4613 11600 4618 11656
rect 4674 11600 17866 11656
rect 17922 11600 17927 11656
rect 4613 11598 17927 11600
rect 4613 11595 4679 11598
rect 17861 11595 17927 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2865 11250 2931 11253
rect 62 11248 2931 11250
rect 62 11192 2870 11248
rect 2926 11192 2931 11248
rect 62 11190 2931 11192
rect 2865 11187 2931 11190
rect 5610 10912 5930 10913
rect 0 10840 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10784 110 10840
rect 166 10784 480 10840
rect 0 10752 480 10784
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5610 9824 5930 9825
rect 0 9752 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 0 9696 110 9752
rect 166 9696 480 9752
rect 0 9664 480 9696
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 1669 8938 1735 8941
rect 9489 8938 9555 8941
rect 1669 8936 9555 8938
rect 1669 8880 1674 8936
rect 1730 8880 9494 8936
rect 9550 8880 9555 8936
rect 1669 8878 9555 8880
rect 1669 8875 1735 8878
rect 9489 8875 9555 8878
rect 0 8800 480 8832
rect 0 8744 110 8800
rect 166 8744 480 8800
rect 0 8712 480 8744
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 13629 7986 13695 7989
rect 25957 7986 26023 7989
rect 13629 7984 26023 7986
rect 13629 7928 13634 7984
rect 13690 7928 25962 7984
rect 26018 7928 26023 7984
rect 13629 7926 26023 7928
rect 13629 7923 13695 7926
rect 25957 7923 26023 7926
rect 0 7712 480 7744
rect 0 7656 110 7712
rect 166 7656 480 7712
rect 0 7624 480 7656
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6624 480 6656
rect 0 6568 110 6624
rect 166 6568 480 6624
rect 0 6536 480 6568
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 1577 6218 1643 6221
rect 11881 6218 11947 6221
rect 1577 6216 11947 6218
rect 1577 6160 1582 6216
rect 1638 6160 11886 6216
rect 11942 6160 11947 6216
rect 1577 6158 11947 6160
rect 1577 6155 1643 6158
rect 11881 6155 11947 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5672 480 5704
rect 0 5616 110 5672
rect 166 5616 480 5672
rect 0 5584 480 5616
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 13261 5266 13327 5269
rect 22461 5266 22527 5269
rect 13261 5264 22527 5266
rect 13261 5208 13266 5264
rect 13322 5208 22466 5264
rect 22522 5208 22527 5264
rect 13261 5206 22527 5208
rect 13261 5203 13327 5206
rect 22461 5203 22527 5206
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4584 480 4616
rect 0 4528 110 4584
rect 166 4528 480 4584
rect 0 4496 480 4528
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3496 480 3528
rect 0 3440 110 3496
rect 166 3440 480 3496
rect 0 3408 480 3440
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 1393 2954 1459 2957
rect 14457 2954 14523 2957
rect 1393 2952 14523 2954
rect 1393 2896 1398 2952
rect 1454 2896 14462 2952
rect 14518 2896 14523 2952
rect 1393 2894 14523 2896
rect 1393 2891 1459 2894
rect 14457 2891 14523 2894
rect 1301 2818 1367 2821
rect 62 2816 1367 2818
rect 62 2760 1306 2816
rect 1362 2760 1367 2816
rect 62 2758 1367 2760
rect 62 2576 122 2758
rect 1301 2755 1367 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2456 480 2576
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 1209 2002 1275 2005
rect 62 2000 1275 2002
rect 62 1944 1214 2000
rect 1270 1944 1275 2000
rect 62 1942 1275 1944
rect 62 1488 122 1942
rect 1209 1939 1275 1942
rect 0 1368 480 1488
rect 2129 1050 2195 1053
rect 62 1048 2195 1050
rect 62 992 2134 1048
rect 2190 992 2195 1048
rect 62 990 2195 992
rect 62 536 122 990
rect 2129 987 2195 990
rect 0 416 480 536
<< via3 >>
rect 6684 27508 6748 27572
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 2820 23428 2884 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 17724 22748 17788 22812
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 6132 22068 6196 22132
rect 18828 22068 18892 22132
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 2820 12004 2884 12068
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 6683 27572 6749 27573
rect 6683 27508 6684 27572
rect 6748 27508 6749 27572
rect 6683 27507 6749 27508
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 2819 23492 2885 23493
rect 2819 23428 2820 23492
rect 2884 23428 2885 23492
rect 2819 23427 2885 23428
rect 2822 12069 2882 23427
rect 5610 22880 5931 23904
rect 6686 22898 6746 27507
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 2819 12068 2885 12069
rect 2819 12004 2820 12068
rect 2884 12004 2885 12068
rect 2819 12003 2885 12004
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 6598 22662 6834 22898
rect 6046 22132 6282 22218
rect 6046 22068 6132 22132
rect 6132 22068 6196 22132
rect 6196 22068 6282 22132
rect 6046 21982 6282 22068
rect 17638 22812 17874 22898
rect 17638 22748 17724 22812
rect 17724 22748 17788 22812
rect 17788 22748 17874 22812
rect 17638 22662 17874 22748
rect 18742 22132 18978 22218
rect 18742 22068 18828 22132
rect 18828 22068 18892 22132
rect 18892 22068 18978 22132
rect 18742 21982 18978 22068
<< metal5 >>
rect 6556 22898 17916 22940
rect 6556 22662 6598 22898
rect 6834 22662 17638 22898
rect 17874 22662 17916 22898
rect 6556 22620 17916 22662
rect 6004 22218 19020 22260
rect 6004 21982 6046 22218
rect 6282 21982 18742 22218
rect 18978 21982 19020 22218
rect 6004 21940 19020 21982
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_17
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_21 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_14 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_18
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_55
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_6
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_10
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_17
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_69
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 406 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 682 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_6
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_10
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_17
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_17
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _101_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 314 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _233_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_14
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 406 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _103_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_25
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_136
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 1472 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_13
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_17
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _213_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_35
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_39
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _166_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 406 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_13
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_14
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _150_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_19_146
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_175
timestamp 1586364061
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_148
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_17
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_25
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_130
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_164
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_168
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_25
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 314 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_142
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 130 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_52
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_75
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_160
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_37
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 406 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_8
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_18
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_22
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_26
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_42
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 314 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_85
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 406 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_151
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_164
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_177
timestamp 1586364061
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_201
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_216
timestamp 1586364061
transform 1 0 20976 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_228
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_55
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_77
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_116
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_132
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 590 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_162
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_177
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 866 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_194
timestamp 1586364061
transform 1 0 18952 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_52
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_169
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_177
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_216
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_228
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_66
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 314 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_180
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_197
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_209
timestamp 1586364061
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_13
timestamp 1586364061
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_30
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_52
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_nor3_4  _170_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 406 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_85
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_102
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_144
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_164
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_200
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_204
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_255
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_267
timestamp 1586364061
transform 1 0 25668 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_275
timestamp 1586364061
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_12
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_16
timestamp 1586364061
transform 1 0 2576 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_50
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_114
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_124
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_173
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_177
timestamp 1586364061
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_201
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 24380 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_257
timestamp 1586364061
transform 1 0 24748 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_269
timestamp 1586364061
transform 1 0 25852 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_8
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 866 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_20
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_24
timestamp 1586364061
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 406 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_36
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 1234 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 5520 0 -1 21216
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_42
timestamp 1586364061
transform 1 0 4968 0 -1 21216
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_61
timestamp 1586364061
transform 1 0 6716 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_65
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_99
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_103
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_122
timestamp 1586364061
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_140
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 590 592
use scs8hd_decap_3  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_168
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 590 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_183
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_187
timestamp 1586364061
transform 1 0 18308 0 -1 21216
box -38 -48 406 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_33_204
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_200
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 20608 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_215
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_212
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_227
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_239
timestamp 1586364061
transform 1 0 23092 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 3496 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_20
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 590 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_65
timestamp 1586364061
transform 1 0 7084 0 1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_90
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_97
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_102
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_139
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_191
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_198
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_202
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_206
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_222
timestamp 1586364061
transform 1 0 21528 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_234
timestamp 1586364061
transform 1 0 22632 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_242
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_51
timestamp 1586364061
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_55
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 590 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_61
timestamp 1586364061
transform 1 0 6716 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_97
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_130
timestamp 1586364061
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_8  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_189
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_200
timestamp 1586364061
transform 1 0 19504 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 21344 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_212
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_219
timestamp 1586364061
transform 1 0 21252 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 22448 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_236
timestamp 1586364061
transform 1 0 22816 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_248
timestamp 1586364061
transform 1 0 23920 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_260
timestamp 1586364061
transform 1 0 25024 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_272
timestamp 1586364061
transform 1 0 26128 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_17
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_21
timestamp 1586364061
transform 1 0 3036 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_38
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_90
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_94
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_107
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_115
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_139
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_174
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_178
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_187
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 20056 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_198
timestamp 1586364061
transform 1 0 19320 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_202
timestamp 1586364061
transform 1 0 19688 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_209
timestamp 1586364061
transform 1 0 20332 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_221
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_233
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_241
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 1932 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_22
timestamp 1586364061
transform 1 0 3128 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_36
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_59
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_69
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  FILLER_38_98
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_110
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_114
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_127
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_131
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_189
timestamp 1586364061
transform 1 0 18492 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_200
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_212
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_10
timestamp 1586364061
transform 1 0 2024 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_20
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_18
timestamp 1586364061
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_14
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_24
timestamp 1586364061
transform 1 0 3312 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_43
timestamp 1586364061
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_55
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_58
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_76
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_80
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_70
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_93
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_132
timestamp 1586364061
transform 1 0 13248 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_139
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_156
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_160
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_167
timestamp 1586364061
transform 1 0 16468 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_171
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 18308 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 18124 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_189
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_6  FILLER_40_191
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 590 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 19228 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_201
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_205
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_212
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_261
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_265
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 314 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_17
timestamp 1586364061
transform 1 0 2668 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_21
timestamp 1586364061
transform 1 0 3036 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 590 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_71
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_75
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_90
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 406 592
use scs8hd_decap_6  FILLER_41_96
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 590 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_102
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 130 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_164
timestamp 1586364061
transform 1 0 16192 0 1 24480
box -38 -48 406 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 16928 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_170
timestamp 1586364061
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_187
timestamp 1586364061
transform 1 0 18308 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_191
timestamp 1586364061
transform 1 0 18676 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_198
timestamp 1586364061
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_202
timestamp 1586364061
transform 1 0 19688 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_206
timestamp 1586364061
transform 1 0 20056 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_218
timestamp 1586364061
transform 1 0 21160 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_230
timestamp 1586364061
transform 1 0 22264 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_242
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_6
timestamp 1586364061
transform 1 0 1656 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_40
timestamp 1586364061
transform 1 0 4784 0 -1 25568
box -38 -48 406 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_53
timestamp 1586364061
transform 1 0 5980 0 -1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_61
timestamp 1586364061
transform 1 0 6716 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 7728 0 -1 25568
box -38 -48 866 592
use scs8hd_fill_1  FILLER_42_71
timestamp 1586364061
transform 1 0 7636 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_81
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_103
timestamp 1586364061
transform 1 0 10580 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_114
timestamp 1586364061
transform 1 0 11592 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_122
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_142
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_154
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_160
timestamp 1586364061
transform 1 0 15824 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_171
timestamp 1586364061
transform 1 0 16836 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_183
timestamp 1586364061
transform 1 0 17940 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_190
timestamp 1586364061
transform 1 0 18584 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_201
timestamp 1586364061
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_213
timestamp 1586364061
transform 1 0 20700 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5262 0 5318 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8758 0 8814 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 12254 0 12310 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15750 0 15806 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 19246 0 19302 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 22742 0 22798 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 7 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[2]
port 8 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[3]
port 9 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[4]
port 10 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[5]
port 11 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[6]
port 12 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[7]
port 13 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 14 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[0]
port 15 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[1]
port 16 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[2]
port 17 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[3]
port 18 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[4]
port 19 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[5]
port 20 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[6]
port 21 nsew default tristate
rlabel metal3 s 0 26256 480 26376 6 chanx_left_out[7]
port 22 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 chanx_left_out[8]
port 23 nsew default tristate
rlabel metal2 s 478 27520 534 28000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 1490 27520 1546 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 8758 27520 8814 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 21178 27520 21234 28000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 22190 27520 22246 28000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 26330 27520 26386 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 27342 27520 27398 28000 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 data_in
port 42 nsew default input
rlabel metal2 s 1766 0 1822 480 6 enable
port 43 nsew default input
rlabel metal3 s 0 15920 480 16040 6 left_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 0 17008 480 17128 6 left_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal3 s 0 17960 480 18080 6 left_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 0 10752 480 10872 6 left_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 0 11704 480 11824 6 left_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 0 12792 480 12912 6 left_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal3 s 0 13880 480 14000 6 left_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 0 14832 480 14952 6 left_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 0 9664 480 9784 6 left_top_grid_pin_10_
port 52 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 top_left_grid_pin_13_
port 53 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 top_right_grid_pin_11_
port 54 nsew default input
rlabel metal2 s 17038 27520 17094 28000 6 top_right_grid_pin_13_
port 55 nsew default input
rlabel metal2 s 18050 27520 18106 28000 6 top_right_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 top_right_grid_pin_1_
port 57 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 top_right_grid_pin_3_
port 58 nsew default input
rlabel metal2 s 12898 27520 12954 28000 6 top_right_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 top_right_grid_pin_7_
port 60 nsew default input
rlabel metal2 s 14922 27520 14978 28000 6 top_right_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
