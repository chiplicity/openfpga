magic
tech EFS8A
magscale 1 2
timestamp 1603801403
<< locali >>
rect 12909 16643 12943 16745
rect 9505 13923 9539 14025
<< viali >>
rect 12817 25449 12851 25483
rect 13921 25449 13955 25483
rect 8620 25313 8654 25347
rect 9816 25313 9850 25347
rect 11621 25313 11655 25347
rect 12633 25313 12667 25347
rect 13737 25313 13771 25347
rect 15828 25313 15862 25347
rect 8723 25109 8757 25143
rect 9919 25109 9953 25143
rect 11437 25109 11471 25143
rect 14289 25109 14323 25143
rect 15899 25109 15933 25143
rect 9229 24905 9263 24939
rect 9781 24905 9815 24939
rect 16313 24905 16347 24939
rect 7849 24769 7883 24803
rect 14565 24769 14599 24803
rect 15577 24769 15611 24803
rect 7364 24701 7398 24735
rect 8677 24701 8711 24735
rect 10425 24701 10459 24735
rect 10609 24701 10643 24735
rect 12541 24701 12575 24735
rect 13461 24701 13495 24735
rect 15761 24701 15795 24735
rect 11621 24633 11655 24667
rect 12449 24633 12483 24667
rect 14289 24633 14323 24667
rect 14381 24633 14415 24667
rect 7435 24565 7469 24599
rect 8493 24565 8527 24599
rect 8861 24565 8895 24599
rect 10977 24565 11011 24599
rect 12265 24565 12299 24599
rect 14013 24565 14047 24599
rect 15945 24565 15979 24599
rect 16865 24565 16899 24599
rect 14565 24361 14599 24395
rect 17049 24361 17083 24395
rect 11437 24293 11471 24327
rect 13001 24293 13035 24327
rect 4144 24225 4178 24259
rect 6596 24225 6630 24259
rect 8125 24225 8159 24259
rect 9781 24225 9815 24259
rect 15393 24225 15427 24259
rect 16865 24225 16899 24259
rect 18220 24225 18254 24259
rect 24568 24225 24602 24259
rect 11345 24157 11379 24191
rect 11989 24157 12023 24191
rect 12909 24157 12943 24191
rect 13185 24157 13219 24191
rect 15301 24157 15335 24191
rect 13829 24089 13863 24123
rect 18291 24089 18325 24123
rect 4215 24021 4249 24055
rect 6699 24021 6733 24055
rect 8033 24021 8067 24055
rect 8861 24021 8895 24055
rect 9965 24021 9999 24055
rect 12541 24021 12575 24055
rect 24639 24021 24673 24055
rect 3709 23817 3743 23851
rect 5273 23817 5307 23851
rect 6561 23817 6595 23851
rect 7665 23817 7699 23851
rect 9689 23817 9723 23851
rect 11345 23817 11379 23851
rect 15853 23817 15887 23851
rect 18521 23817 18555 23851
rect 18981 23817 19015 23851
rect 19809 23817 19843 23851
rect 21511 23817 21545 23851
rect 21925 23817 21959 23851
rect 25513 23817 25547 23851
rect 4169 23749 4203 23783
rect 20913 23749 20947 23783
rect 25145 23749 25179 23783
rect 8677 23681 8711 23715
rect 9137 23681 9171 23715
rect 10517 23681 10551 23715
rect 12909 23681 12943 23715
rect 14565 23681 14599 23715
rect 14841 23681 14875 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 3224 23613 3258 23647
rect 4772 23613 4806 23647
rect 7481 23613 7515 23647
rect 8125 23613 8159 23647
rect 11621 23613 11655 23647
rect 16129 23613 16163 23647
rect 18128 23613 18162 23647
rect 19324 23613 19358 23647
rect 20428 23613 20462 23647
rect 21440 23613 21474 23647
rect 24660 23613 24694 23647
rect 1547 23545 1581 23579
rect 4859 23545 4893 23579
rect 7389 23545 7423 23579
rect 8769 23545 8803 23579
rect 10241 23545 10275 23579
rect 10333 23545 10367 23579
rect 12541 23545 12575 23579
rect 12633 23545 12667 23579
rect 14657 23545 14691 23579
rect 16037 23545 16071 23579
rect 3295 23477 3329 23511
rect 8493 23477 8527 23511
rect 9965 23477 9999 23511
rect 12173 23477 12207 23511
rect 13461 23477 13495 23511
rect 14381 23477 14415 23511
rect 15485 23477 15519 23511
rect 17049 23477 17083 23511
rect 18199 23477 18233 23511
rect 19395 23477 19429 23511
rect 20499 23477 20533 23511
rect 24731 23477 24765 23511
rect 10793 23273 10827 23307
rect 12909 23273 12943 23307
rect 17325 23273 17359 23307
rect 7757 23205 7791 23239
rect 7849 23205 7883 23239
rect 8401 23205 8435 23239
rect 9781 23205 9815 23239
rect 9873 23205 9907 23239
rect 11437 23205 11471 23239
rect 13829 23205 13863 23239
rect 14381 23205 14415 23239
rect 15761 23205 15795 23239
rect 1476 23137 1510 23171
rect 2488 23137 2522 23171
rect 5641 23137 5675 23171
rect 6720 23137 6754 23171
rect 12541 23137 12575 23171
rect 17141 23137 17175 23171
rect 18296 23137 18330 23171
rect 11345 23069 11379 23103
rect 11621 23069 11655 23103
rect 13737 23069 13771 23103
rect 15669 23069 15703 23103
rect 16313 23069 16347 23103
rect 18383 23069 18417 23103
rect 10333 23001 10367 23035
rect 11161 23001 11195 23035
rect 1547 22933 1581 22967
rect 2559 22933 2593 22967
rect 6791 22933 6825 22967
rect 8677 22933 8711 22967
rect 3249 22729 3283 22763
rect 7113 22729 7147 22763
rect 8033 22729 8067 22763
rect 9781 22729 9815 22763
rect 11805 22729 11839 22763
rect 12265 22729 12299 22763
rect 13737 22729 13771 22763
rect 17233 22729 17267 22763
rect 9137 22661 9171 22695
rect 10057 22661 10091 22695
rect 3571 22593 3605 22627
rect 7481 22593 7515 22627
rect 8585 22593 8619 22627
rect 10609 22593 10643 22627
rect 10885 22593 10919 22627
rect 12541 22593 12575 22627
rect 13185 22593 13219 22627
rect 14381 22593 14415 22627
rect 14841 22593 14875 22627
rect 16221 22593 16255 22627
rect 16497 22593 16531 22627
rect 1444 22525 1478 22559
rect 2237 22525 2271 22559
rect 2488 22525 2522 22559
rect 3468 22525 3502 22559
rect 3893 22525 3927 22559
rect 1547 22457 1581 22491
rect 8677 22457 8711 22491
rect 10977 22457 11011 22491
rect 11529 22457 11563 22491
rect 12633 22457 12667 22491
rect 14473 22457 14507 22491
rect 16037 22457 16071 22491
rect 16313 22457 16347 22491
rect 1961 22389 1995 22423
rect 2559 22389 2593 22423
rect 2973 22389 3007 22423
rect 8309 22389 8343 22423
rect 14105 22389 14139 22423
rect 15577 22389 15611 22423
rect 18061 22389 18095 22423
rect 18521 22389 18555 22423
rect 7757 22185 7791 22219
rect 8309 22185 8343 22219
rect 11897 22185 11931 22219
rect 13645 22185 13679 22219
rect 14657 22185 14691 22219
rect 16221 22185 16255 22219
rect 11069 22117 11103 22151
rect 11621 22117 11655 22151
rect 13185 22117 13219 22151
rect 16497 22117 16531 22151
rect 17877 22117 17911 22151
rect 2028 22049 2062 22083
rect 3040 22049 3074 22083
rect 6009 22049 6043 22083
rect 7088 22049 7122 22083
rect 8585 22049 8619 22083
rect 9940 22049 9974 22083
rect 12449 22049 12483 22083
rect 13001 22049 13035 22083
rect 14232 22049 14266 22083
rect 14335 22049 14369 22083
rect 15336 22049 15370 22083
rect 15439 22049 15473 22083
rect 18245 22049 18279 22083
rect 10977 21981 11011 22015
rect 16405 21981 16439 22015
rect 16681 21981 16715 22015
rect 7159 21913 7193 21947
rect 10011 21913 10045 21947
rect 10425 21913 10459 21947
rect 2099 21845 2133 21879
rect 3111 21845 3145 21879
rect 6193 21845 6227 21879
rect 15761 21845 15795 21879
rect 6561 21641 6595 21675
rect 8953 21641 8987 21675
rect 9321 21641 9355 21675
rect 10701 21641 10735 21675
rect 12265 21641 12299 21675
rect 13461 21641 13495 21675
rect 14197 21641 14231 21675
rect 15117 21641 15151 21675
rect 15761 21641 15795 21675
rect 16129 21641 16163 21675
rect 18245 21641 18279 21675
rect 2559 21573 2593 21607
rect 5917 21573 5951 21607
rect 16865 21573 16899 21607
rect 6929 21505 6963 21539
rect 7481 21505 7515 21539
rect 16313 21505 16347 21539
rect 17233 21505 17267 21539
rect 1444 21437 1478 21471
rect 1869 21437 1903 21471
rect 2488 21437 2522 21471
rect 2881 21437 2915 21471
rect 3468 21437 3502 21471
rect 3893 21437 3927 21471
rect 4480 21437 4514 21471
rect 4905 21437 4939 21471
rect 5733 21437 5767 21471
rect 7849 21437 7883 21471
rect 8217 21437 8251 21471
rect 8401 21437 8435 21471
rect 9540 21437 9574 21471
rect 10333 21437 10367 21471
rect 10977 21437 11011 21471
rect 11345 21437 11379 21471
rect 12725 21437 12759 21471
rect 12909 21437 12943 21471
rect 14565 21437 14599 21471
rect 15301 21437 15335 21471
rect 1547 21369 1581 21403
rect 3571 21369 3605 21403
rect 11529 21369 11563 21403
rect 11897 21369 11931 21403
rect 16405 21369 16439 21403
rect 2329 21301 2363 21335
rect 3249 21301 3283 21335
rect 4583 21301 4617 21335
rect 6193 21301 6227 21335
rect 8033 21301 8067 21335
rect 9643 21301 9677 21335
rect 12725 21301 12759 21335
rect 8769 21097 8803 21131
rect 10885 21097 10919 21131
rect 11943 21097 11977 21131
rect 13737 21097 13771 21131
rect 14013 21097 14047 21131
rect 15117 21097 15151 21131
rect 16221 21097 16255 21131
rect 16589 21097 16623 21131
rect 17601 21097 17635 21131
rect 6469 21029 6503 21063
rect 8170 21029 8204 21063
rect 10327 21029 10361 21063
rect 11529 21029 11563 21063
rect 13179 21029 13213 21063
rect 15622 21029 15656 21063
rect 1444 20961 1478 20995
rect 4721 20961 4755 20995
rect 11872 20961 11906 20995
rect 12817 20961 12851 20995
rect 17417 20961 17451 20995
rect 2421 20893 2455 20927
rect 6377 20893 6411 20927
rect 7849 20893 7883 20927
rect 9965 20893 9999 20927
rect 15301 20893 15335 20927
rect 6929 20825 6963 20859
rect 1547 20757 1581 20791
rect 4813 20757 4847 20791
rect 7389 20757 7423 20791
rect 7757 20757 7791 20791
rect 11253 20757 11287 20791
rect 12541 20757 12575 20791
rect 2237 20553 2271 20587
rect 4629 20553 4663 20587
rect 8953 20553 8987 20587
rect 10701 20553 10735 20587
rect 11897 20553 11931 20587
rect 14933 20553 14967 20587
rect 17417 20553 17451 20587
rect 18199 20553 18233 20587
rect 14657 20485 14691 20519
rect 16129 20485 16163 20519
rect 1961 20417 1995 20451
rect 7573 20417 7607 20451
rect 8033 20417 8067 20451
rect 13737 20417 13771 20451
rect 15577 20417 15611 20451
rect 16865 20417 16899 20451
rect 1460 20349 1494 20383
rect 2456 20349 2490 20383
rect 2881 20349 2915 20383
rect 5089 20349 5123 20383
rect 5825 20349 5859 20383
rect 9781 20349 9815 20383
rect 10977 20349 11011 20383
rect 18128 20349 18162 20383
rect 18521 20349 18555 20383
rect 1547 20281 1581 20315
rect 5917 20281 5951 20315
rect 7941 20281 7975 20315
rect 8395 20281 8429 20315
rect 9321 20281 9355 20315
rect 9689 20281 9723 20315
rect 10143 20281 10177 20315
rect 14099 20281 14133 20315
rect 15669 20281 15703 20315
rect 16497 20281 16531 20315
rect 2559 20213 2593 20247
rect 3433 20213 3467 20247
rect 6377 20213 6411 20247
rect 6837 20213 6871 20247
rect 12725 20213 12759 20247
rect 13277 20213 13311 20247
rect 13645 20213 13679 20247
rect 15301 20213 15335 20247
rect 2789 20009 2823 20043
rect 4445 20009 4479 20043
rect 6377 20009 6411 20043
rect 8125 20009 8159 20043
rect 8769 20009 8803 20043
rect 9965 20009 9999 20043
rect 10701 20009 10735 20043
rect 11345 20009 11379 20043
rect 12817 20009 12851 20043
rect 13921 20009 13955 20043
rect 1777 19941 1811 19975
rect 1869 19941 1903 19975
rect 4721 19941 4755 19975
rect 4813 19941 4847 19975
rect 5365 19941 5399 19975
rect 6929 19941 6963 19975
rect 7481 19941 7515 19975
rect 13363 19941 13397 19975
rect 15761 19941 15795 19975
rect 17325 19941 17359 19975
rect 18705 19941 18739 19975
rect 8309 19873 8343 19907
rect 9965 19873 9999 19907
rect 10149 19873 10183 19907
rect 11529 19873 11563 19907
rect 11805 19873 11839 19907
rect 18797 19873 18831 19907
rect 6837 19805 6871 19839
rect 9505 19805 9539 19839
rect 13001 19805 13035 19839
rect 15669 19805 15703 19839
rect 16129 19805 16163 19839
rect 17233 19805 17267 19839
rect 17877 19805 17911 19839
rect 2329 19737 2363 19771
rect 14381 19737 14415 19771
rect 5733 19669 5767 19703
rect 8493 19669 8527 19703
rect 11161 19669 11195 19703
rect 12449 19669 12483 19703
rect 16589 19669 16623 19703
rect 4353 19465 4387 19499
rect 6285 19465 6319 19499
rect 9781 19465 9815 19499
rect 11897 19465 11931 19499
rect 12173 19465 12207 19499
rect 15669 19465 15703 19499
rect 17417 19465 17451 19499
rect 19073 19465 19107 19499
rect 15945 19397 15979 19431
rect 2329 19329 2363 19363
rect 14473 19329 14507 19363
rect 15117 19329 15151 19363
rect 2697 19261 2731 19295
rect 3065 19261 3099 19295
rect 3801 19261 3835 19295
rect 4813 19261 4847 19295
rect 6837 19261 6871 19295
rect 7757 19261 7791 19295
rect 8677 19261 8711 19295
rect 9045 19261 9079 19295
rect 10609 19261 10643 19295
rect 11529 19261 11563 19295
rect 12449 19261 12483 19295
rect 12909 19261 12943 19295
rect 13185 19261 13219 19295
rect 13829 19261 13863 19295
rect 18061 19261 18095 19295
rect 18153 19261 18187 19295
rect 1685 19193 1719 19227
rect 1777 19193 1811 19227
rect 3157 19193 3191 19227
rect 5175 19193 5209 19227
rect 6561 19193 6595 19227
rect 7199 19193 7233 19227
rect 10517 19193 10551 19227
rect 10971 19193 11005 19227
rect 14289 19193 14323 19227
rect 14565 19193 14599 19227
rect 16497 19193 16531 19227
rect 16589 19193 16623 19227
rect 17141 19193 17175 19227
rect 17877 19193 17911 19227
rect 4721 19125 4755 19159
rect 5733 19125 5767 19159
rect 8401 19125 8435 19159
rect 8677 19125 8711 19159
rect 10149 19125 10183 19159
rect 13553 19125 13587 19159
rect 1685 18921 1719 18955
rect 2973 18921 3007 18955
rect 6745 18921 6779 18955
rect 7205 18921 7239 18955
rect 7573 18921 7607 18955
rect 8585 18921 8619 18955
rect 9781 18921 9815 18955
rect 12265 18921 12299 18955
rect 13185 18921 13219 18955
rect 15761 18921 15795 18955
rect 16957 18921 16991 18955
rect 2145 18853 2179 18887
rect 4629 18853 4663 18887
rect 11707 18853 11741 18887
rect 16037 18853 16071 18887
rect 16589 18853 16623 18887
rect 17233 18853 17267 18887
rect 17601 18853 17635 18887
rect 18153 18853 18187 18887
rect 6009 18785 6043 18819
rect 7757 18785 7791 18819
rect 8033 18785 8067 18819
rect 9965 18785 9999 18819
rect 10241 18785 10275 18819
rect 11345 18785 11379 18819
rect 13093 18785 13127 18819
rect 13553 18785 13587 18819
rect 2053 18717 2087 18751
rect 3341 18717 3375 18751
rect 4537 18717 4571 18751
rect 15945 18717 15979 18751
rect 17509 18717 17543 18751
rect 18981 18717 19015 18751
rect 2605 18649 2639 18683
rect 5089 18649 5123 18683
rect 9413 18649 9447 18683
rect 5549 18581 5583 18615
rect 6193 18581 6227 18615
rect 9137 18581 9171 18615
rect 10793 18581 10827 18615
rect 11253 18581 11287 18615
rect 14105 18581 14139 18615
rect 4537 18377 4571 18411
rect 7389 18377 7423 18411
rect 9505 18377 9539 18411
rect 13093 18377 13127 18411
rect 14841 18377 14875 18411
rect 17877 18377 17911 18411
rect 2421 18309 2455 18343
rect 9210 18309 9244 18343
rect 10747 18309 10781 18343
rect 10885 18309 10919 18343
rect 15209 18309 15243 18343
rect 16313 18309 16347 18343
rect 1869 18241 1903 18275
rect 3433 18241 3467 18275
rect 3801 18241 3835 18275
rect 6653 18241 6687 18275
rect 9413 18241 9447 18275
rect 10977 18241 11011 18275
rect 11345 18241 11379 18275
rect 15761 18241 15795 18275
rect 16773 18241 16807 18275
rect 18061 18241 18095 18275
rect 5549 18173 5583 18207
rect 7757 18173 7791 18207
rect 8033 18173 8067 18207
rect 9275 18173 9309 18207
rect 12265 18173 12299 18207
rect 12449 18173 12483 18207
rect 13921 18173 13955 18207
rect 18153 18173 18187 18207
rect 1685 18105 1719 18139
rect 1961 18105 1995 18139
rect 3249 18105 3283 18139
rect 3525 18105 3559 18139
rect 4905 18105 4939 18139
rect 8585 18105 8619 18139
rect 9045 18105 9079 18139
rect 10609 18105 10643 18139
rect 11713 18105 11747 18139
rect 14242 18105 14276 18139
rect 15577 18105 15611 18139
rect 15853 18105 15887 18139
rect 2789 18037 2823 18071
rect 6101 18037 6135 18071
rect 7573 18037 7607 18071
rect 8861 18037 8895 18071
rect 10057 18037 10091 18071
rect 10425 18037 10459 18071
rect 12633 18037 12667 18071
rect 13737 18037 13771 18071
rect 17509 18037 17543 18071
rect 2789 17833 2823 17867
rect 3433 17833 3467 17867
rect 4537 17833 4571 17867
rect 7481 17833 7515 17867
rect 8493 17833 8527 17867
rect 9505 17833 9539 17867
rect 10333 17833 10367 17867
rect 10701 17833 10735 17867
rect 11345 17833 11379 17867
rect 12173 17833 12207 17867
rect 13185 17833 13219 17867
rect 14381 17833 14415 17867
rect 16221 17833 16255 17867
rect 17509 17833 17543 17867
rect 18153 17833 18187 17867
rect 1777 17765 1811 17799
rect 1869 17765 1903 17799
rect 2421 17765 2455 17799
rect 5226 17765 5260 17799
rect 7935 17765 7969 17799
rect 13823 17765 13857 17799
rect 15663 17765 15697 17799
rect 9689 17697 9723 17731
rect 11897 17697 11931 17731
rect 12449 17697 12483 17731
rect 17325 17697 17359 17731
rect 18680 17697 18714 17731
rect 4905 17629 4939 17663
rect 7573 17629 7607 17663
rect 10057 17629 10091 17663
rect 13461 17629 13495 17663
rect 14657 17629 14691 17663
rect 15301 17629 15335 17663
rect 9965 17561 9999 17595
rect 5825 17493 5859 17527
rect 7113 17493 7147 17527
rect 9137 17493 9171 17527
rect 9854 17493 9888 17527
rect 11805 17493 11839 17527
rect 18751 17493 18785 17527
rect 1777 17289 1811 17323
rect 3709 17289 3743 17323
rect 6653 17289 6687 17323
rect 8493 17289 8527 17323
rect 8861 17289 8895 17323
rect 10701 17289 10735 17323
rect 11069 17289 11103 17323
rect 12081 17289 12115 17323
rect 13645 17289 13679 17323
rect 16681 17289 16715 17323
rect 17141 17289 17175 17323
rect 18245 17289 18279 17323
rect 2973 17221 3007 17255
rect 5917 17221 5951 17255
rect 18705 17221 18739 17255
rect 1961 17153 1995 17187
rect 2605 17153 2639 17187
rect 6193 17153 6227 17187
rect 7573 17153 7607 17187
rect 9873 17153 9907 17187
rect 13277 17153 13311 17187
rect 3341 17085 3375 17119
rect 4077 17085 4111 17119
rect 4537 17085 4571 17119
rect 4997 17085 5031 17119
rect 9321 17085 9355 17119
rect 9781 17085 9815 17119
rect 10885 17085 10919 17119
rect 11345 17085 11379 17119
rect 12817 17085 12851 17119
rect 13093 17085 13127 17119
rect 14105 17085 14139 17119
rect 14657 17085 14691 17119
rect 14841 17085 14875 17119
rect 15761 17085 15795 17119
rect 17877 17085 17911 17119
rect 18061 17085 18095 17119
rect 2053 17017 2087 17051
rect 5359 17017 5393 17051
rect 7113 17017 7147 17051
rect 7481 17017 7515 17051
rect 7935 17017 7969 17051
rect 9229 17017 9263 17051
rect 15301 17017 15335 17051
rect 16082 17017 16116 17051
rect 4905 16949 4939 16983
rect 10333 16949 10367 16983
rect 11805 16949 11839 16983
rect 13921 16949 13955 16983
rect 15669 16949 15703 16983
rect 1685 16745 1719 16779
rect 2513 16745 2547 16779
rect 4261 16745 4295 16779
rect 5273 16745 5307 16779
rect 9321 16745 9355 16779
rect 9873 16745 9907 16779
rect 12541 16745 12575 16779
rect 12909 16745 12943 16779
rect 13553 16745 13587 16779
rect 14657 16745 14691 16779
rect 15853 16745 15887 16779
rect 3433 16677 3467 16711
rect 4721 16677 4755 16711
rect 11069 16677 11103 16711
rect 11805 16677 11839 16711
rect 13829 16677 13863 16711
rect 15485 16677 15519 16711
rect 16405 16677 16439 16711
rect 17969 16677 18003 16711
rect 2237 16609 2271 16643
rect 3065 16609 3099 16643
rect 4077 16609 4111 16643
rect 4997 16609 5031 16643
rect 5365 16609 5399 16643
rect 6009 16609 6043 16643
rect 6193 16609 6227 16643
rect 7757 16609 7791 16643
rect 7849 16609 7883 16643
rect 9689 16609 9723 16643
rect 12633 16609 12667 16643
rect 12909 16609 12943 16643
rect 13185 16609 13219 16643
rect 19349 16609 19383 16643
rect 11437 16541 11471 16575
rect 13737 16541 13771 16575
rect 14381 16541 14415 16575
rect 16313 16541 16347 16575
rect 16957 16541 16991 16575
rect 17877 16541 17911 16575
rect 8217 16473 8251 16507
rect 8585 16473 8619 16507
rect 18429 16473 18463 16507
rect 8861 16405 8895 16439
rect 10517 16405 10551 16439
rect 10793 16405 10827 16439
rect 11234 16405 11268 16439
rect 11345 16405 11379 16439
rect 12081 16405 12115 16439
rect 12817 16405 12851 16439
rect 19533 16405 19567 16439
rect 2513 16201 2547 16235
rect 4353 16201 4387 16235
rect 9321 16201 9355 16235
rect 9873 16201 9907 16235
rect 11069 16201 11103 16235
rect 17877 16201 17911 16235
rect 18613 16201 18647 16235
rect 19349 16201 19383 16235
rect 3801 16133 3835 16167
rect 5549 16133 5583 16167
rect 9137 16133 9171 16167
rect 10701 16133 10735 16167
rect 17049 16133 17083 16167
rect 1593 16065 1627 16099
rect 3249 16065 3283 16099
rect 6653 16065 6687 16099
rect 8769 16065 8803 16099
rect 9229 16065 9263 16099
rect 10793 16065 10827 16099
rect 13277 16065 13311 16099
rect 15945 16065 15979 16099
rect 16497 16065 16531 16099
rect 18061 16065 18095 16099
rect 4721 15997 4755 16031
rect 5089 15997 5123 16031
rect 5641 15997 5675 16031
rect 5825 15997 5859 16031
rect 7573 15997 7607 16031
rect 7849 15997 7883 16031
rect 8401 15997 8435 16031
rect 9008 15997 9042 16031
rect 10572 15997 10606 16031
rect 12817 15997 12851 16031
rect 13093 15997 13127 16031
rect 14105 15997 14139 16031
rect 1685 15929 1719 15963
rect 2237 15929 2271 15963
rect 3065 15929 3099 15963
rect 3341 15929 3375 15963
rect 8861 15929 8895 15963
rect 10425 15929 10459 15963
rect 11529 15929 11563 15963
rect 14013 15929 14047 15963
rect 14467 15929 14501 15963
rect 16313 15929 16347 15963
rect 16589 15929 16623 15963
rect 6285 15861 6319 15895
rect 7205 15861 7239 15895
rect 7573 15861 7607 15895
rect 10241 15861 10275 15895
rect 11805 15861 11839 15895
rect 12173 15861 12207 15895
rect 13645 15861 13679 15895
rect 15025 15861 15059 15895
rect 15577 15861 15611 15895
rect 3249 15657 3283 15691
rect 3893 15657 3927 15691
rect 4261 15657 4295 15691
rect 5273 15657 5307 15691
rect 5549 15657 5583 15691
rect 7481 15657 7515 15691
rect 10609 15657 10643 15691
rect 14473 15657 14507 15691
rect 2329 15589 2363 15623
rect 2421 15589 2455 15623
rect 11529 15589 11563 15623
rect 12265 15589 12299 15623
rect 15663 15589 15697 15623
rect 17049 15589 17083 15623
rect 4077 15521 4111 15555
rect 5733 15521 5767 15555
rect 6285 15521 6319 15555
rect 7665 15521 7699 15555
rect 7849 15521 7883 15555
rect 8217 15521 8251 15555
rect 9965 15521 9999 15555
rect 11676 15521 11710 15555
rect 13093 15521 13127 15555
rect 13553 15521 13587 15555
rect 16221 15521 16255 15555
rect 17509 15521 17543 15555
rect 2973 15453 3007 15487
rect 6377 15453 6411 15487
rect 10333 15453 10367 15487
rect 11897 15453 11931 15487
rect 13737 15453 13771 15487
rect 15301 15453 15335 15487
rect 16589 15453 16623 15487
rect 8953 15385 8987 15419
rect 10241 15385 10275 15419
rect 1685 15317 1719 15351
rect 1961 15317 1995 15351
rect 4905 15317 4939 15351
rect 7021 15317 7055 15351
rect 9413 15317 9447 15351
rect 10103 15317 10137 15351
rect 11069 15317 11103 15351
rect 11805 15317 11839 15351
rect 12633 15317 12667 15351
rect 12909 15317 12943 15351
rect 14105 15317 14139 15351
rect 1777 15113 1811 15147
rect 4905 15113 4939 15147
rect 6193 15113 6227 15147
rect 6653 15113 6687 15147
rect 8033 15113 8067 15147
rect 8309 15113 8343 15147
rect 12081 15113 12115 15147
rect 13921 15113 13955 15147
rect 15393 15113 15427 15147
rect 17509 15113 17543 15147
rect 2973 15045 3007 15079
rect 16589 15045 16623 15079
rect 3433 14977 3467 15011
rect 4537 14977 4571 15011
rect 4997 14977 5031 15011
rect 13645 14977 13679 15011
rect 2145 14909 2179 14943
rect 2605 14909 2639 14943
rect 5917 14909 5951 14943
rect 7021 14909 7055 14943
rect 9137 14909 9171 14943
rect 10517 14909 10551 14943
rect 10977 14909 11011 14943
rect 12909 14909 12943 14943
rect 13461 14909 13495 14943
rect 14289 14909 14323 14943
rect 14657 14909 14691 14943
rect 15761 14909 15795 14943
rect 16681 14909 16715 14943
rect 17141 14909 17175 14943
rect 3157 14841 3191 14875
rect 3249 14841 3283 14875
rect 5318 14841 5352 14875
rect 9781 14841 9815 14875
rect 10609 14841 10643 14875
rect 4077 14773 4111 14807
rect 7205 14773 7239 14807
rect 8861 14773 8895 14807
rect 10057 14773 10091 14807
rect 11713 14773 11747 14807
rect 12725 14773 12759 14807
rect 16221 14773 16255 14807
rect 16865 14773 16899 14807
rect 3249 14569 3283 14603
rect 3893 14569 3927 14603
rect 5181 14569 5215 14603
rect 6653 14569 6687 14603
rect 7757 14569 7791 14603
rect 10793 14569 10827 14603
rect 12725 14569 12759 14603
rect 13461 14569 13495 14603
rect 14013 14569 14047 14603
rect 16129 14569 16163 14603
rect 16865 14569 16899 14603
rect 6095 14501 6129 14535
rect 9505 14501 9539 14535
rect 9689 14501 9723 14535
rect 12817 14501 12851 14535
rect 15853 14501 15887 14535
rect 2513 14433 2547 14467
rect 2973 14433 3007 14467
rect 4169 14433 4203 14467
rect 5733 14433 5767 14467
rect 7665 14433 7699 14467
rect 8217 14433 8251 14467
rect 9919 14433 9953 14467
rect 11529 14433 11563 14467
rect 11989 14433 12023 14467
rect 12964 14433 12998 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 16681 14433 16715 14467
rect 1685 14365 1719 14399
rect 1869 14365 1903 14399
rect 7205 14365 7239 14399
rect 7573 14365 7607 14399
rect 10057 14365 10091 14399
rect 13185 14365 13219 14399
rect 9137 14297 9171 14331
rect 11345 14297 11379 14331
rect 13093 14297 13127 14331
rect 4353 14229 4387 14263
rect 5549 14229 5583 14263
rect 8769 14229 8803 14263
rect 9836 14229 9870 14263
rect 10149 14229 10183 14263
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 2605 14025 2639 14059
rect 4169 14025 4203 14059
rect 5733 14025 5767 14059
rect 8125 14025 8159 14059
rect 9137 14025 9171 14059
rect 9505 14025 9539 14059
rect 11345 14025 11379 14059
rect 14289 14025 14323 14059
rect 15761 14025 15795 14059
rect 16681 14025 16715 14059
rect 4721 13957 4755 13991
rect 6009 13957 6043 13991
rect 8953 13957 8987 13991
rect 10149 13957 10183 13991
rect 12265 13957 12299 13991
rect 13553 13957 13587 13991
rect 14178 13957 14212 13991
rect 2237 13889 2271 13923
rect 3157 13889 3191 13923
rect 3433 13889 3467 13923
rect 8585 13889 8619 13923
rect 9045 13889 9079 13923
rect 9505 13889 9539 13923
rect 14381 13889 14415 13923
rect 14473 13889 14507 13923
rect 15393 13889 15427 13923
rect 16037 13889 16071 13923
rect 2973 13821 3007 13855
rect 4813 13821 4847 13855
rect 6469 13821 6503 13855
rect 7389 13821 7423 13855
rect 7665 13821 7699 13855
rect 8824 13821 8858 13855
rect 10241 13821 10275 13855
rect 10701 13821 10735 13855
rect 13093 13821 13127 13855
rect 15577 13821 15611 13855
rect 1593 13753 1627 13787
rect 1685 13753 1719 13787
rect 3249 13753 3283 13787
rect 5134 13753 5168 13787
rect 8677 13753 8711 13787
rect 11805 13753 11839 13787
rect 13185 13753 13219 13787
rect 14013 13753 14047 13787
rect 7205 13685 7239 13719
rect 9689 13685 9723 13719
rect 10333 13685 10367 13719
rect 13829 13685 13863 13719
rect 1409 13481 1443 13515
rect 5733 13481 5767 13515
rect 6101 13481 6135 13515
rect 7205 13481 7239 13515
rect 9137 13481 9171 13515
rect 11345 13481 11379 13515
rect 12173 13481 12207 13515
rect 12817 13481 12851 13515
rect 13185 13481 13219 13515
rect 14105 13481 14139 13515
rect 2605 13413 2639 13447
rect 5134 13413 5168 13447
rect 7481 13413 7515 13447
rect 15577 13413 15611 13447
rect 9505 13345 9539 13379
rect 9965 13345 9999 13379
rect 10112 13345 10146 13379
rect 11529 13345 11563 13379
rect 13093 13345 13127 13379
rect 13645 13345 13679 13379
rect 2513 13277 2547 13311
rect 4813 13277 4847 13311
rect 7389 13277 7423 13311
rect 7665 13277 7699 13311
rect 10333 13277 10367 13311
rect 11897 13277 11931 13311
rect 3065 13209 3099 13243
rect 10425 13209 10459 13243
rect 1961 13141 1995 13175
rect 8401 13141 8435 13175
rect 8677 13141 8711 13175
rect 10241 13141 10275 13175
rect 10977 13141 11011 13175
rect 11667 13141 11701 13175
rect 11805 13141 11839 13175
rect 3341 12937 3375 12971
rect 4905 12937 4939 12971
rect 5549 12937 5583 12971
rect 7021 12937 7055 12971
rect 8125 12937 8159 12971
rect 8769 12937 8803 12971
rect 9689 12937 9723 12971
rect 11897 12937 11931 12971
rect 12587 12937 12621 12971
rect 13093 12937 13127 12971
rect 14841 12937 14875 12971
rect 1777 12869 1811 12903
rect 2881 12869 2915 12903
rect 10057 12869 10091 12903
rect 12725 12869 12759 12903
rect 13829 12869 13863 12903
rect 14197 12869 14231 12903
rect 4169 12801 4203 12835
rect 6653 12801 6687 12835
rect 7205 12801 7239 12835
rect 8401 12801 8435 12835
rect 12817 12801 12851 12835
rect 5365 12733 5399 12767
rect 5917 12733 5951 12767
rect 10609 12733 10643 12767
rect 10885 12733 10919 12767
rect 11621 12733 11655 12767
rect 14013 12733 14047 12767
rect 14473 12733 14507 12767
rect 2329 12665 2363 12699
rect 2421 12665 2455 12699
rect 3893 12665 3927 12699
rect 3985 12665 4019 12699
rect 7526 12665 7560 12699
rect 8953 12665 8987 12699
rect 12449 12665 12483 12699
rect 13461 12665 13495 12699
rect 2145 12597 2179 12631
rect 3709 12597 3743 12631
rect 5273 12597 5307 12631
rect 10701 12597 10735 12631
rect 4629 12393 4663 12427
rect 4813 12393 4847 12427
rect 6837 12393 6871 12427
rect 7297 12393 7331 12427
rect 9413 12393 9447 12427
rect 9965 12393 9999 12427
rect 11621 12393 11655 12427
rect 11989 12393 12023 12427
rect 12449 12393 12483 12427
rect 13553 12393 13587 12427
rect 13921 12393 13955 12427
rect 1409 12325 1443 12359
rect 7986 12325 8020 12359
rect 10787 12325 10821 12359
rect 13185 12325 13219 12359
rect 2513 12257 2547 12291
rect 2973 12257 3007 12291
rect 3893 12257 3927 12291
rect 4721 12257 4755 12291
rect 5273 12257 5307 12291
rect 6653 12257 6687 12291
rect 12173 12257 12207 12291
rect 12725 12257 12759 12291
rect 3157 12189 3191 12223
rect 7665 12189 7699 12223
rect 10425 12189 10459 12223
rect 1869 12053 1903 12087
rect 2237 12053 2271 12087
rect 6561 12053 6595 12087
rect 8585 12053 8619 12087
rect 8861 12053 8895 12087
rect 11345 12053 11379 12087
rect 2881 11849 2915 11883
rect 5917 11849 5951 11883
rect 7941 11849 7975 11883
rect 9781 11849 9815 11883
rect 11897 11849 11931 11883
rect 12173 11849 12207 11883
rect 12909 11849 12943 11883
rect 13277 11849 13311 11883
rect 12633 11781 12667 11815
rect 3065 11713 3099 11747
rect 3341 11713 3375 11747
rect 4629 11713 4663 11747
rect 7573 11713 7607 11747
rect 8493 11713 8527 11747
rect 10609 11645 10643 11679
rect 12449 11645 12483 11679
rect 1501 11577 1535 11611
rect 1593 11577 1627 11611
rect 2145 11577 2179 11611
rect 3157 11577 3191 11611
rect 4537 11577 4571 11611
rect 4950 11577 4984 11611
rect 6929 11577 6963 11611
rect 7021 11577 7055 11611
rect 8585 11577 8619 11611
rect 9137 11577 9171 11611
rect 10149 11577 10183 11611
rect 10517 11577 10551 11611
rect 10971 11577 11005 11611
rect 2513 11509 2547 11543
rect 4169 11509 4203 11543
rect 5549 11509 5583 11543
rect 6285 11509 6319 11543
rect 6653 11509 6687 11543
rect 8309 11509 8343 11543
rect 11529 11509 11563 11543
rect 3341 11305 3375 11339
rect 6469 11305 6503 11339
rect 6929 11305 6963 11339
rect 7389 11305 7423 11339
rect 8953 11305 8987 11339
rect 11253 11305 11287 11339
rect 2145 11237 2179 11271
rect 4899 11237 4933 11271
rect 7665 11237 7699 11271
rect 8217 11237 8251 11271
rect 10425 11237 10459 11271
rect 11989 11237 12023 11271
rect 4537 11169 4571 11203
rect 6285 11169 6319 11203
rect 2053 11101 2087 11135
rect 2697 11101 2731 11135
rect 7573 11101 7607 11135
rect 10333 11101 10367 11135
rect 11897 11101 11931 11135
rect 1593 11033 1627 11067
rect 2973 11033 3007 11067
rect 5457 11033 5491 11067
rect 6193 11033 6227 11067
rect 10885 11033 10919 11067
rect 12449 11033 12483 11067
rect 8493 10965 8527 10999
rect 10149 10965 10183 10999
rect 12817 10965 12851 10999
rect 3341 10761 3375 10795
rect 3617 10761 3651 10795
rect 4537 10761 4571 10795
rect 6009 10761 6043 10795
rect 8658 10761 8692 10795
rect 2513 10693 2547 10727
rect 8401 10693 8435 10727
rect 8769 10693 8803 10727
rect 2881 10625 2915 10659
rect 4169 10625 4203 10659
rect 5733 10625 5767 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 12173 10625 12207 10659
rect 3433 10557 3467 10591
rect 4905 10557 4939 10591
rect 5181 10557 5215 10591
rect 6929 10557 6963 10591
rect 7297 10557 7331 10591
rect 8493 10557 8527 10591
rect 10793 10557 10827 10591
rect 11161 10557 11195 10591
rect 12817 10557 12851 10591
rect 1961 10489 1995 10523
rect 2053 10489 2087 10523
rect 10149 10489 10183 10523
rect 10241 10489 10275 10523
rect 12449 10489 12483 10523
rect 1777 10421 1811 10455
rect 4721 10421 4755 10455
rect 6561 10421 6595 10455
rect 6929 10421 6963 10455
rect 7941 10421 7975 10455
rect 9965 10421 9999 10455
rect 11897 10421 11931 10455
rect 2053 10217 2087 10251
rect 4445 10217 4479 10251
rect 4629 10217 4663 10251
rect 7573 10217 7607 10251
rect 8769 10217 8803 10251
rect 9321 10217 9355 10251
rect 9965 10217 9999 10251
rect 10517 10217 10551 10251
rect 7849 10149 7883 10183
rect 11161 10149 11195 10183
rect 11713 10149 11747 10183
rect 12541 10149 12575 10183
rect 2881 10081 2915 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 6101 10081 6135 10115
rect 6561 10081 6595 10115
rect 12633 10081 12667 10115
rect 1409 10013 1443 10047
rect 2421 10013 2455 10047
rect 6837 10013 6871 10047
rect 7205 10013 7239 10047
rect 7757 10013 7791 10047
rect 8401 10013 8435 10047
rect 11069 10013 11103 10047
rect 3525 9877 3559 9911
rect 4353 9673 4387 9707
rect 5641 9673 5675 9707
rect 6101 9673 6135 9707
rect 6561 9673 6595 9707
rect 8677 9673 8711 9707
rect 9367 9673 9401 9707
rect 9505 9673 9539 9707
rect 11805 9673 11839 9707
rect 12633 9673 12667 9707
rect 1593 9605 1627 9639
rect 2421 9605 2455 9639
rect 3985 9605 4019 9639
rect 9137 9605 9171 9639
rect 9689 9605 9723 9639
rect 11253 9605 11287 9639
rect 2973 9537 3007 9571
rect 3341 9537 3375 9571
rect 4445 9537 4479 9571
rect 7297 9537 7331 9571
rect 9597 9537 9631 9571
rect 1409 9469 1443 9503
rect 5365 9469 5399 9503
rect 10701 9469 10735 9503
rect 10885 9469 10919 9503
rect 2789 9401 2823 9435
rect 3065 9401 3099 9435
rect 4807 9401 4841 9435
rect 7618 9401 7652 9435
rect 9229 9401 9263 9435
rect 2053 9333 2087 9367
rect 7113 9333 7147 9367
rect 8217 9333 8251 9367
rect 4353 9129 4387 9163
rect 6285 9129 6319 9163
rect 8033 9129 8067 9163
rect 11069 9129 11103 9163
rect 2421 9061 2455 9095
rect 2973 9061 3007 9095
rect 4807 9061 4841 9095
rect 6790 9061 6824 9095
rect 7757 9061 7791 9095
rect 1685 8993 1719 9027
rect 4445 8993 4479 9027
rect 9781 8993 9815 9027
rect 11320 8993 11354 9027
rect 2329 8925 2363 8959
rect 6469 8925 6503 8959
rect 8217 8925 8251 8959
rect 9689 8925 9723 8959
rect 3709 8857 3743 8891
rect 3249 8789 3283 8823
rect 5365 8789 5399 8823
rect 7389 8789 7423 8823
rect 9229 8789 9263 8823
rect 11391 8789 11425 8823
rect 1593 8585 1627 8619
rect 2145 8585 2179 8619
rect 3709 8585 3743 8619
rect 5181 8585 5215 8619
rect 5871 8585 5905 8619
rect 8125 8585 8159 8619
rect 9781 8585 9815 8619
rect 11345 8585 11379 8619
rect 3249 8517 3283 8551
rect 6469 8517 6503 8551
rect 2697 8449 2731 8483
rect 4077 8449 4111 8483
rect 4537 8449 4571 8483
rect 7113 8449 7147 8483
rect 7481 8449 7515 8483
rect 8677 8449 8711 8483
rect 8953 8449 8987 8483
rect 1409 8381 1443 8415
rect 5641 8381 5675 8415
rect 5768 8381 5802 8415
rect 2513 8313 2547 8347
rect 2789 8313 2823 8347
rect 4261 8313 4295 8347
rect 4353 8313 4387 8347
rect 7205 8313 7239 8347
rect 8493 8313 8527 8347
rect 8769 8313 8803 8347
rect 1409 8041 1443 8075
rect 2237 8041 2271 8075
rect 2881 8041 2915 8075
rect 4353 8041 4387 8075
rect 6561 8041 6595 8075
rect 7665 8041 7699 8075
rect 8355 8041 8389 8075
rect 6837 7973 6871 8007
rect 3065 7905 3099 7939
rect 4353 7905 4387 7939
rect 7389 7905 7423 7939
rect 8284 7905 8318 7939
rect 6745 7837 6779 7871
rect 3249 7497 3283 7531
rect 3617 7497 3651 7531
rect 3893 7497 3927 7531
rect 4353 7497 4387 7531
rect 8309 7497 8343 7531
rect 4951 7429 4985 7463
rect 2145 7361 2179 7395
rect 6653 7361 6687 7395
rect 6837 7361 6871 7395
rect 2053 7293 2087 7327
rect 2697 7293 2731 7327
rect 3709 7293 3743 7327
rect 4848 7293 4882 7327
rect 5273 7293 5307 7327
rect 7389 7293 7423 7327
rect 6193 7157 6227 7191
rect 6929 6953 6963 6987
rect 1409 6817 1443 6851
rect 2053 6817 2087 6851
rect 3040 6817 3074 6851
rect 3111 6681 3145 6715
rect 7757 6613 7791 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 2651 6409 2685 6443
rect 3341 6409 3375 6443
rect 8125 6273 8159 6307
rect 1409 6205 1443 6239
rect 2548 6205 2582 6239
rect 2973 6205 3007 6239
rect 7757 6205 7791 6239
rect 8401 6205 8435 6239
rect 2421 6137 2455 6171
rect 7665 6137 7699 6171
rect 1547 5865 1581 5899
rect 2559 5865 2593 5899
rect 1476 5729 1510 5763
rect 2488 5729 2522 5763
rect 7665 5729 7699 5763
rect 8033 5525 8067 5559
rect 2237 5321 2271 5355
rect 2605 5321 2639 5355
rect 8033 5321 8067 5355
rect 1547 5185 1581 5219
rect 8677 5185 8711 5219
rect 1444 5117 1478 5151
rect 1869 5117 1903 5151
rect 8125 5117 8159 5151
rect 8309 5117 8343 5151
rect 7573 4981 7607 5015
rect 8953 4981 8987 5015
rect 1547 4777 1581 4811
rect 1444 4641 1478 4675
rect 1593 4233 1627 4267
rect 1547 3689 1581 3723
rect 1444 3553 1478 3587
rect 1547 3145 1581 3179
rect 2237 3077 2271 3111
rect 1476 2941 1510 2975
rect 1869 2941 1903 2975
rect 1547 2601 1581 2635
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 2488 2465 2522 2499
rect 2881 2465 2915 2499
rect 2559 2329 2593 2363
<< metal1 >>
rect 4062 26256 4068 26308
rect 4120 26296 4126 26308
rect 6546 26296 6552 26308
rect 4120 26268 6552 26296
rect 4120 26256 4126 26268
rect 6546 26256 6552 26268
rect 6604 26256 6610 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 12894 25480 12900 25492
rect 12851 25452 12900 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 12894 25440 12900 25452
rect 12952 25440 12958 25492
rect 13906 25480 13912 25492
rect 13867 25452 13912 25480
rect 13906 25440 13912 25452
rect 13964 25440 13970 25492
rect 4062 25304 4068 25356
rect 4120 25344 4126 25356
rect 8608 25347 8666 25353
rect 8608 25344 8620 25347
rect 4120 25316 8620 25344
rect 4120 25304 4126 25316
rect 8608 25313 8620 25316
rect 8654 25344 8666 25347
rect 9214 25344 9220 25356
rect 8654 25316 9220 25344
rect 8654 25313 8666 25316
rect 8608 25307 8666 25313
rect 9214 25304 9220 25316
rect 9272 25304 9278 25356
rect 9766 25304 9772 25356
rect 9824 25353 9830 25356
rect 9824 25347 9862 25353
rect 9850 25313 9862 25347
rect 11606 25344 11612 25356
rect 11567 25316 11612 25344
rect 9824 25307 9862 25313
rect 9824 25304 9830 25307
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 12618 25344 12624 25356
rect 12579 25316 12624 25344
rect 12618 25304 12624 25316
rect 12676 25304 12682 25356
rect 13725 25347 13783 25353
rect 13725 25313 13737 25347
rect 13771 25344 13783 25347
rect 13814 25344 13820 25356
rect 13771 25316 13820 25344
rect 13771 25313 13783 25316
rect 13725 25307 13783 25313
rect 13814 25304 13820 25316
rect 13872 25304 13878 25356
rect 15816 25347 15874 25353
rect 15816 25313 15828 25347
rect 15862 25344 15874 25347
rect 16298 25344 16304 25356
rect 15862 25316 16304 25344
rect 15862 25313 15874 25316
rect 15816 25307 15874 25313
rect 16298 25304 16304 25316
rect 16356 25304 16362 25356
rect 8711 25143 8769 25149
rect 8711 25109 8723 25143
rect 8757 25140 8769 25143
rect 9674 25140 9680 25152
rect 8757 25112 9680 25140
rect 8757 25109 8769 25112
rect 8711 25103 8769 25109
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 9907 25143 9965 25149
rect 9907 25109 9919 25143
rect 9953 25140 9965 25143
rect 10686 25140 10692 25152
rect 9953 25112 10692 25140
rect 9953 25109 9965 25112
rect 9907 25103 9965 25109
rect 10686 25100 10692 25112
rect 10744 25100 10750 25152
rect 11422 25140 11428 25152
rect 11383 25112 11428 25140
rect 11422 25100 11428 25112
rect 11480 25100 11486 25152
rect 14274 25140 14280 25152
rect 14235 25112 14280 25140
rect 14274 25100 14280 25112
rect 14332 25100 14338 25152
rect 15746 25100 15752 25152
rect 15804 25140 15810 25152
rect 15887 25143 15945 25149
rect 15887 25140 15899 25143
rect 15804 25112 15899 25140
rect 15804 25100 15810 25112
rect 15887 25109 15899 25112
rect 15933 25109 15945 25143
rect 15887 25103 15945 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 9214 24936 9220 24948
rect 9175 24908 9220 24936
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 9766 24936 9772 24948
rect 9727 24908 9772 24936
rect 9766 24896 9772 24908
rect 9824 24896 9830 24948
rect 16298 24936 16304 24948
rect 16259 24908 16304 24936
rect 16298 24896 16304 24908
rect 16356 24896 16362 24948
rect 7837 24803 7895 24809
rect 7837 24769 7849 24803
rect 7883 24800 7895 24803
rect 8754 24800 8760 24812
rect 7883 24772 8760 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 7352 24735 7410 24741
rect 7352 24701 7364 24735
rect 7398 24732 7410 24735
rect 7852 24732 7880 24763
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 14366 24760 14372 24812
rect 14424 24800 14430 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 14424 24772 14565 24800
rect 14424 24760 14430 24772
rect 14553 24769 14565 24772
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 14734 24760 14740 24812
rect 14792 24800 14798 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 14792 24772 15577 24800
rect 14792 24760 14798 24772
rect 15565 24769 15577 24772
rect 15611 24800 15623 24803
rect 15611 24772 15792 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 8665 24735 8723 24741
rect 8665 24732 8677 24735
rect 7398 24704 7880 24732
rect 8496 24704 8677 24732
rect 7398 24701 7410 24704
rect 7352 24695 7410 24701
rect 7006 24556 7012 24608
rect 7064 24596 7070 24608
rect 7423 24599 7481 24605
rect 7423 24596 7435 24599
rect 7064 24568 7435 24596
rect 7064 24556 7070 24568
rect 7423 24565 7435 24568
rect 7469 24565 7481 24599
rect 7423 24559 7481 24565
rect 8294 24556 8300 24608
rect 8352 24596 8358 24608
rect 8496 24605 8524 24704
rect 8665 24701 8677 24704
rect 8711 24701 8723 24735
rect 8665 24695 8723 24701
rect 9858 24692 9864 24744
rect 9916 24732 9922 24744
rect 10413 24735 10471 24741
rect 10413 24732 10425 24735
rect 9916 24704 10425 24732
rect 9916 24692 9922 24704
rect 10413 24701 10425 24704
rect 10459 24732 10471 24735
rect 10597 24735 10655 24741
rect 10597 24732 10609 24735
rect 10459 24704 10609 24732
rect 10459 24701 10471 24704
rect 10413 24695 10471 24701
rect 10597 24701 10609 24704
rect 10643 24701 10655 24735
rect 10597 24695 10655 24701
rect 12529 24735 12587 24741
rect 12529 24701 12541 24735
rect 12575 24701 12587 24735
rect 12529 24695 12587 24701
rect 11606 24664 11612 24676
rect 11519 24636 11612 24664
rect 11606 24624 11612 24636
rect 11664 24664 11670 24676
rect 12158 24664 12164 24676
rect 11664 24636 12164 24664
rect 11664 24624 11670 24636
rect 12158 24624 12164 24636
rect 12216 24624 12222 24676
rect 12434 24664 12440 24676
rect 12395 24636 12440 24664
rect 12434 24624 12440 24636
rect 12492 24624 12498 24676
rect 8481 24599 8539 24605
rect 8481 24596 8493 24599
rect 8352 24568 8493 24596
rect 8352 24556 8358 24568
rect 8481 24565 8493 24568
rect 8527 24565 8539 24599
rect 8846 24596 8852 24608
rect 8807 24568 8852 24596
rect 8481 24559 8539 24565
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 10962 24596 10968 24608
rect 10923 24568 10968 24596
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 12250 24596 12256 24608
rect 12163 24568 12256 24596
rect 12250 24556 12256 24568
rect 12308 24596 12314 24608
rect 12544 24596 12572 24695
rect 12618 24692 12624 24744
rect 12676 24732 12682 24744
rect 15764 24741 15792 24772
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 12676 24704 13461 24732
rect 12676 24692 12682 24704
rect 13449 24701 13461 24704
rect 13495 24701 13507 24735
rect 13449 24695 13507 24701
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24701 15807 24735
rect 15749 24695 15807 24701
rect 14274 24664 14280 24676
rect 14235 24636 14280 24664
rect 14274 24624 14280 24636
rect 14332 24624 14338 24676
rect 14369 24667 14427 24673
rect 14369 24633 14381 24667
rect 14415 24633 14427 24667
rect 14369 24627 14427 24633
rect 12308 24568 12572 24596
rect 12308 24556 12314 24568
rect 13630 24556 13636 24608
rect 13688 24596 13694 24608
rect 14001 24599 14059 24605
rect 14001 24596 14013 24599
rect 13688 24568 14013 24596
rect 13688 24556 13694 24568
rect 14001 24565 14013 24568
rect 14047 24596 14059 24599
rect 14384 24596 14412 24627
rect 14047 24568 14412 24596
rect 14047 24565 14059 24568
rect 14001 24559 14059 24565
rect 14826 24556 14832 24608
rect 14884 24596 14890 24608
rect 15933 24599 15991 24605
rect 15933 24596 15945 24599
rect 14884 24568 15945 24596
rect 14884 24556 14890 24568
rect 15933 24565 15945 24568
rect 15979 24565 15991 24599
rect 16850 24596 16856 24608
rect 16811 24568 16856 24596
rect 15933 24559 15991 24565
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 14550 24392 14556 24404
rect 14511 24364 14556 24392
rect 14550 24352 14556 24364
rect 14608 24352 14614 24404
rect 15930 24352 15936 24404
rect 15988 24392 15994 24404
rect 17037 24395 17095 24401
rect 17037 24392 17049 24395
rect 15988 24364 17049 24392
rect 15988 24352 15994 24364
rect 17037 24361 17049 24364
rect 17083 24361 17095 24395
rect 17037 24355 17095 24361
rect 11422 24324 11428 24336
rect 11383 24296 11428 24324
rect 11422 24284 11428 24296
rect 11480 24284 11486 24336
rect 12250 24284 12256 24336
rect 12308 24324 12314 24336
rect 12989 24327 13047 24333
rect 12989 24324 13001 24327
rect 12308 24296 13001 24324
rect 12308 24284 12314 24296
rect 12989 24293 13001 24296
rect 13035 24293 13047 24327
rect 12989 24287 13047 24293
rect 4154 24265 4160 24268
rect 4132 24259 4160 24265
rect 4132 24256 4144 24259
rect 4067 24228 4144 24256
rect 4132 24225 4144 24228
rect 4212 24256 4218 24268
rect 5442 24256 5448 24268
rect 4212 24228 5448 24256
rect 4132 24219 4160 24225
rect 4154 24216 4160 24219
rect 4212 24216 4218 24228
rect 5442 24216 5448 24228
rect 5500 24216 5506 24268
rect 6546 24216 6552 24268
rect 6604 24265 6610 24268
rect 6604 24259 6642 24265
rect 6630 24225 6642 24259
rect 8110 24256 8116 24268
rect 8071 24228 8116 24256
rect 6604 24219 6642 24225
rect 6604 24216 6610 24219
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 9766 24256 9772 24268
rect 9727 24228 9772 24256
rect 9766 24216 9772 24228
rect 9824 24216 9830 24268
rect 15378 24256 15384 24268
rect 15339 24228 15384 24256
rect 15378 24216 15384 24228
rect 15436 24216 15442 24268
rect 16574 24216 16580 24268
rect 16632 24256 16638 24268
rect 18230 24265 18236 24268
rect 16853 24259 16911 24265
rect 16853 24256 16865 24259
rect 16632 24228 16865 24256
rect 16632 24216 16638 24228
rect 16853 24225 16865 24228
rect 16899 24225 16911 24259
rect 16853 24219 16911 24225
rect 18208 24259 18236 24265
rect 18208 24225 18220 24259
rect 18208 24219 18236 24225
rect 18230 24216 18236 24219
rect 18288 24216 18294 24268
rect 24556 24259 24614 24265
rect 24556 24225 24568 24259
rect 24602 24256 24614 24259
rect 25130 24256 25136 24268
rect 24602 24228 25136 24256
rect 24602 24225 24614 24228
rect 24556 24219 24614 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24188 11391 24191
rect 11606 24188 11612 24200
rect 11379 24160 11612 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 11977 24191 12035 24197
rect 11977 24157 11989 24191
rect 12023 24188 12035 24191
rect 12894 24188 12900 24200
rect 12023 24160 12900 24188
rect 12023 24157 12035 24160
rect 11977 24151 12035 24157
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 13170 24188 13176 24200
rect 13131 24160 13176 24188
rect 13170 24148 13176 24160
rect 13228 24148 13234 24200
rect 14642 24148 14648 24200
rect 14700 24188 14706 24200
rect 15289 24191 15347 24197
rect 15289 24188 15301 24191
rect 14700 24160 15301 24188
rect 14700 24148 14706 24160
rect 15289 24157 15301 24160
rect 15335 24157 15347 24191
rect 15289 24151 15347 24157
rect 12342 24080 12348 24132
rect 12400 24120 12406 24132
rect 13814 24120 13820 24132
rect 12400 24092 13820 24120
rect 12400 24080 12406 24092
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 18279 24123 18337 24129
rect 18279 24120 18291 24123
rect 18012 24092 18291 24120
rect 18012 24080 18018 24092
rect 18279 24089 18291 24092
rect 18325 24089 18337 24123
rect 18279 24083 18337 24089
rect 4203 24055 4261 24061
rect 4203 24021 4215 24055
rect 4249 24052 4261 24055
rect 4890 24052 4896 24064
rect 4249 24024 4896 24052
rect 4249 24021 4261 24024
rect 4203 24015 4261 24021
rect 4890 24012 4896 24024
rect 4948 24012 4954 24064
rect 6687 24055 6745 24061
rect 6687 24021 6699 24055
rect 6733 24052 6745 24055
rect 6822 24052 6828 24064
rect 6733 24024 6828 24052
rect 6733 24021 6745 24024
rect 6687 24015 6745 24021
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 8018 24052 8024 24064
rect 7979 24024 8024 24052
rect 8018 24012 8024 24024
rect 8076 24012 8082 24064
rect 8846 24052 8852 24064
rect 8807 24024 8852 24052
rect 8846 24012 8852 24024
rect 8904 24012 8910 24064
rect 9950 24052 9956 24064
rect 9911 24024 9956 24052
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 12526 24052 12532 24064
rect 12487 24024 12532 24052
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 24627 24055 24685 24061
rect 24627 24052 24639 24055
rect 23624 24024 24639 24052
rect 23624 24012 23630 24024
rect 24627 24021 24639 24024
rect 24673 24021 24685 24055
rect 24627 24015 24685 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 3697 23851 3755 23857
rect 3697 23817 3709 23851
rect 3743 23848 3755 23851
rect 4614 23848 4620 23860
rect 3743 23820 4620 23848
rect 3743 23817 3755 23820
rect 3697 23811 3755 23817
rect 1394 23604 1400 23656
rect 1452 23653 1458 23656
rect 1452 23647 1490 23653
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1452 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 3212 23647 3270 23653
rect 3212 23613 3224 23647
rect 3258 23644 3270 23647
rect 3712 23644 3740 23811
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 5258 23848 5264 23860
rect 5219 23820 5264 23848
rect 5258 23808 5264 23820
rect 5316 23808 5322 23860
rect 6546 23848 6552 23860
rect 6507 23820 6552 23848
rect 6546 23808 6552 23820
rect 6604 23808 6610 23860
rect 7653 23851 7711 23857
rect 7653 23817 7665 23851
rect 7699 23848 7711 23851
rect 7742 23848 7748 23860
rect 7699 23820 7748 23848
rect 7699 23817 7711 23820
rect 7653 23811 7711 23817
rect 7742 23808 7748 23820
rect 7800 23808 7806 23860
rect 9677 23851 9735 23857
rect 9677 23817 9689 23851
rect 9723 23848 9735 23851
rect 9766 23848 9772 23860
rect 9723 23820 9772 23848
rect 9723 23817 9735 23820
rect 9677 23811 9735 23817
rect 9766 23808 9772 23820
rect 9824 23848 9830 23860
rect 11054 23848 11060 23860
rect 9824 23820 11060 23848
rect 9824 23808 9830 23820
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 11333 23851 11391 23857
rect 11333 23817 11345 23851
rect 11379 23848 11391 23851
rect 11422 23848 11428 23860
rect 11379 23820 11428 23848
rect 11379 23817 11391 23820
rect 11333 23811 11391 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 13814 23808 13820 23860
rect 13872 23848 13878 23860
rect 15841 23851 15899 23857
rect 15841 23848 15853 23851
rect 13872 23820 15853 23848
rect 13872 23808 13878 23820
rect 15841 23817 15853 23820
rect 15887 23817 15899 23851
rect 15841 23811 15899 23817
rect 4154 23780 4160 23792
rect 4115 23752 4160 23780
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 3258 23616 3740 23644
rect 4760 23647 4818 23653
rect 3258 23613 3270 23616
rect 3212 23607 3270 23613
rect 4760 23613 4772 23647
rect 4806 23644 4818 23647
rect 5276 23644 5304 23808
rect 8846 23780 8852 23792
rect 8680 23752 8852 23780
rect 8680 23721 8708 23752
rect 8846 23740 8852 23752
rect 8904 23780 8910 23792
rect 8904 23752 10548 23780
rect 8904 23740 8910 23752
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 9122 23712 9128 23724
rect 9083 23684 9128 23712
rect 8665 23675 8723 23681
rect 9122 23672 9128 23684
rect 9180 23672 9186 23724
rect 10520 23721 10548 23752
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 12158 23672 12164 23724
rect 12216 23712 12222 23724
rect 12618 23712 12624 23724
rect 12216 23684 12624 23712
rect 12216 23672 12222 23684
rect 12618 23672 12624 23684
rect 12676 23672 12682 23724
rect 12894 23712 12900 23724
rect 12855 23684 12900 23712
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 14550 23712 14556 23724
rect 14511 23684 14556 23712
rect 14550 23672 14556 23684
rect 14608 23672 14614 23724
rect 14826 23712 14832 23724
rect 14787 23684 14832 23712
rect 14826 23672 14832 23684
rect 14884 23672 14890 23724
rect 4806 23616 5304 23644
rect 7469 23647 7527 23653
rect 4806 23613 4818 23616
rect 4760 23607 4818 23613
rect 7469 23613 7481 23647
rect 7515 23644 7527 23647
rect 8110 23644 8116 23656
rect 7515 23616 7549 23644
rect 8023 23616 8116 23644
rect 7515 23613 7527 23616
rect 7469 23607 7527 23613
rect 1452 23604 1458 23607
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 2682 23576 2688 23588
rect 1581 23548 2688 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 2682 23536 2688 23548
rect 2740 23536 2746 23588
rect 4847 23579 4905 23585
rect 4847 23545 4859 23579
rect 4893 23576 4905 23579
rect 5258 23576 5264 23588
rect 4893 23548 5264 23576
rect 4893 23545 4905 23548
rect 4847 23539 4905 23545
rect 5258 23536 5264 23548
rect 5316 23536 5322 23588
rect 7377 23579 7435 23585
rect 7377 23545 7389 23579
rect 7423 23576 7435 23579
rect 7484 23576 7512 23607
rect 8110 23604 8116 23616
rect 8168 23644 8174 23656
rect 8478 23644 8484 23656
rect 8168 23616 8484 23644
rect 8168 23604 8174 23616
rect 8478 23604 8484 23616
rect 8536 23604 8542 23656
rect 11606 23644 11612 23656
rect 11567 23616 11612 23644
rect 11606 23604 11612 23616
rect 11664 23604 11670 23656
rect 15856 23644 15884 23811
rect 18230 23808 18236 23860
rect 18288 23848 18294 23860
rect 18509 23851 18567 23857
rect 18509 23848 18521 23851
rect 18288 23820 18521 23848
rect 18288 23808 18294 23820
rect 18509 23817 18521 23820
rect 18555 23817 18567 23851
rect 18966 23848 18972 23860
rect 18927 23820 18972 23848
rect 18509 23811 18567 23817
rect 18966 23808 18972 23820
rect 19024 23808 19030 23860
rect 19797 23851 19855 23857
rect 19797 23817 19809 23851
rect 19843 23848 19855 23851
rect 21174 23848 21180 23860
rect 19843 23820 21180 23848
rect 19843 23817 19855 23820
rect 19797 23811 19855 23817
rect 16117 23647 16175 23653
rect 16117 23644 16129 23647
rect 15856 23616 16129 23644
rect 16117 23613 16129 23616
rect 16163 23613 16175 23647
rect 16117 23607 16175 23613
rect 18116 23647 18174 23653
rect 18116 23613 18128 23647
rect 18162 23644 18174 23647
rect 18966 23644 18972 23656
rect 18162 23616 18972 23644
rect 18162 23613 18174 23616
rect 18116 23607 18174 23613
rect 18966 23604 18972 23616
rect 19024 23604 19030 23656
rect 19312 23647 19370 23653
rect 19312 23613 19324 23647
rect 19358 23644 19370 23647
rect 19812 23644 19840 23811
rect 21174 23808 21180 23820
rect 21232 23808 21238 23860
rect 21266 23808 21272 23860
rect 21324 23848 21330 23860
rect 21499 23851 21557 23857
rect 21499 23848 21511 23851
rect 21324 23820 21511 23848
rect 21324 23808 21330 23820
rect 21499 23817 21511 23820
rect 21545 23817 21557 23851
rect 21910 23848 21916 23860
rect 21871 23820 21916 23848
rect 21499 23811 21557 23817
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 25498 23848 25504 23860
rect 25459 23820 25504 23848
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 20901 23783 20959 23789
rect 20901 23749 20913 23783
rect 20947 23780 20959 23783
rect 22002 23780 22008 23792
rect 20947 23752 22008 23780
rect 20947 23749 20959 23752
rect 20901 23743 20959 23749
rect 19358 23616 19840 23644
rect 20416 23647 20474 23653
rect 19358 23613 19370 23616
rect 19312 23607 19370 23613
rect 20416 23613 20428 23647
rect 20462 23644 20474 23647
rect 20916 23644 20944 23743
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 25130 23780 25136 23792
rect 25043 23752 25136 23780
rect 25130 23740 25136 23752
rect 25188 23780 25194 23792
rect 26142 23780 26148 23792
rect 25188 23752 26148 23780
rect 25188 23740 25194 23752
rect 26142 23740 26148 23752
rect 26200 23740 26206 23792
rect 20462 23616 20944 23644
rect 21428 23647 21486 23653
rect 20462 23613 20474 23616
rect 20416 23607 20474 23613
rect 21428 23613 21440 23647
rect 21474 23644 21486 23647
rect 21910 23644 21916 23656
rect 21474 23616 21916 23644
rect 21474 23613 21486 23616
rect 21428 23607 21486 23613
rect 21910 23604 21916 23616
rect 21968 23604 21974 23656
rect 24648 23647 24706 23653
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 25498 23644 25504 23656
rect 24694 23616 25504 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 8386 23576 8392 23588
rect 7423 23548 8392 23576
rect 7423 23545 7435 23548
rect 7377 23539 7435 23545
rect 8386 23536 8392 23548
rect 8444 23536 8450 23588
rect 8757 23579 8815 23585
rect 8757 23545 8769 23579
rect 8803 23545 8815 23579
rect 8757 23539 8815 23545
rect 10229 23579 10287 23585
rect 10229 23545 10241 23579
rect 10275 23545 10287 23579
rect 10229 23539 10287 23545
rect 3142 23468 3148 23520
rect 3200 23508 3206 23520
rect 3283 23511 3341 23517
rect 3283 23508 3295 23511
rect 3200 23480 3295 23508
rect 3200 23468 3206 23480
rect 3283 23477 3295 23480
rect 3329 23477 3341 23511
rect 3283 23471 3341 23477
rect 8481 23511 8539 23517
rect 8481 23477 8493 23511
rect 8527 23508 8539 23511
rect 8570 23508 8576 23520
rect 8527 23480 8576 23508
rect 8527 23477 8539 23480
rect 8481 23471 8539 23477
rect 8570 23468 8576 23480
rect 8628 23508 8634 23520
rect 8772 23508 8800 23539
rect 8628 23480 8800 23508
rect 8628 23468 8634 23480
rect 9858 23468 9864 23520
rect 9916 23508 9922 23520
rect 9953 23511 10011 23517
rect 9953 23508 9965 23511
rect 9916 23480 9965 23508
rect 9916 23468 9922 23480
rect 9953 23477 9965 23480
rect 9999 23508 10011 23511
rect 10134 23508 10140 23520
rect 9999 23480 10140 23508
rect 9999 23477 10011 23480
rect 9953 23471 10011 23477
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 10244 23508 10272 23539
rect 10318 23536 10324 23588
rect 10376 23576 10382 23588
rect 12526 23576 12532 23588
rect 10376 23548 10421 23576
rect 12487 23548 12532 23576
rect 10376 23536 10382 23548
rect 12526 23536 12532 23548
rect 12584 23536 12590 23588
rect 12618 23536 12624 23588
rect 12676 23576 12682 23588
rect 12676 23548 12721 23576
rect 12676 23536 12682 23548
rect 14642 23536 14648 23588
rect 14700 23576 14706 23588
rect 14700 23548 14745 23576
rect 14700 23536 14706 23548
rect 15194 23536 15200 23588
rect 15252 23576 15258 23588
rect 16025 23579 16083 23585
rect 16025 23576 16037 23579
rect 15252 23548 16037 23576
rect 15252 23536 15258 23548
rect 16025 23545 16037 23548
rect 16071 23545 16083 23579
rect 16025 23539 16083 23545
rect 10778 23508 10784 23520
rect 10244 23480 10784 23508
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 12158 23508 12164 23520
rect 12119 23480 12164 23508
rect 12158 23468 12164 23480
rect 12216 23468 12222 23520
rect 12250 23468 12256 23520
rect 12308 23508 12314 23520
rect 13449 23511 13507 23517
rect 13449 23508 13461 23511
rect 12308 23480 13461 23508
rect 12308 23468 12314 23480
rect 13449 23477 13461 23480
rect 13495 23477 13507 23511
rect 13449 23471 13507 23477
rect 14369 23511 14427 23517
rect 14369 23477 14381 23511
rect 14415 23508 14427 23511
rect 14660 23508 14688 23536
rect 14415 23480 14688 23508
rect 14415 23477 14427 23480
rect 14369 23471 14427 23477
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15436 23480 15485 23508
rect 15436 23468 15442 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17037 23511 17095 23517
rect 17037 23508 17049 23511
rect 16632 23480 17049 23508
rect 16632 23468 16638 23480
rect 17037 23477 17049 23480
rect 17083 23477 17095 23511
rect 17037 23471 17095 23477
rect 17954 23468 17960 23520
rect 18012 23508 18018 23520
rect 18187 23511 18245 23517
rect 18187 23508 18199 23511
rect 18012 23480 18199 23508
rect 18012 23468 18018 23480
rect 18187 23477 18199 23480
rect 18233 23477 18245 23511
rect 18187 23471 18245 23477
rect 19334 23468 19340 23520
rect 19392 23517 19398 23520
rect 19392 23511 19441 23517
rect 19392 23477 19395 23511
rect 19429 23477 19441 23511
rect 19392 23471 19441 23477
rect 19392 23468 19398 23471
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 20487 23511 20545 23517
rect 20487 23508 20499 23511
rect 19576 23480 20499 23508
rect 19576 23468 19582 23480
rect 20487 23477 20499 23480
rect 20533 23477 20545 23511
rect 20487 23471 20545 23477
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 23532 23480 24731 23508
rect 23532 23468 23538 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 9674 23264 9680 23316
rect 9732 23264 9738 23316
rect 10778 23304 10784 23316
rect 10739 23276 10784 23304
rect 10778 23264 10784 23276
rect 10836 23264 10842 23316
rect 12894 23304 12900 23316
rect 12855 23276 12900 23304
rect 12894 23264 12900 23276
rect 12952 23264 12958 23316
rect 15102 23304 15108 23316
rect 13832 23276 15108 23304
rect 6914 23196 6920 23248
rect 6972 23236 6978 23248
rect 7742 23236 7748 23248
rect 6972 23208 7748 23236
rect 6972 23196 6978 23208
rect 7742 23196 7748 23208
rect 7800 23196 7806 23248
rect 7837 23239 7895 23245
rect 7837 23205 7849 23239
rect 7883 23236 7895 23239
rect 8018 23236 8024 23248
rect 7883 23208 8024 23236
rect 7883 23205 7895 23208
rect 7837 23199 7895 23205
rect 8018 23196 8024 23208
rect 8076 23196 8082 23248
rect 8389 23239 8447 23245
rect 8389 23205 8401 23239
rect 8435 23236 8447 23239
rect 8846 23236 8852 23248
rect 8435 23208 8852 23236
rect 8435 23205 8447 23208
rect 8389 23199 8447 23205
rect 8846 23196 8852 23208
rect 8904 23196 8910 23248
rect 9692 23236 9720 23264
rect 9769 23239 9827 23245
rect 9769 23236 9781 23239
rect 9692 23208 9781 23236
rect 9769 23205 9781 23208
rect 9815 23205 9827 23239
rect 9769 23199 9827 23205
rect 9861 23239 9919 23245
rect 9861 23205 9873 23239
rect 9907 23236 9919 23239
rect 9950 23236 9956 23248
rect 9907 23208 9956 23236
rect 9907 23205 9919 23208
rect 9861 23199 9919 23205
rect 9950 23196 9956 23208
rect 10008 23196 10014 23248
rect 11054 23196 11060 23248
rect 11112 23236 11118 23248
rect 11425 23239 11483 23245
rect 11425 23236 11437 23239
rect 11112 23208 11437 23236
rect 11112 23196 11118 23208
rect 11425 23205 11437 23208
rect 11471 23236 11483 23239
rect 11790 23236 11796 23248
rect 11471 23208 11796 23236
rect 11471 23205 11483 23208
rect 11425 23199 11483 23205
rect 11790 23196 11796 23208
rect 11848 23196 11854 23248
rect 13722 23196 13728 23248
rect 13780 23236 13786 23248
rect 13832 23245 13860 23276
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 17034 23264 17040 23316
rect 17092 23304 17098 23316
rect 17313 23307 17371 23313
rect 17313 23304 17325 23307
rect 17092 23276 17325 23304
rect 17092 23264 17098 23276
rect 17313 23273 17325 23276
rect 17359 23273 17371 23307
rect 17313 23267 17371 23273
rect 13817 23239 13875 23245
rect 13817 23236 13829 23239
rect 13780 23208 13829 23236
rect 13780 23196 13786 23208
rect 13817 23205 13829 23208
rect 13863 23205 13875 23239
rect 14366 23236 14372 23248
rect 14327 23208 14372 23236
rect 13817 23199 13875 23205
rect 14366 23196 14372 23208
rect 14424 23196 14430 23248
rect 15286 23196 15292 23248
rect 15344 23236 15350 23248
rect 15749 23239 15807 23245
rect 15749 23236 15761 23239
rect 15344 23208 15761 23236
rect 15344 23196 15350 23208
rect 15749 23205 15761 23208
rect 15795 23205 15807 23239
rect 15749 23199 15807 23205
rect 1464 23171 1522 23177
rect 1464 23137 1476 23171
rect 1510 23168 1522 23171
rect 2038 23168 2044 23180
rect 1510 23140 2044 23168
rect 1510 23137 1522 23140
rect 1464 23131 1522 23137
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2476 23171 2534 23177
rect 2476 23137 2488 23171
rect 2522 23168 2534 23171
rect 2774 23168 2780 23180
rect 2522 23140 2780 23168
rect 2522 23137 2534 23140
rect 2476 23131 2534 23137
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 5626 23168 5632 23180
rect 5587 23140 5632 23168
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 6708 23171 6766 23177
rect 6708 23137 6720 23171
rect 6754 23168 6766 23171
rect 7098 23168 7104 23180
rect 6754 23140 7104 23168
rect 6754 23137 6766 23140
rect 6708 23131 6766 23137
rect 7098 23128 7104 23140
rect 7156 23168 7162 23180
rect 7558 23168 7564 23180
rect 7156 23140 7564 23168
rect 7156 23128 7162 23140
rect 7558 23128 7564 23140
rect 7616 23128 7622 23180
rect 12526 23168 12532 23180
rect 12487 23140 12532 23168
rect 12526 23128 12532 23140
rect 12584 23128 12590 23180
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23137 17187 23171
rect 17129 23131 17187 23137
rect 18284 23171 18342 23177
rect 18284 23137 18296 23171
rect 18330 23168 18342 23171
rect 18506 23168 18512 23180
rect 18330 23140 18512 23168
rect 18330 23137 18342 23140
rect 18284 23131 18342 23137
rect 11330 23100 11336 23112
rect 11291 23072 11336 23100
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 11609 23103 11667 23109
rect 11609 23069 11621 23103
rect 11655 23069 11667 23103
rect 11609 23063 11667 23069
rect 10321 23035 10379 23041
rect 10321 23001 10333 23035
rect 10367 23032 10379 23035
rect 10870 23032 10876 23044
rect 10367 23004 10876 23032
rect 10367 23001 10379 23004
rect 10321 22995 10379 23001
rect 10870 22992 10876 23004
rect 10928 23032 10934 23044
rect 11149 23035 11207 23041
rect 11149 23032 11161 23035
rect 10928 23004 11161 23032
rect 10928 22992 10934 23004
rect 11149 23001 11161 23004
rect 11195 23032 11207 23035
rect 11624 23032 11652 23063
rect 13538 23060 13544 23112
rect 13596 23100 13602 23112
rect 13725 23103 13783 23109
rect 13725 23100 13737 23103
rect 13596 23072 13737 23100
rect 13596 23060 13602 23072
rect 13725 23069 13737 23072
rect 13771 23069 13783 23103
rect 13725 23063 13783 23069
rect 15657 23103 15715 23109
rect 15657 23069 15669 23103
rect 15703 23069 15715 23103
rect 16298 23100 16304 23112
rect 16259 23072 16304 23100
rect 15657 23063 15715 23069
rect 11195 23004 11652 23032
rect 11195 23001 11207 23004
rect 11149 22995 11207 23001
rect 15562 22992 15568 23044
rect 15620 23032 15626 23044
rect 15672 23032 15700 23063
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 17144 23100 17172 23131
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 17218 23100 17224 23112
rect 17131 23072 17224 23100
rect 17218 23060 17224 23072
rect 17276 23100 17282 23112
rect 18371 23103 18429 23109
rect 18371 23100 18383 23103
rect 17276 23072 18383 23100
rect 17276 23060 17282 23072
rect 18371 23069 18383 23072
rect 18417 23069 18429 23103
rect 18371 23063 18429 23069
rect 15620 23004 15700 23032
rect 15620 22992 15626 23004
rect 1578 22973 1584 22976
rect 1535 22967 1584 22973
rect 1535 22933 1547 22967
rect 1581 22933 1584 22967
rect 1535 22927 1584 22933
rect 1578 22924 1584 22927
rect 1636 22924 1642 22976
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 2547 22967 2605 22973
rect 2547 22964 2559 22967
rect 1728 22936 2559 22964
rect 1728 22924 1734 22936
rect 2547 22933 2559 22936
rect 2593 22933 2605 22967
rect 2547 22927 2605 22933
rect 6086 22924 6092 22976
rect 6144 22964 6150 22976
rect 6779 22967 6837 22973
rect 6779 22964 6791 22967
rect 6144 22936 6791 22964
rect 6144 22924 6150 22936
rect 6779 22933 6791 22936
rect 6825 22933 6837 22967
rect 8662 22964 8668 22976
rect 8623 22936 8668 22964
rect 6779 22927 6837 22933
rect 8662 22924 8668 22936
rect 8720 22924 8726 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 3237 22763 3295 22769
rect 3237 22760 3249 22763
rect 2832 22732 3249 22760
rect 2832 22720 2838 22732
rect 3237 22729 3249 22732
rect 3283 22729 3295 22763
rect 7098 22760 7104 22772
rect 7059 22732 7104 22760
rect 3237 22723 3295 22729
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 8018 22760 8024 22772
rect 7979 22732 8024 22760
rect 8018 22720 8024 22732
rect 8076 22720 8082 22772
rect 9769 22763 9827 22769
rect 9769 22729 9781 22763
rect 9815 22760 9827 22763
rect 9950 22760 9956 22772
rect 9815 22732 9956 22760
rect 9815 22729 9827 22732
rect 9769 22723 9827 22729
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 11790 22760 11796 22772
rect 11751 22732 11796 22760
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12434 22760 12440 22772
rect 12299 22732 12440 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 13722 22760 13728 22772
rect 13683 22732 13728 22760
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 17218 22760 17224 22772
rect 17179 22732 17224 22760
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 9122 22692 9128 22704
rect 9083 22664 9128 22692
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 9674 22652 9680 22704
rect 9732 22692 9738 22704
rect 10045 22695 10103 22701
rect 10045 22692 10057 22695
rect 9732 22664 10057 22692
rect 9732 22652 9738 22664
rect 10045 22661 10057 22664
rect 10091 22661 10103 22695
rect 10045 22655 10103 22661
rect 2866 22584 2872 22636
rect 2924 22624 2930 22636
rect 3559 22627 3617 22633
rect 3559 22624 3571 22627
rect 2924 22596 3571 22624
rect 2924 22584 2930 22596
rect 3559 22593 3571 22596
rect 3605 22593 3617 22627
rect 3559 22587 3617 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22624 7527 22627
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 7515 22596 8585 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 8573 22593 8585 22596
rect 8619 22624 8631 22627
rect 8662 22624 8668 22636
rect 8619 22596 8668 22624
rect 8619 22593 8631 22596
rect 8573 22587 8631 22593
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 10597 22627 10655 22633
rect 10597 22624 10609 22627
rect 9824 22596 10609 22624
rect 9824 22584 9830 22596
rect 10597 22593 10609 22596
rect 10643 22593 10655 22627
rect 10870 22624 10876 22636
rect 10831 22596 10876 22624
rect 10597 22587 10655 22593
rect 1394 22516 1400 22568
rect 1452 22565 1458 22568
rect 1452 22559 1490 22565
rect 1478 22556 1490 22559
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 1478 22528 2237 22556
rect 1478 22525 1490 22528
rect 1452 22519 1490 22525
rect 2225 22525 2237 22528
rect 2271 22525 2283 22559
rect 2225 22519 2283 22525
rect 2476 22559 2534 22565
rect 2476 22525 2488 22559
rect 2522 22556 2534 22559
rect 2522 22528 3004 22556
rect 2522 22525 2534 22528
rect 2476 22519 2534 22525
rect 1452 22516 1458 22519
rect 1535 22491 1593 22497
rect 1535 22457 1547 22491
rect 1581 22488 1593 22491
rect 2682 22488 2688 22500
rect 1581 22460 2688 22488
rect 1581 22457 1593 22460
rect 1535 22451 1593 22457
rect 2682 22448 2688 22460
rect 2740 22448 2746 22500
rect 1949 22423 2007 22429
rect 1949 22389 1961 22423
rect 1995 22420 2007 22423
rect 2038 22420 2044 22432
rect 1995 22392 2044 22420
rect 1995 22389 2007 22392
rect 1949 22383 2007 22389
rect 2038 22380 2044 22392
rect 2096 22380 2102 22432
rect 2406 22380 2412 22432
rect 2464 22420 2470 22432
rect 2976 22429 3004 22528
rect 3326 22516 3332 22568
rect 3384 22556 3390 22568
rect 3456 22559 3514 22565
rect 3456 22556 3468 22559
rect 3384 22528 3468 22556
rect 3384 22516 3390 22528
rect 3456 22525 3468 22528
rect 3502 22556 3514 22559
rect 3881 22559 3939 22565
rect 3881 22556 3893 22559
rect 3502 22528 3893 22556
rect 3502 22525 3514 22528
rect 3456 22519 3514 22525
rect 3881 22525 3893 22528
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 8665 22491 8723 22497
rect 8665 22457 8677 22491
rect 8711 22457 8723 22491
rect 10612 22488 10640 22587
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 12526 22624 12532 22636
rect 12487 22596 12532 22624
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 12618 22584 12624 22636
rect 12676 22624 12682 22636
rect 13170 22624 13176 22636
rect 12676 22596 13176 22624
rect 12676 22584 12682 22596
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 14826 22624 14832 22636
rect 14787 22596 14832 22624
rect 14826 22584 14832 22596
rect 14884 22584 14890 22636
rect 16206 22624 16212 22636
rect 16167 22596 16212 22624
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 16298 22584 16304 22636
rect 16356 22624 16362 22636
rect 16485 22627 16543 22633
rect 16485 22624 16497 22627
rect 16356 22596 16497 22624
rect 16356 22584 16362 22596
rect 16485 22593 16497 22596
rect 16531 22593 16543 22627
rect 16485 22587 16543 22593
rect 10870 22488 10876 22500
rect 10612 22460 10876 22488
rect 8665 22451 8723 22457
rect 2547 22423 2605 22429
rect 2547 22420 2559 22423
rect 2464 22392 2559 22420
rect 2464 22380 2470 22392
rect 2547 22389 2559 22392
rect 2593 22389 2605 22423
rect 2547 22383 2605 22389
rect 2961 22423 3019 22429
rect 2961 22389 2973 22423
rect 3007 22420 3019 22423
rect 3510 22420 3516 22432
rect 3007 22392 3516 22420
rect 3007 22389 3019 22392
rect 2961 22383 3019 22389
rect 3510 22380 3516 22392
rect 3568 22380 3574 22432
rect 8294 22420 8300 22432
rect 8255 22392 8300 22420
rect 8294 22380 8300 22392
rect 8352 22420 8358 22432
rect 8680 22420 8708 22451
rect 10870 22448 10876 22460
rect 10928 22488 10934 22500
rect 10965 22491 11023 22497
rect 10965 22488 10977 22491
rect 10928 22460 10977 22488
rect 10928 22448 10934 22460
rect 10965 22457 10977 22460
rect 11011 22457 11023 22491
rect 10965 22451 11023 22457
rect 11517 22491 11575 22497
rect 11517 22457 11529 22491
rect 11563 22488 11575 22491
rect 11606 22488 11612 22500
rect 11563 22460 11612 22488
rect 11563 22457 11575 22460
rect 11517 22451 11575 22457
rect 11606 22448 11612 22460
rect 11664 22448 11670 22500
rect 12621 22491 12679 22497
rect 12621 22457 12633 22491
rect 12667 22457 12679 22491
rect 14458 22488 14464 22500
rect 14371 22460 14464 22488
rect 12621 22451 12679 22457
rect 8352 22392 8708 22420
rect 8352 22380 8358 22392
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12636 22420 12664 22451
rect 14458 22448 14464 22460
rect 14516 22448 14522 22500
rect 15654 22448 15660 22500
rect 15712 22488 15718 22500
rect 16025 22491 16083 22497
rect 16025 22488 16037 22491
rect 15712 22460 16037 22488
rect 15712 22448 15718 22460
rect 16025 22457 16037 22460
rect 16071 22488 16083 22491
rect 16301 22491 16359 22497
rect 16301 22488 16313 22491
rect 16071 22460 16313 22488
rect 16071 22457 16083 22460
rect 16025 22451 16083 22457
rect 16301 22457 16313 22460
rect 16347 22457 16359 22491
rect 16301 22451 16359 22457
rect 12492 22392 12664 22420
rect 12492 22380 12498 22392
rect 13906 22380 13912 22432
rect 13964 22420 13970 22432
rect 14093 22423 14151 22429
rect 14093 22420 14105 22423
rect 13964 22392 14105 22420
rect 13964 22380 13970 22392
rect 14093 22389 14105 22392
rect 14139 22420 14151 22423
rect 14476 22420 14504 22448
rect 14139 22392 14504 22420
rect 14139 22389 14151 22392
rect 14093 22383 14151 22389
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 15565 22423 15623 22429
rect 15565 22420 15577 22423
rect 15344 22392 15577 22420
rect 15344 22380 15350 22392
rect 15565 22389 15577 22392
rect 15611 22389 15623 22423
rect 18046 22420 18052 22432
rect 18007 22392 18052 22420
rect 15565 22383 15623 22389
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 18506 22420 18512 22432
rect 18467 22392 18512 22420
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 7742 22216 7748 22228
rect 7703 22188 7748 22216
rect 7742 22176 7748 22188
rect 7800 22176 7806 22228
rect 8294 22216 8300 22228
rect 8255 22188 8300 22216
rect 8294 22176 8300 22188
rect 8352 22176 8358 22228
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 11882 22216 11888 22228
rect 11388 22188 11888 22216
rect 11388 22176 11394 22188
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 13633 22219 13691 22225
rect 13633 22216 13645 22219
rect 13596 22188 13645 22216
rect 13596 22176 13602 22188
rect 13633 22185 13645 22188
rect 13679 22185 13691 22219
rect 13633 22179 13691 22185
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 14645 22219 14703 22225
rect 14645 22216 14657 22219
rect 14424 22188 14657 22216
rect 14424 22176 14430 22188
rect 14645 22185 14657 22188
rect 14691 22185 14703 22219
rect 16206 22216 16212 22228
rect 16167 22188 16212 22216
rect 14645 22179 14703 22185
rect 16206 22176 16212 22188
rect 16264 22176 16270 22228
rect 11054 22148 11060 22160
rect 11015 22120 11060 22148
rect 11054 22108 11060 22120
rect 11112 22108 11118 22160
rect 11606 22148 11612 22160
rect 11567 22120 11612 22148
rect 11606 22108 11612 22120
rect 11664 22108 11670 22160
rect 13173 22151 13231 22157
rect 13173 22117 13185 22151
rect 13219 22148 13231 22151
rect 13814 22148 13820 22160
rect 13219 22120 13820 22148
rect 13219 22117 13231 22120
rect 13173 22111 13231 22117
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 16482 22148 16488 22160
rect 16443 22120 16488 22148
rect 16482 22108 16488 22120
rect 16540 22148 16546 22160
rect 17865 22151 17923 22157
rect 17865 22148 17877 22151
rect 16540 22120 17877 22148
rect 16540 22108 16546 22120
rect 17865 22117 17877 22120
rect 17911 22117 17923 22151
rect 17865 22111 17923 22117
rect 2016 22083 2074 22089
rect 2016 22049 2028 22083
rect 2062 22080 2074 22083
rect 2314 22080 2320 22092
rect 2062 22052 2320 22080
rect 2062 22049 2074 22052
rect 2016 22043 2074 22049
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 3050 22089 3056 22092
rect 3028 22083 3056 22089
rect 3028 22049 3040 22083
rect 3028 22043 3056 22049
rect 3050 22040 3056 22043
rect 3108 22040 3114 22092
rect 5997 22083 6055 22089
rect 5997 22049 6009 22083
rect 6043 22080 6055 22083
rect 6546 22080 6552 22092
rect 6043 22052 6552 22080
rect 6043 22049 6055 22052
rect 5997 22043 6055 22049
rect 6546 22040 6552 22052
rect 6604 22040 6610 22092
rect 7076 22083 7134 22089
rect 7076 22049 7088 22083
rect 7122 22080 7134 22083
rect 7466 22080 7472 22092
rect 7122 22052 7472 22080
rect 7122 22049 7134 22052
rect 7076 22043 7134 22049
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 8570 22080 8576 22092
rect 8531 22052 8576 22080
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 9928 22083 9986 22089
rect 9928 22049 9940 22083
rect 9974 22080 9986 22083
rect 9974 22052 10456 22080
rect 9974 22049 9986 22052
rect 9928 22043 9986 22049
rect 7147 21947 7205 21953
rect 7147 21913 7159 21947
rect 7193 21944 7205 21947
rect 8202 21944 8208 21956
rect 7193 21916 8208 21944
rect 7193 21913 7205 21916
rect 7147 21907 7205 21913
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 10042 21953 10048 21956
rect 9999 21947 10048 21953
rect 9999 21913 10011 21947
rect 10045 21913 10048 21947
rect 9999 21907 10048 21913
rect 10042 21904 10048 21907
rect 10100 21904 10106 21956
rect 10428 21953 10456 22052
rect 12434 22040 12440 22092
rect 12492 22080 12498 22092
rect 12986 22080 12992 22092
rect 12492 22052 12537 22080
rect 12947 22052 12992 22080
rect 12492 22040 12498 22052
rect 12986 22040 12992 22052
rect 13044 22040 13050 22092
rect 14182 22040 14188 22092
rect 14240 22089 14246 22092
rect 14240 22083 14278 22089
rect 14266 22049 14278 22083
rect 14240 22043 14278 22049
rect 14323 22083 14381 22089
rect 14323 22049 14335 22083
rect 14369 22080 14381 22083
rect 14734 22080 14740 22092
rect 14369 22052 14740 22080
rect 14369 22049 14381 22052
rect 14323 22043 14381 22049
rect 14240 22040 14246 22043
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 15470 22089 15476 22092
rect 15324 22083 15382 22089
rect 15324 22080 15336 22083
rect 15304 22049 15336 22080
rect 15370 22049 15382 22083
rect 15304 22043 15382 22049
rect 15427 22083 15476 22089
rect 15427 22049 15439 22083
rect 15473 22049 15476 22083
rect 15427 22043 15476 22049
rect 10778 21972 10784 22024
rect 10836 22012 10842 22024
rect 10965 22015 11023 22021
rect 10965 22012 10977 22015
rect 10836 21984 10977 22012
rect 10836 21972 10842 21984
rect 10965 21981 10977 21984
rect 11011 21981 11023 22015
rect 15304 22012 15332 22043
rect 15470 22040 15476 22043
rect 15528 22040 15534 22092
rect 18230 22080 18236 22092
rect 18191 22052 18236 22080
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 15304 21984 15424 22012
rect 10965 21975 11023 21981
rect 15396 21956 15424 21984
rect 16022 21972 16028 22024
rect 16080 22012 16086 22024
rect 16390 22012 16396 22024
rect 16080 21984 16396 22012
rect 16080 21972 16086 21984
rect 16390 21972 16396 21984
rect 16448 21972 16454 22024
rect 16666 22012 16672 22024
rect 16627 21984 16672 22012
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 10413 21947 10471 21953
rect 10413 21913 10425 21947
rect 10459 21944 10471 21947
rect 11606 21944 11612 21956
rect 10459 21916 11612 21944
rect 10459 21913 10471 21916
rect 10413 21907 10471 21913
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 15378 21904 15384 21956
rect 15436 21904 15442 21956
rect 2130 21885 2136 21888
rect 2087 21879 2136 21885
rect 2087 21845 2099 21879
rect 2133 21845 2136 21879
rect 2087 21839 2136 21845
rect 2130 21836 2136 21839
rect 2188 21836 2194 21888
rect 3099 21879 3157 21885
rect 3099 21845 3111 21879
rect 3145 21876 3157 21879
rect 3970 21876 3976 21888
rect 3145 21848 3976 21876
rect 3145 21845 3157 21848
rect 3099 21839 3157 21845
rect 3970 21836 3976 21848
rect 4028 21836 4034 21888
rect 6178 21876 6184 21888
rect 6139 21848 6184 21876
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 15562 21836 15568 21888
rect 15620 21876 15626 21888
rect 15749 21879 15807 21885
rect 15749 21876 15761 21879
rect 15620 21848 15761 21876
rect 15620 21836 15626 21848
rect 15749 21845 15761 21848
rect 15795 21845 15807 21879
rect 15749 21839 15807 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 6546 21672 6552 21684
rect 6507 21644 6552 21672
rect 6546 21632 6552 21644
rect 6604 21632 6610 21684
rect 8570 21632 8576 21684
rect 8628 21672 8634 21684
rect 8941 21675 8999 21681
rect 8941 21672 8953 21675
rect 8628 21644 8953 21672
rect 8628 21632 8634 21644
rect 8941 21641 8953 21644
rect 8987 21641 8999 21675
rect 8941 21635 8999 21641
rect 9122 21632 9128 21684
rect 9180 21672 9186 21684
rect 9309 21675 9367 21681
rect 9309 21672 9321 21675
rect 9180 21644 9321 21672
rect 9180 21632 9186 21644
rect 9309 21641 9321 21644
rect 9355 21641 9367 21675
rect 9309 21635 9367 21641
rect 10689 21675 10747 21681
rect 10689 21641 10701 21675
rect 10735 21672 10747 21675
rect 10962 21672 10968 21684
rect 10735 21644 10968 21672
rect 10735 21641 10747 21644
rect 10689 21635 10747 21641
rect 1946 21564 1952 21616
rect 2004 21604 2010 21616
rect 2547 21607 2605 21613
rect 2547 21604 2559 21607
rect 2004 21576 2559 21604
rect 2004 21564 2010 21576
rect 2547 21573 2559 21576
rect 2593 21573 2605 21607
rect 2547 21567 2605 21573
rect 5905 21607 5963 21613
rect 5905 21573 5917 21607
rect 5951 21604 5963 21607
rect 5951 21576 7144 21604
rect 5951 21573 5963 21576
rect 5905 21567 5963 21573
rect 6914 21496 6920 21548
rect 6972 21536 6978 21548
rect 6972 21508 7017 21536
rect 6972 21496 6978 21508
rect 1394 21428 1400 21480
rect 1452 21477 1458 21480
rect 2498 21477 2504 21480
rect 1452 21471 1490 21477
rect 1478 21468 1490 21471
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1478 21440 1869 21468
rect 1478 21437 1490 21440
rect 1452 21431 1490 21437
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 2476 21471 2504 21477
rect 2476 21437 2488 21471
rect 2556 21468 2562 21480
rect 2869 21471 2927 21477
rect 2869 21468 2881 21471
rect 2556 21440 2881 21468
rect 2476 21431 2504 21437
rect 1452 21428 1458 21431
rect 2498 21428 2504 21431
rect 2556 21428 2562 21440
rect 2869 21437 2881 21440
rect 2915 21437 2927 21471
rect 2869 21431 2927 21437
rect 3418 21428 3424 21480
rect 3476 21477 3482 21480
rect 3476 21471 3514 21477
rect 3502 21468 3514 21471
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3502 21440 3893 21468
rect 3502 21437 3514 21440
rect 3476 21431 3514 21437
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 3881 21431 3939 21437
rect 3476 21428 3482 21431
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 4468 21471 4526 21477
rect 4468 21468 4480 21471
rect 4396 21440 4480 21468
rect 4396 21428 4402 21440
rect 4468 21437 4480 21440
rect 4514 21468 4526 21471
rect 4893 21471 4951 21477
rect 4893 21468 4905 21471
rect 4514 21440 4905 21468
rect 4514 21437 4526 21440
rect 4468 21431 4526 21437
rect 4893 21437 4905 21440
rect 4939 21437 4951 21471
rect 4893 21431 4951 21437
rect 5721 21471 5779 21477
rect 5721 21437 5733 21471
rect 5767 21468 5779 21471
rect 7116 21468 7144 21576
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 7515 21508 8432 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 5767 21440 6040 21468
rect 7116 21440 7849 21468
rect 5767 21437 5779 21440
rect 5721 21431 5779 21437
rect 1535 21403 1593 21409
rect 1535 21369 1547 21403
rect 1581 21400 1593 21403
rect 2682 21400 2688 21412
rect 1581 21372 2688 21400
rect 1581 21369 1593 21372
rect 1535 21363 1593 21369
rect 2682 21360 2688 21372
rect 2740 21360 2746 21412
rect 3559 21403 3617 21409
rect 3559 21369 3571 21403
rect 3605 21400 3617 21403
rect 4154 21400 4160 21412
rect 3605 21372 4160 21400
rect 3605 21369 3617 21372
rect 3559 21363 3617 21369
rect 4154 21360 4160 21372
rect 4212 21360 4218 21412
rect 6012 21344 6040 21440
rect 7837 21437 7849 21440
rect 7883 21468 7895 21471
rect 8202 21468 8208 21480
rect 7883 21440 8208 21468
rect 7883 21437 7895 21440
rect 7837 21431 7895 21437
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 8404 21477 8432 21508
rect 8389 21471 8447 21477
rect 8389 21437 8401 21471
rect 8435 21468 8447 21471
rect 8754 21468 8760 21480
rect 8435 21440 8760 21468
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 9324 21468 9352 21635
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12253 21675 12311 21681
rect 12253 21672 12265 21675
rect 12124 21644 12265 21672
rect 12124 21632 12130 21644
rect 12253 21641 12265 21644
rect 12299 21672 12311 21675
rect 12434 21672 12440 21684
rect 12299 21644 12440 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 12986 21632 12992 21684
rect 13044 21672 13050 21684
rect 13449 21675 13507 21681
rect 13449 21672 13461 21675
rect 13044 21644 13461 21672
rect 13044 21632 13050 21644
rect 13449 21641 13461 21644
rect 13495 21641 13507 21675
rect 14182 21672 14188 21684
rect 14095 21644 14188 21672
rect 13449 21635 13507 21641
rect 14182 21632 14188 21644
rect 14240 21672 14246 21684
rect 14826 21672 14832 21684
rect 14240 21644 14832 21672
rect 14240 21632 14246 21644
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15105 21675 15163 21681
rect 15105 21641 15117 21675
rect 15151 21672 15163 21675
rect 15286 21672 15292 21684
rect 15151 21644 15292 21672
rect 15151 21641 15163 21644
rect 15105 21635 15163 21641
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 15749 21675 15807 21681
rect 15749 21641 15761 21675
rect 15795 21672 15807 21675
rect 16022 21672 16028 21684
rect 15795 21644 16028 21672
rect 15795 21641 15807 21644
rect 15749 21635 15807 21641
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 16117 21675 16175 21681
rect 16117 21641 16129 21675
rect 16163 21672 16175 21675
rect 16482 21672 16488 21684
rect 16163 21644 16488 21672
rect 16163 21641 16175 21644
rect 16117 21635 16175 21641
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 18230 21672 18236 21684
rect 18191 21644 18236 21672
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 12802 21604 12808 21616
rect 10980 21576 12808 21604
rect 9528 21471 9586 21477
rect 9528 21468 9540 21471
rect 9324 21440 9540 21468
rect 9528 21437 9540 21440
rect 9574 21437 9586 21471
rect 9528 21431 9586 21437
rect 10042 21428 10048 21480
rect 10100 21468 10106 21480
rect 10980 21477 11008 21576
rect 12802 21564 12808 21576
rect 12860 21564 12866 21616
rect 13004 21536 13032 21632
rect 15378 21564 15384 21616
rect 15436 21604 15442 21616
rect 16666 21604 16672 21616
rect 15436 21576 16672 21604
rect 15436 21564 15442 21576
rect 16666 21564 16672 21576
rect 16724 21604 16730 21616
rect 16853 21607 16911 21613
rect 16853 21604 16865 21607
rect 16724 21576 16865 21604
rect 16724 21564 16730 21576
rect 16853 21573 16865 21576
rect 16899 21573 16911 21607
rect 16853 21567 16911 21573
rect 16298 21536 16304 21548
rect 11440 21508 13032 21536
rect 16259 21508 16304 21536
rect 11440 21480 11468 21508
rect 16298 21496 16304 21508
rect 16356 21536 16362 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 16356 21508 17233 21536
rect 16356 21496 16362 21508
rect 17221 21505 17233 21508
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 10321 21471 10379 21477
rect 10321 21468 10333 21471
rect 10100 21440 10333 21468
rect 10100 21428 10106 21440
rect 10321 21437 10333 21440
rect 10367 21468 10379 21471
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 10367 21440 10977 21468
rect 10367 21437 10379 21440
rect 10321 21431 10379 21437
rect 10965 21437 10977 21440
rect 11011 21437 11023 21471
rect 10965 21431 11023 21437
rect 11333 21471 11391 21477
rect 11333 21437 11345 21471
rect 11379 21468 11391 21471
rect 11422 21468 11428 21480
rect 11379 21440 11428 21468
rect 11379 21437 11391 21440
rect 11333 21431 11391 21437
rect 11422 21428 11428 21440
rect 11480 21428 11486 21480
rect 12713 21471 12771 21477
rect 12713 21437 12725 21471
rect 12759 21468 12771 21471
rect 12802 21468 12808 21480
rect 12759 21440 12808 21468
rect 12759 21437 12771 21440
rect 12713 21431 12771 21437
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 12897 21471 12955 21477
rect 12897 21437 12909 21471
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 14642 21468 14648 21480
rect 14599 21440 14648 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 11514 21400 11520 21412
rect 11475 21372 11520 21400
rect 11514 21360 11520 21372
rect 11572 21360 11578 21412
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 12618 21400 12624 21412
rect 11931 21372 12624 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 12618 21360 12624 21372
rect 12676 21400 12682 21412
rect 12912 21400 12940 21431
rect 14642 21428 14648 21440
rect 14700 21468 14706 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 14700 21440 15301 21468
rect 14700 21428 14706 21440
rect 15289 21437 15301 21440
rect 15335 21468 15347 21471
rect 15654 21468 15660 21480
rect 15335 21440 15660 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 15654 21428 15660 21440
rect 15712 21428 15718 21480
rect 12676 21372 12940 21400
rect 16393 21403 16451 21409
rect 12676 21360 12682 21372
rect 16393 21369 16405 21403
rect 16439 21369 16451 21403
rect 16393 21363 16451 21369
rect 2314 21332 2320 21344
rect 2275 21304 2320 21332
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3237 21335 3295 21341
rect 3237 21332 3249 21335
rect 3108 21304 3249 21332
rect 3108 21292 3114 21304
rect 3237 21301 3249 21304
rect 3283 21301 3295 21335
rect 3237 21295 3295 21301
rect 4571 21335 4629 21341
rect 4571 21301 4583 21335
rect 4617 21332 4629 21335
rect 5442 21332 5448 21344
rect 4617 21304 5448 21332
rect 4617 21301 4629 21304
rect 4571 21295 4629 21301
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 5994 21292 6000 21344
rect 6052 21332 6058 21344
rect 6181 21335 6239 21341
rect 6181 21332 6193 21335
rect 6052 21304 6193 21332
rect 6052 21292 6058 21304
rect 6181 21301 6193 21304
rect 6227 21301 6239 21335
rect 8018 21332 8024 21344
rect 7979 21304 8024 21332
rect 6181 21295 6239 21301
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 8386 21292 8392 21344
rect 8444 21332 8450 21344
rect 9631 21335 9689 21341
rect 9631 21332 9643 21335
rect 8444 21304 9643 21332
rect 8444 21292 8450 21304
rect 9631 21301 9643 21304
rect 9677 21301 9689 21335
rect 12710 21332 12716 21344
rect 12671 21304 12716 21332
rect 9631 21295 9689 21301
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 16408 21332 16436 21363
rect 16574 21332 16580 21344
rect 16408 21304 16580 21332
rect 16574 21292 16580 21304
rect 16632 21332 16638 21344
rect 18230 21332 18236 21344
rect 16632 21304 18236 21332
rect 16632 21292 16638 21304
rect 18230 21292 18236 21304
rect 18288 21292 18294 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 8570 21088 8576 21140
rect 8628 21128 8634 21140
rect 8757 21131 8815 21137
rect 8757 21128 8769 21131
rect 8628 21100 8769 21128
rect 8628 21088 8634 21100
rect 8757 21097 8769 21100
rect 8803 21097 8815 21131
rect 10870 21128 10876 21140
rect 10831 21100 10876 21128
rect 8757 21091 8815 21097
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 11931 21131 11989 21137
rect 11931 21097 11943 21131
rect 11977 21128 11989 21131
rect 12342 21128 12348 21140
rect 11977 21100 12348 21128
rect 11977 21097 11989 21100
rect 11931 21091 11989 21097
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 13630 21088 13636 21140
rect 13688 21128 13694 21140
rect 13725 21131 13783 21137
rect 13725 21128 13737 21131
rect 13688 21100 13737 21128
rect 13688 21088 13694 21100
rect 13725 21097 13737 21100
rect 13771 21097 13783 21131
rect 13998 21128 14004 21140
rect 13959 21100 14004 21128
rect 13725 21091 13783 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 15105 21131 15163 21137
rect 15105 21097 15117 21131
rect 15151 21128 15163 21131
rect 15378 21128 15384 21140
rect 15151 21100 15384 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 16209 21131 16267 21137
rect 16209 21097 16221 21131
rect 16255 21128 16267 21131
rect 16574 21128 16580 21140
rect 16255 21100 16580 21128
rect 16255 21097 16267 21100
rect 16209 21091 16267 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17589 21131 17647 21137
rect 17589 21097 17601 21131
rect 17635 21128 17647 21131
rect 17862 21128 17868 21140
rect 17635 21100 17868 21128
rect 17635 21097 17647 21100
rect 17589 21091 17647 21097
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 6454 21060 6460 21072
rect 6415 21032 6460 21060
rect 6454 21020 6460 21032
rect 6512 21020 6518 21072
rect 8110 21020 8116 21072
rect 8168 21069 8174 21072
rect 8168 21063 8216 21069
rect 8168 21029 8170 21063
rect 8204 21029 8216 21063
rect 8168 21023 8216 21029
rect 10315 21063 10373 21069
rect 10315 21029 10327 21063
rect 10361 21060 10373 21063
rect 10594 21060 10600 21072
rect 10361 21032 10600 21060
rect 10361 21029 10373 21032
rect 10315 21023 10373 21029
rect 8168 21020 8174 21023
rect 10594 21020 10600 21032
rect 10652 21020 10658 21072
rect 10778 21020 10784 21072
rect 10836 21060 10842 21072
rect 11517 21063 11575 21069
rect 11517 21060 11529 21063
rect 10836 21032 11529 21060
rect 10836 21020 10842 21032
rect 11517 21029 11529 21032
rect 11563 21029 11575 21063
rect 11517 21023 11575 21029
rect 13167 21063 13225 21069
rect 13167 21029 13179 21063
rect 13213 21060 13225 21063
rect 13262 21060 13268 21072
rect 13213 21032 13268 21060
rect 13213 21029 13225 21032
rect 13167 21023 13225 21029
rect 13262 21020 13268 21032
rect 13320 21020 13326 21072
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 15610 21063 15668 21069
rect 15610 21060 15622 21063
rect 15528 21032 15622 21060
rect 15528 21020 15534 21032
rect 15610 21029 15622 21032
rect 15656 21029 15668 21063
rect 15610 21023 15668 21029
rect 1394 20952 1400 21004
rect 1452 21001 1458 21004
rect 1452 20995 1490 21001
rect 1478 20961 1490 20995
rect 4706 20992 4712 21004
rect 4667 20964 4712 20992
rect 1452 20955 1490 20961
rect 1452 20952 1458 20955
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 11882 21001 11888 21004
rect 11860 20995 11888 21001
rect 11860 20992 11872 20995
rect 11795 20964 11872 20992
rect 11860 20961 11872 20964
rect 11940 20992 11946 21004
rect 12342 20992 12348 21004
rect 11940 20964 12348 20992
rect 11860 20955 11888 20961
rect 11882 20952 11888 20955
rect 11940 20952 11946 20964
rect 12342 20952 12348 20964
rect 12400 20952 12406 21004
rect 12710 20952 12716 21004
rect 12768 20992 12774 21004
rect 12805 20995 12863 21001
rect 12805 20992 12817 20995
rect 12768 20964 12817 20992
rect 12768 20952 12774 20964
rect 12805 20961 12817 20964
rect 12851 20961 12863 20995
rect 17402 20992 17408 21004
rect 17363 20964 17408 20992
rect 12805 20955 12863 20961
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 1578 20884 1584 20936
rect 1636 20924 1642 20936
rect 2409 20927 2467 20933
rect 2409 20924 2421 20927
rect 1636 20896 2421 20924
rect 1636 20884 1642 20896
rect 2409 20893 2421 20896
rect 2455 20893 2467 20927
rect 6362 20924 6368 20936
rect 6323 20896 6368 20924
rect 2409 20887 2467 20893
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 7837 20927 7895 20933
rect 7837 20893 7849 20927
rect 7883 20893 7895 20927
rect 9950 20924 9956 20936
rect 9911 20896 9956 20924
rect 7837 20887 7895 20893
rect 6917 20859 6975 20865
rect 6917 20825 6929 20859
rect 6963 20825 6975 20859
rect 6917 20819 6975 20825
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 2498 20788 2504 20800
rect 1581 20760 2504 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 2498 20748 2504 20760
rect 2556 20748 2562 20800
rect 4614 20748 4620 20800
rect 4672 20788 4678 20800
rect 4801 20791 4859 20797
rect 4801 20788 4813 20791
rect 4672 20760 4813 20788
rect 4672 20748 4678 20760
rect 4801 20757 4813 20760
rect 4847 20757 4859 20791
rect 6932 20788 6960 20819
rect 7377 20791 7435 20797
rect 7377 20788 7389 20791
rect 6932 20760 7389 20788
rect 4801 20751 4859 20757
rect 7377 20757 7389 20760
rect 7423 20788 7435 20791
rect 7466 20788 7472 20800
rect 7423 20760 7472 20788
rect 7423 20757 7435 20760
rect 7377 20751 7435 20757
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 7745 20791 7803 20797
rect 7745 20757 7757 20791
rect 7791 20788 7803 20791
rect 7852 20788 7880 20887
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 8202 20788 8208 20800
rect 7791 20760 8208 20788
rect 7791 20757 7803 20760
rect 7745 20751 7803 20757
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 11241 20791 11299 20797
rect 11241 20757 11253 20791
rect 11287 20788 11299 20791
rect 11422 20788 11428 20800
rect 11287 20760 11428 20788
rect 11287 20757 11299 20760
rect 11241 20751 11299 20757
rect 11422 20748 11428 20760
rect 11480 20748 11486 20800
rect 12529 20791 12587 20797
rect 12529 20757 12541 20791
rect 12575 20788 12587 20791
rect 12802 20788 12808 20800
rect 12575 20760 12808 20788
rect 12575 20757 12587 20760
rect 12529 20751 12587 20757
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1394 20544 1400 20596
rect 1452 20584 1458 20596
rect 2225 20587 2283 20593
rect 2225 20584 2237 20587
rect 1452 20556 2237 20584
rect 1452 20544 1458 20556
rect 2225 20553 2237 20556
rect 2271 20553 2283 20587
rect 2225 20547 2283 20553
rect 4617 20587 4675 20593
rect 4617 20553 4629 20587
rect 4663 20584 4675 20587
rect 4706 20584 4712 20596
rect 4663 20556 4712 20584
rect 4663 20553 4675 20556
rect 4617 20547 4675 20553
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 8478 20544 8484 20596
rect 8536 20584 8542 20596
rect 8941 20587 8999 20593
rect 8941 20584 8953 20587
rect 8536 20556 8953 20584
rect 8536 20544 8542 20556
rect 8941 20553 8953 20556
rect 8987 20553 8999 20587
rect 8941 20547 8999 20553
rect 10689 20587 10747 20593
rect 10689 20553 10701 20587
rect 10735 20584 10747 20587
rect 10962 20584 10968 20596
rect 10735 20556 10968 20584
rect 10735 20553 10747 20556
rect 10689 20547 10747 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11882 20584 11888 20596
rect 11843 20556 11888 20584
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14921 20587 14979 20593
rect 14921 20584 14933 20587
rect 13872 20556 14933 20584
rect 13872 20544 13878 20556
rect 14921 20553 14933 20556
rect 14967 20584 14979 20587
rect 15286 20584 15292 20596
rect 14967 20556 15292 20584
rect 14967 20553 14979 20556
rect 14921 20547 14979 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 17402 20584 17408 20596
rect 17363 20556 17408 20584
rect 17402 20544 17408 20556
rect 17460 20584 17466 20596
rect 18187 20587 18245 20593
rect 18187 20584 18199 20587
rect 17460 20556 18199 20584
rect 17460 20544 17466 20556
rect 18187 20553 18199 20556
rect 18233 20553 18245 20587
rect 18187 20547 18245 20553
rect 14642 20516 14648 20528
rect 14603 20488 14648 20516
rect 14642 20476 14648 20488
rect 14700 20476 14706 20528
rect 16114 20516 16120 20528
rect 16075 20488 16120 20516
rect 16114 20476 16120 20488
rect 16172 20476 16178 20528
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2682 20448 2688 20460
rect 1995 20420 2688 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 1448 20383 1506 20389
rect 1448 20349 1460 20383
rect 1494 20380 1506 20383
rect 1964 20380 1992 20411
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20448 7619 20451
rect 8018 20448 8024 20460
rect 7607 20420 8024 20448
rect 7607 20417 7619 20420
rect 7561 20411 7619 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 13722 20448 13728 20460
rect 13683 20420 13728 20448
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 15562 20448 15568 20460
rect 15475 20420 15568 20448
rect 15562 20408 15568 20420
rect 15620 20448 15626 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 15620 20420 16865 20448
rect 15620 20408 15626 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 1494 20352 1992 20380
rect 1494 20349 1506 20352
rect 1448 20343 1506 20349
rect 2314 20340 2320 20392
rect 2372 20380 2378 20392
rect 2444 20383 2502 20389
rect 2444 20380 2456 20383
rect 2372 20352 2456 20380
rect 2372 20340 2378 20352
rect 2444 20349 2456 20352
rect 2490 20380 2502 20383
rect 2869 20383 2927 20389
rect 2869 20380 2881 20383
rect 2490 20352 2881 20380
rect 2490 20349 2502 20352
rect 2444 20343 2502 20349
rect 2869 20349 2881 20352
rect 2915 20349 2927 20383
rect 2869 20343 2927 20349
rect 5077 20383 5135 20389
rect 5077 20349 5089 20383
rect 5123 20380 5135 20383
rect 5813 20383 5871 20389
rect 5813 20380 5825 20383
rect 5123 20352 5825 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5813 20349 5825 20352
rect 5859 20380 5871 20383
rect 9766 20380 9772 20392
rect 5859 20352 6408 20380
rect 9679 20352 9772 20380
rect 5859 20349 5871 20352
rect 5813 20343 5871 20349
rect 1535 20315 1593 20321
rect 1535 20281 1547 20315
rect 1581 20312 1593 20315
rect 2222 20312 2228 20324
rect 1581 20284 2228 20312
rect 1581 20281 1593 20284
rect 1535 20275 1593 20281
rect 2222 20272 2228 20284
rect 2280 20272 2286 20324
rect 5902 20312 5908 20324
rect 5863 20284 5908 20312
rect 5902 20272 5908 20284
rect 5960 20272 5966 20324
rect 2547 20247 2605 20253
rect 2547 20213 2559 20247
rect 2593 20244 2605 20247
rect 2682 20244 2688 20256
rect 2593 20216 2688 20244
rect 2593 20213 2605 20216
rect 2547 20207 2605 20213
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 3418 20244 3424 20256
rect 3379 20216 3424 20244
rect 3418 20204 3424 20216
rect 3476 20204 3482 20256
rect 6380 20253 6408 20352
rect 9766 20340 9772 20352
rect 9824 20380 9830 20392
rect 18138 20389 18144 20392
rect 10965 20383 11023 20389
rect 10965 20380 10977 20383
rect 9824 20352 10977 20380
rect 9824 20340 9830 20352
rect 10965 20349 10977 20352
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 18116 20383 18144 20389
rect 18116 20349 18128 20383
rect 18196 20380 18202 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18196 20352 18521 20380
rect 18116 20343 18144 20349
rect 18138 20340 18144 20343
rect 18196 20340 18202 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 7929 20315 7987 20321
rect 7929 20281 7941 20315
rect 7975 20312 7987 20315
rect 8110 20312 8116 20324
rect 7975 20284 8116 20312
rect 7975 20281 7987 20284
rect 7929 20275 7987 20281
rect 8110 20272 8116 20284
rect 8168 20312 8174 20324
rect 8383 20315 8441 20321
rect 8383 20312 8395 20315
rect 8168 20284 8395 20312
rect 8168 20272 8174 20284
rect 8383 20281 8395 20284
rect 8429 20312 8441 20315
rect 9309 20315 9367 20321
rect 9309 20312 9321 20315
rect 8429 20284 9321 20312
rect 8429 20281 8441 20284
rect 8383 20275 8441 20281
rect 9309 20281 9321 20284
rect 9355 20312 9367 20315
rect 9677 20315 9735 20321
rect 9677 20312 9689 20315
rect 9355 20284 9689 20312
rect 9355 20281 9367 20284
rect 9309 20275 9367 20281
rect 9677 20281 9689 20284
rect 9723 20312 9735 20315
rect 10131 20315 10189 20321
rect 10131 20312 10143 20315
rect 9723 20284 10143 20312
rect 9723 20281 9735 20284
rect 9677 20275 9735 20281
rect 10131 20281 10143 20284
rect 10177 20312 10189 20315
rect 10686 20312 10692 20324
rect 10177 20284 10692 20312
rect 10177 20281 10189 20284
rect 10131 20275 10189 20281
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 14087 20315 14145 20321
rect 14087 20281 14099 20315
rect 14133 20281 14145 20315
rect 14087 20275 14145 20281
rect 6365 20247 6423 20253
rect 6365 20213 6377 20247
rect 6411 20244 6423 20247
rect 6454 20244 6460 20256
rect 6411 20216 6460 20244
rect 6411 20213 6423 20216
rect 6365 20207 6423 20213
rect 6454 20204 6460 20216
rect 6512 20204 6518 20256
rect 6822 20244 6828 20256
rect 6783 20216 6828 20244
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 12713 20247 12771 20253
rect 12713 20213 12725 20247
rect 12759 20244 12771 20247
rect 13078 20244 13084 20256
rect 12759 20216 13084 20244
rect 12759 20213 12771 20216
rect 12713 20207 12771 20213
rect 13078 20204 13084 20216
rect 13136 20204 13142 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 13630 20244 13636 20256
rect 13320 20216 13636 20244
rect 13320 20204 13326 20216
rect 13630 20204 13636 20216
rect 13688 20244 13694 20256
rect 14108 20244 14136 20275
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 15657 20315 15715 20321
rect 15657 20312 15669 20315
rect 14884 20284 15669 20312
rect 14884 20272 14890 20284
rect 15657 20281 15669 20284
rect 15703 20312 15715 20315
rect 16485 20315 16543 20321
rect 16485 20312 16497 20315
rect 15703 20284 16497 20312
rect 15703 20281 15715 20284
rect 15657 20275 15715 20281
rect 16485 20281 16497 20284
rect 16531 20312 16543 20315
rect 18782 20312 18788 20324
rect 16531 20284 18788 20312
rect 16531 20281 16543 20284
rect 16485 20275 16543 20281
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 13688 20216 15301 20244
rect 13688 20204 13694 20216
rect 15289 20213 15301 20216
rect 15335 20244 15347 20247
rect 15470 20244 15476 20256
rect 15335 20216 15476 20244
rect 15335 20213 15347 20216
rect 15289 20207 15347 20213
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2777 20043 2835 20049
rect 2777 20040 2789 20043
rect 1780 20012 2789 20040
rect 1780 19981 1808 20012
rect 2777 20009 2789 20012
rect 2823 20040 2835 20043
rect 2866 20040 2872 20052
rect 2823 20012 2872 20040
rect 2823 20009 2835 20012
rect 2777 20003 2835 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 4212 20012 4445 20040
rect 4212 20000 4218 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 6362 20040 6368 20052
rect 4433 20003 4491 20009
rect 5368 20012 6368 20040
rect 1765 19975 1823 19981
rect 1765 19941 1777 19975
rect 1811 19941 1823 19975
rect 1765 19935 1823 19941
rect 1857 19975 1915 19981
rect 1857 19941 1869 19975
rect 1903 19972 1915 19975
rect 2590 19972 2596 19984
rect 1903 19944 2596 19972
rect 1903 19941 1915 19944
rect 1857 19935 1915 19941
rect 2590 19932 2596 19944
rect 2648 19932 2654 19984
rect 4448 19972 4476 20003
rect 4709 19975 4767 19981
rect 4709 19972 4721 19975
rect 4448 19944 4721 19972
rect 4709 19941 4721 19944
rect 4755 19941 4767 19975
rect 4709 19935 4767 19941
rect 4798 19932 4804 19984
rect 4856 19972 4862 19984
rect 4856 19944 4901 19972
rect 4856 19932 4862 19944
rect 5074 19932 5080 19984
rect 5132 19972 5138 19984
rect 5368 19981 5396 20012
rect 6362 20000 6368 20012
rect 6420 20000 6426 20052
rect 6730 20000 6736 20052
rect 6788 20000 6794 20052
rect 8110 20040 8116 20052
rect 8071 20012 8116 20040
rect 8110 20000 8116 20012
rect 8168 20000 8174 20052
rect 8754 20040 8760 20052
rect 8715 20012 8760 20040
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 9950 20040 9956 20052
rect 9911 20012 9956 20040
rect 9950 20000 9956 20012
rect 10008 20040 10014 20052
rect 10689 20043 10747 20049
rect 10689 20040 10701 20043
rect 10008 20012 10701 20040
rect 10008 20000 10014 20012
rect 10689 20009 10701 20012
rect 10735 20009 10747 20043
rect 11330 20040 11336 20052
rect 11291 20012 11336 20040
rect 10689 20003 10747 20009
rect 11330 20000 11336 20012
rect 11388 20000 11394 20052
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 12805 20043 12863 20049
rect 12805 20040 12817 20043
rect 12768 20012 12817 20040
rect 12768 20000 12774 20012
rect 12805 20009 12817 20012
rect 12851 20009 12863 20043
rect 13906 20040 13912 20052
rect 13867 20012 13912 20040
rect 12805 20003 12863 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 15764 20012 18736 20040
rect 5353 19975 5411 19981
rect 5353 19972 5365 19975
rect 5132 19944 5365 19972
rect 5132 19932 5138 19944
rect 5353 19941 5365 19944
rect 5399 19941 5411 19975
rect 5353 19935 5411 19941
rect 5902 19932 5908 19984
rect 5960 19972 5966 19984
rect 6748 19972 6776 20000
rect 6917 19975 6975 19981
rect 6917 19972 6929 19975
rect 5960 19944 6929 19972
rect 5960 19932 5966 19944
rect 6917 19941 6929 19944
rect 6963 19941 6975 19975
rect 7466 19972 7472 19984
rect 7427 19944 7472 19972
rect 6917 19935 6975 19941
rect 7466 19932 7472 19944
rect 7524 19932 7530 19984
rect 12066 19972 12072 19984
rect 9968 19944 12072 19972
rect 9968 19916 9996 19944
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19904 8355 19907
rect 8386 19904 8392 19916
rect 8343 19876 8392 19904
rect 8343 19873 8355 19876
rect 8297 19867 8355 19873
rect 6270 19796 6276 19848
rect 6328 19836 6334 19848
rect 6822 19836 6828 19848
rect 6328 19808 6828 19836
rect 6328 19796 6334 19808
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 2314 19768 2320 19780
rect 2275 19740 2320 19768
rect 2314 19728 2320 19740
rect 2372 19728 2378 19780
rect 6546 19728 6552 19780
rect 6604 19768 6610 19780
rect 8312 19768 8340 19867
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 9950 19904 9956 19916
rect 9863 19876 9956 19904
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 11532 19913 11560 19944
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 13351 19975 13409 19981
rect 13351 19941 13363 19975
rect 13397 19972 13409 19975
rect 13630 19972 13636 19984
rect 13397 19944 13636 19972
rect 13397 19941 13409 19944
rect 13351 19935 13409 19941
rect 13630 19932 13636 19944
rect 13688 19932 13694 19984
rect 15654 19932 15660 19984
rect 15712 19972 15718 19984
rect 15764 19981 15792 20012
rect 15749 19975 15807 19981
rect 15749 19972 15761 19975
rect 15712 19944 15761 19972
rect 15712 19932 15718 19944
rect 15749 19941 15761 19944
rect 15795 19941 15807 19975
rect 17310 19972 17316 19984
rect 17271 19944 17316 19972
rect 15749 19935 15807 19941
rect 17310 19932 17316 19944
rect 17368 19932 17374 19984
rect 18708 19981 18736 20012
rect 18693 19975 18751 19981
rect 18693 19941 18705 19975
rect 18739 19941 18751 19975
rect 18693 19935 18751 19941
rect 11517 19907 11575 19913
rect 11517 19873 11529 19907
rect 11563 19873 11575 19907
rect 11790 19904 11796 19916
rect 11751 19876 11796 19904
rect 11517 19867 11575 19873
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 18782 19904 18788 19916
rect 18743 19876 18788 19904
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 10152 19836 10180 19864
rect 12986 19836 12992 19848
rect 9539 19808 10180 19836
rect 12947 19808 12992 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 15470 19796 15476 19848
rect 15528 19836 15534 19848
rect 15657 19839 15715 19845
rect 15657 19836 15669 19839
rect 15528 19808 15669 19836
rect 15528 19796 15534 19808
rect 15657 19805 15669 19808
rect 15703 19805 15715 19839
rect 16114 19836 16120 19848
rect 16075 19808 16120 19836
rect 15657 19799 15715 19805
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19805 17279 19839
rect 17221 19799 17279 19805
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19836 17923 19839
rect 18138 19836 18144 19848
rect 17911 19808 18144 19836
rect 17911 19805 17923 19808
rect 17865 19799 17923 19805
rect 14366 19768 14372 19780
rect 6604 19740 8340 19768
rect 14327 19740 14372 19768
rect 6604 19728 6610 19740
rect 14366 19728 14372 19740
rect 14424 19728 14430 19780
rect 17126 19728 17132 19780
rect 17184 19768 17190 19780
rect 17236 19768 17264 19799
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 17184 19740 17264 19768
rect 17184 19728 17190 19740
rect 5721 19703 5779 19709
rect 5721 19669 5733 19703
rect 5767 19700 5779 19703
rect 6362 19700 6368 19712
rect 5767 19672 6368 19700
rect 5767 19669 5779 19672
rect 5721 19663 5779 19669
rect 6362 19660 6368 19672
rect 6420 19660 6426 19712
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8662 19700 8668 19712
rect 8527 19672 8668 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 11146 19700 11152 19712
rect 11059 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19700 11210 19712
rect 12342 19700 12348 19712
rect 11204 19672 12348 19700
rect 11204 19660 11210 19672
rect 12342 19660 12348 19672
rect 12400 19660 12406 19712
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 16574 19700 16580 19712
rect 12492 19672 12537 19700
rect 16535 19672 16580 19700
rect 12492 19660 12498 19672
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 4341 19499 4399 19505
rect 4341 19465 4353 19499
rect 4387 19496 4399 19499
rect 4798 19496 4804 19508
rect 4387 19468 4804 19496
rect 4387 19465 4399 19468
rect 4341 19459 4399 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 6270 19496 6276 19508
rect 6231 19468 6276 19496
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 9769 19499 9827 19505
rect 9769 19465 9781 19499
rect 9815 19496 9827 19499
rect 9950 19496 9956 19508
rect 9815 19468 9956 19496
rect 9815 19465 9827 19468
rect 9769 19459 9827 19465
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 2314 19360 2320 19372
rect 1912 19332 2320 19360
rect 1912 19320 1918 19332
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 8680 19332 9168 19360
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2648 19264 2697 19292
rect 2648 19252 2654 19264
rect 2685 19261 2697 19264
rect 2731 19292 2743 19295
rect 3053 19295 3111 19301
rect 3053 19292 3065 19295
rect 2731 19264 3065 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 3053 19261 3065 19264
rect 3099 19292 3111 19295
rect 3786 19292 3792 19304
rect 3099 19264 3792 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19292 4859 19295
rect 4982 19292 4988 19304
rect 4847 19264 4988 19292
rect 4847 19261 4859 19264
rect 4801 19255 4859 19261
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 6822 19292 6828 19304
rect 6783 19264 6828 19292
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 7742 19292 7748 19304
rect 7703 19264 7748 19292
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 8570 19252 8576 19304
rect 8628 19292 8634 19304
rect 8680 19301 8708 19332
rect 8665 19295 8723 19301
rect 8665 19292 8677 19295
rect 8628 19264 8677 19292
rect 8628 19252 8634 19264
rect 8665 19261 8677 19264
rect 8711 19261 8723 19295
rect 8665 19255 8723 19261
rect 8754 19252 8760 19304
rect 8812 19292 8818 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8812 19264 9045 19292
rect 8812 19252 8818 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9140 19292 9168 19332
rect 9784 19292 9812 19459
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 11885 19499 11943 19505
rect 11885 19465 11897 19499
rect 11931 19496 11943 19499
rect 12066 19496 12072 19508
rect 11931 19468 12072 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 12066 19456 12072 19468
rect 12124 19496 12130 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 12124 19468 12173 19496
rect 12124 19456 12130 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 15654 19496 15660 19508
rect 15615 19468 15660 19496
rect 12161 19459 12219 19465
rect 11146 19360 11152 19372
rect 10980 19332 11152 19360
rect 9140 19264 9812 19292
rect 10597 19295 10655 19301
rect 9033 19255 9091 19261
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 10980 19292 11008 19332
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 12176 19360 12204 19459
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 17310 19456 17316 19508
rect 17368 19496 17374 19508
rect 17405 19499 17463 19505
rect 17405 19496 17417 19499
rect 17368 19468 17417 19496
rect 17368 19456 17374 19468
rect 17405 19465 17417 19468
rect 17451 19465 17463 19499
rect 17405 19459 17463 19465
rect 18782 19456 18788 19508
rect 18840 19496 18846 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 18840 19468 19073 19496
rect 18840 19456 18846 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 14366 19388 14372 19440
rect 14424 19428 14430 19440
rect 14424 19400 14504 19428
rect 14424 19388 14430 19400
rect 14476 19369 14504 19400
rect 15470 19388 15476 19440
rect 15528 19428 15534 19440
rect 15933 19431 15991 19437
rect 15933 19428 15945 19431
rect 15528 19400 15945 19428
rect 15528 19388 15534 19400
rect 15933 19397 15945 19400
rect 15979 19397 15991 19431
rect 15933 19391 15991 19397
rect 14461 19363 14519 19369
rect 12176 19332 12388 19360
rect 10643 19264 11008 19292
rect 11517 19295 11575 19301
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 11517 19261 11529 19295
rect 11563 19292 11575 19295
rect 12158 19292 12164 19304
rect 11563 19264 12164 19292
rect 11563 19261 11575 19264
rect 11517 19255 11575 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12360 19292 12388 19332
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19360 15163 19363
rect 15562 19360 15568 19372
rect 15151 19332 15568 19360
rect 15151 19329 15163 19332
rect 15105 19323 15163 19329
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12360 19264 12449 19292
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12584 19264 12909 19292
rect 12584 19252 12590 19264
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 12986 19252 12992 19304
rect 13044 19292 13050 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 13044 19264 13185 19292
rect 13044 19252 13050 19264
rect 13173 19261 13185 19264
rect 13219 19292 13231 19295
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13219 19264 13829 19292
rect 13219 19261 13231 19264
rect 13173 19255 13231 19261
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 13817 19255 13875 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19261 18199 19295
rect 18141 19255 18199 19261
rect 1670 19224 1676 19236
rect 1583 19196 1676 19224
rect 1670 19184 1676 19196
rect 1728 19184 1734 19236
rect 1762 19184 1768 19236
rect 1820 19224 1826 19236
rect 3145 19227 3203 19233
rect 3145 19224 3157 19227
rect 1820 19196 3157 19224
rect 1820 19184 1826 19196
rect 3145 19193 3157 19196
rect 3191 19193 3203 19227
rect 5163 19227 5221 19233
rect 5163 19224 5175 19227
rect 3145 19187 3203 19193
rect 4724 19196 5175 19224
rect 1688 19156 1716 19184
rect 4724 19168 4752 19196
rect 5163 19193 5175 19196
rect 5209 19224 5221 19227
rect 6549 19227 6607 19233
rect 6549 19224 6561 19227
rect 5209 19196 6561 19224
rect 5209 19193 5221 19196
rect 5163 19187 5221 19193
rect 6549 19193 6561 19196
rect 6595 19224 6607 19227
rect 7187 19227 7245 19233
rect 7187 19224 7199 19227
rect 6595 19196 7199 19224
rect 6595 19193 6607 19196
rect 6549 19187 6607 19193
rect 7187 19193 7199 19196
rect 7233 19224 7245 19227
rect 8110 19224 8116 19236
rect 7233 19196 8116 19224
rect 7233 19193 7245 19196
rect 7187 19187 7245 19193
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 10505 19227 10563 19233
rect 8260 19196 8708 19224
rect 8260 19184 8266 19196
rect 1946 19156 1952 19168
rect 1688 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 4706 19156 4712 19168
rect 4667 19128 4712 19156
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 5721 19159 5779 19165
rect 5721 19156 5733 19159
rect 4856 19128 5733 19156
rect 4856 19116 4862 19128
rect 5721 19125 5733 19128
rect 5767 19125 5779 19159
rect 8386 19156 8392 19168
rect 8347 19128 8392 19156
rect 5721 19119 5779 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 8680 19165 8708 19196
rect 10505 19193 10517 19227
rect 10551 19224 10563 19227
rect 10686 19224 10692 19236
rect 10551 19196 10692 19224
rect 10551 19193 10563 19196
rect 10505 19187 10563 19193
rect 10686 19184 10692 19196
rect 10744 19224 10750 19236
rect 10959 19227 11017 19233
rect 10959 19224 10971 19227
rect 10744 19196 10971 19224
rect 10744 19184 10750 19196
rect 10959 19193 10971 19196
rect 11005 19224 11017 19227
rect 11698 19224 11704 19236
rect 11005 19196 11704 19224
rect 11005 19193 11017 19196
rect 10959 19187 11017 19193
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 14277 19227 14335 19233
rect 14277 19193 14289 19227
rect 14323 19224 14335 19227
rect 14550 19224 14556 19236
rect 14323 19196 14556 19224
rect 14323 19193 14335 19196
rect 14277 19187 14335 19193
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 16485 19227 16543 19233
rect 16485 19193 16497 19227
rect 16531 19193 16543 19227
rect 16485 19187 16543 19193
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19125 8723 19159
rect 10134 19156 10140 19168
rect 10095 19128 10140 19156
rect 8665 19119 8723 19125
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 13541 19159 13599 19165
rect 13541 19125 13553 19159
rect 13587 19156 13599 19159
rect 13630 19156 13636 19168
rect 13587 19128 13636 19156
rect 13587 19125 13599 19128
rect 13541 19119 13599 19125
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 16500 19156 16528 19187
rect 16574 19184 16580 19236
rect 16632 19224 16638 19236
rect 17126 19224 17132 19236
rect 16632 19196 16677 19224
rect 17087 19196 17132 19224
rect 16632 19184 16638 19196
rect 17126 19184 17132 19196
rect 17184 19184 17190 19236
rect 17218 19184 17224 19236
rect 17276 19224 17282 19236
rect 17865 19227 17923 19233
rect 17865 19224 17877 19227
rect 17276 19196 17877 19224
rect 17276 19184 17282 19196
rect 17865 19193 17877 19196
rect 17911 19224 17923 19227
rect 18156 19224 18184 19255
rect 17911 19196 18184 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 16942 19156 16948 19168
rect 16500 19128 16948 19156
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1673 18955 1731 18961
rect 1673 18921 1685 18955
rect 1719 18952 1731 18955
rect 1762 18952 1768 18964
rect 1719 18924 1768 18952
rect 1719 18921 1731 18924
rect 1673 18915 1731 18921
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2004 18924 2973 18952
rect 2004 18912 2010 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 6730 18952 6736 18964
rect 6691 18924 6736 18952
rect 2961 18915 3019 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 6880 18924 7205 18952
rect 6880 18912 6886 18924
rect 7193 18921 7205 18924
rect 7239 18952 7251 18955
rect 7561 18955 7619 18961
rect 7561 18952 7573 18955
rect 7239 18924 7573 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7561 18921 7573 18924
rect 7607 18921 7619 18955
rect 8570 18952 8576 18964
rect 8531 18924 8576 18952
rect 7561 18915 7619 18921
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 9766 18952 9772 18964
rect 9727 18924 9772 18952
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 12250 18952 12256 18964
rect 12211 18924 12256 18952
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 12342 18912 12348 18964
rect 12400 18952 12406 18964
rect 13173 18955 13231 18961
rect 13173 18952 13185 18955
rect 12400 18924 13185 18952
rect 12400 18912 12406 18924
rect 13173 18921 13185 18924
rect 13219 18921 13231 18955
rect 15746 18952 15752 18964
rect 15707 18924 15752 18952
rect 13173 18915 13231 18921
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 16942 18952 16948 18964
rect 16903 18924 16948 18952
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 2133 18887 2191 18893
rect 2133 18853 2145 18887
rect 2179 18884 2191 18887
rect 2682 18884 2688 18896
rect 2179 18856 2688 18884
rect 2179 18853 2191 18856
rect 2133 18847 2191 18853
rect 2682 18844 2688 18856
rect 2740 18844 2746 18896
rect 4614 18884 4620 18896
rect 4575 18856 4620 18884
rect 4614 18844 4620 18856
rect 4672 18844 4678 18896
rect 8588 18884 8616 18912
rect 11698 18893 11704 18896
rect 11695 18884 11704 18893
rect 7760 18856 8616 18884
rect 11659 18856 11704 18884
rect 5994 18816 6000 18828
rect 5955 18788 6000 18816
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 7374 18816 7380 18828
rect 6236 18788 7380 18816
rect 6236 18776 6242 18788
rect 7374 18776 7380 18788
rect 7432 18816 7438 18828
rect 7760 18825 7788 18856
rect 11695 18847 11704 18856
rect 11698 18844 11704 18847
rect 11756 18844 11762 18896
rect 16022 18884 16028 18896
rect 15983 18856 16028 18884
rect 16022 18844 16028 18856
rect 16080 18844 16086 18896
rect 16577 18887 16635 18893
rect 16577 18853 16589 18887
rect 16623 18884 16635 18887
rect 17126 18884 17132 18896
rect 16623 18856 17132 18884
rect 16623 18853 16635 18856
rect 16577 18847 16635 18853
rect 17126 18844 17132 18856
rect 17184 18884 17190 18896
rect 17221 18887 17279 18893
rect 17221 18884 17233 18887
rect 17184 18856 17233 18884
rect 17184 18844 17190 18856
rect 17221 18853 17233 18856
rect 17267 18853 17279 18887
rect 17221 18847 17279 18853
rect 17494 18844 17500 18896
rect 17552 18884 17558 18896
rect 17589 18887 17647 18893
rect 17589 18884 17601 18887
rect 17552 18856 17601 18884
rect 17552 18844 17558 18856
rect 17589 18853 17601 18856
rect 17635 18853 17647 18887
rect 18138 18884 18144 18896
rect 18099 18856 18144 18884
rect 17589 18847 17647 18853
rect 18138 18844 18144 18856
rect 18196 18844 18202 18896
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7432 18788 7757 18816
rect 7432 18776 7438 18788
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 8018 18816 8024 18828
rect 7979 18788 8024 18816
rect 7745 18779 7803 18785
rect 8018 18776 8024 18788
rect 8076 18776 8082 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9953 18819 10011 18825
rect 9953 18816 9965 18819
rect 9548 18788 9965 18816
rect 9548 18776 9554 18788
rect 9953 18785 9965 18788
rect 9999 18816 10011 18819
rect 10042 18816 10048 18828
rect 9999 18788 10048 18816
rect 9999 18785 10011 18788
rect 9953 18779 10011 18785
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 10134 18776 10140 18828
rect 10192 18816 10198 18828
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 10192 18788 10241 18816
rect 10192 18776 10198 18788
rect 10229 18785 10241 18788
rect 10275 18816 10287 18819
rect 10870 18816 10876 18828
rect 10275 18788 10876 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11330 18816 11336 18828
rect 11291 18788 11336 18816
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 13078 18816 13084 18828
rect 12860 18788 13084 18816
rect 12860 18776 12866 18788
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 13170 18776 13176 18828
rect 13228 18816 13234 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 13228 18788 13553 18816
rect 13228 18776 13234 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 1762 18708 1768 18760
rect 1820 18748 1826 18760
rect 2041 18751 2099 18757
rect 2041 18748 2053 18751
rect 1820 18720 2053 18748
rect 1820 18708 1826 18720
rect 2041 18717 2053 18720
rect 2087 18748 2099 18751
rect 3329 18751 3387 18757
rect 3329 18748 3341 18751
rect 2087 18720 3341 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 3329 18717 3341 18720
rect 3375 18717 3387 18751
rect 4522 18748 4528 18760
rect 4483 18720 4528 18748
rect 3329 18711 3387 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15344 18720 15945 18748
rect 15344 18708 15350 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 17862 18748 17868 18760
rect 17543 18720 17868 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17862 18708 17868 18720
rect 17920 18748 17926 18760
rect 18969 18751 19027 18757
rect 18969 18748 18981 18751
rect 17920 18720 18981 18748
rect 17920 18708 17926 18720
rect 18969 18717 18981 18720
rect 19015 18717 19027 18751
rect 18969 18711 19027 18717
rect 2590 18680 2596 18692
rect 2551 18652 2596 18680
rect 2590 18640 2596 18652
rect 2648 18640 2654 18692
rect 5074 18680 5080 18692
rect 5035 18652 5080 18680
rect 5074 18640 5080 18652
rect 5132 18640 5138 18692
rect 9030 18640 9036 18692
rect 9088 18680 9094 18692
rect 9401 18683 9459 18689
rect 9401 18680 9413 18683
rect 9088 18652 9413 18680
rect 9088 18640 9094 18652
rect 9401 18649 9413 18652
rect 9447 18649 9459 18683
rect 9401 18643 9459 18649
rect 5534 18612 5540 18624
rect 5495 18584 5540 18612
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 6178 18612 6184 18624
rect 6139 18584 6184 18612
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18612 9183 18615
rect 9214 18612 9220 18624
rect 9171 18584 9220 18612
rect 9171 18581 9183 18584
rect 9125 18575 9183 18581
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 10781 18615 10839 18621
rect 10781 18581 10793 18615
rect 10827 18612 10839 18615
rect 11054 18612 11060 18624
rect 10827 18584 11060 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11238 18612 11244 18624
rect 11199 18584 11244 18612
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13964 18584 14105 18612
rect 13964 18572 13970 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 4525 18411 4583 18417
rect 4525 18377 4537 18411
rect 4571 18408 4583 18411
rect 4614 18408 4620 18420
rect 4571 18380 4620 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 7374 18408 7380 18420
rect 7335 18380 7380 18408
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 8754 18368 8760 18420
rect 8812 18408 8818 18420
rect 9493 18411 9551 18417
rect 9493 18408 9505 18411
rect 8812 18380 9505 18408
rect 8812 18368 8818 18380
rect 9493 18377 9505 18380
rect 9539 18377 9551 18411
rect 13078 18408 13084 18420
rect 13039 18380 13084 18408
rect 9493 18371 9551 18377
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 14826 18408 14832 18420
rect 14787 18380 14832 18408
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 17862 18408 17868 18420
rect 17823 18380 17868 18408
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 2406 18340 2412 18352
rect 2367 18312 2412 18340
rect 2406 18300 2412 18312
rect 2464 18300 2470 18352
rect 9214 18349 9220 18352
rect 9198 18343 9220 18349
rect 9198 18309 9210 18343
rect 9272 18340 9278 18352
rect 10042 18340 10048 18352
rect 9272 18312 10048 18340
rect 9198 18303 9220 18309
rect 9214 18300 9220 18303
rect 9272 18300 9278 18312
rect 10042 18300 10048 18312
rect 10100 18340 10106 18352
rect 10735 18343 10793 18349
rect 10735 18340 10747 18343
rect 10100 18312 10747 18340
rect 10100 18300 10106 18312
rect 10735 18309 10747 18312
rect 10781 18309 10793 18343
rect 10735 18303 10793 18309
rect 10873 18343 10931 18349
rect 10873 18309 10885 18343
rect 10919 18340 10931 18343
rect 11054 18340 11060 18352
rect 10919 18312 11060 18340
rect 10919 18309 10931 18312
rect 10873 18303 10931 18309
rect 11054 18300 11060 18312
rect 11112 18300 11118 18352
rect 15194 18340 15200 18352
rect 15155 18312 15200 18340
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 15562 18300 15568 18352
rect 15620 18340 15626 18352
rect 16301 18343 16359 18349
rect 16301 18340 16313 18343
rect 15620 18312 16313 18340
rect 15620 18300 15626 18312
rect 16301 18309 16313 18312
rect 16347 18309 16359 18343
rect 16301 18303 16359 18309
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18272 1918 18284
rect 2774 18272 2780 18284
rect 1912 18244 2780 18272
rect 1912 18232 1918 18244
rect 2774 18232 2780 18244
rect 2832 18232 2838 18284
rect 3418 18272 3424 18284
rect 3379 18244 3424 18272
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 3786 18272 3792 18284
rect 3747 18244 3792 18272
rect 3786 18232 3792 18244
rect 3844 18272 3850 18284
rect 4062 18272 4068 18284
rect 3844 18244 4068 18272
rect 3844 18232 3850 18244
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 6687 18244 8064 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 8036 18216 8064 18244
rect 8846 18232 8852 18284
rect 8904 18272 8910 18284
rect 9401 18275 9459 18281
rect 9401 18272 9413 18275
rect 8904 18244 9413 18272
rect 8904 18232 8910 18244
rect 9401 18241 9413 18244
rect 9447 18241 9459 18275
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 9401 18235 9459 18241
rect 10796 18244 10977 18272
rect 5534 18204 5540 18216
rect 5495 18176 5540 18204
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 7742 18204 7748 18216
rect 7703 18176 7748 18204
rect 7742 18164 7748 18176
rect 7800 18164 7806 18216
rect 8018 18204 8024 18216
rect 7931 18176 8024 18204
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9263 18207 9321 18213
rect 9263 18204 9275 18207
rect 9180 18176 9275 18204
rect 9180 18164 9186 18176
rect 9263 18173 9275 18176
rect 9309 18173 9321 18207
rect 9263 18167 9321 18173
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18136 1731 18139
rect 1946 18136 1952 18148
rect 1719 18108 1952 18136
rect 1719 18105 1731 18108
rect 1673 18099 1731 18105
rect 1946 18096 1952 18108
rect 2004 18096 2010 18148
rect 3237 18139 3295 18145
rect 3237 18105 3249 18139
rect 3283 18136 3295 18139
rect 3510 18136 3516 18148
rect 3283 18108 3516 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 3510 18096 3516 18108
rect 3568 18096 3574 18148
rect 4890 18136 4896 18148
rect 4851 18108 4896 18136
rect 4890 18096 4896 18108
rect 4948 18096 4954 18148
rect 6362 18096 6368 18148
rect 6420 18136 6426 18148
rect 8036 18136 8064 18164
rect 8573 18139 8631 18145
rect 8573 18136 8585 18139
rect 6420 18108 7604 18136
rect 8036 18108 8585 18136
rect 6420 18096 6426 18108
rect 2682 18028 2688 18080
rect 2740 18068 2746 18080
rect 2777 18071 2835 18077
rect 2777 18068 2789 18071
rect 2740 18040 2789 18068
rect 2740 18028 2746 18040
rect 2777 18037 2789 18040
rect 2823 18037 2835 18071
rect 2777 18031 2835 18037
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 6089 18071 6147 18077
rect 6089 18068 6101 18071
rect 6052 18040 6101 18068
rect 6052 18028 6058 18040
rect 6089 18037 6101 18040
rect 6135 18068 6147 18071
rect 6914 18068 6920 18080
rect 6135 18040 6920 18068
rect 6135 18037 6147 18040
rect 6089 18031 6147 18037
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 7576 18077 7604 18108
rect 8573 18105 8585 18108
rect 8619 18136 8631 18139
rect 8619 18108 8984 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 7561 18071 7619 18077
rect 7561 18037 7573 18071
rect 7607 18037 7619 18071
rect 8846 18068 8852 18080
rect 8807 18040 8852 18068
rect 7561 18031 7619 18037
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 8956 18068 8984 18108
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 10597 18139 10655 18145
rect 10597 18136 10609 18139
rect 9088 18108 10609 18136
rect 9088 18096 9094 18108
rect 10597 18105 10609 18108
rect 10643 18136 10655 18139
rect 10686 18136 10692 18148
rect 10643 18108 10692 18136
rect 10643 18105 10655 18108
rect 10597 18099 10655 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 9582 18068 9588 18080
rect 8956 18040 9588 18068
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 10192 18040 10425 18068
rect 10192 18028 10198 18040
rect 10413 18037 10425 18040
rect 10459 18068 10471 18071
rect 10796 18068 10824 18244
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 11238 18232 11244 18284
rect 11296 18272 11302 18284
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 11296 18244 11345 18272
rect 11296 18232 11302 18244
rect 11333 18241 11345 18244
rect 11379 18272 11391 18275
rect 11790 18272 11796 18284
rect 11379 18244 11796 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 11790 18232 11796 18244
rect 11848 18272 11854 18284
rect 13170 18272 13176 18284
rect 11848 18244 13176 18272
rect 11848 18232 11854 18244
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 15746 18272 15752 18284
rect 15707 18244 15752 18272
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 16022 18232 16028 18284
rect 16080 18272 16086 18284
rect 16761 18275 16819 18281
rect 16761 18272 16773 18275
rect 16080 18244 16773 18272
rect 16080 18232 16086 18244
rect 16761 18241 16773 18244
rect 16807 18272 16819 18275
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 16807 18244 18061 18272
rect 16807 18241 16819 18244
rect 16761 18235 16819 18241
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18204 12311 18207
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12299 18176 12449 18204
rect 12299 18173 12311 18176
rect 12253 18167 12311 18173
rect 12437 18173 12449 18176
rect 12483 18204 12495 18207
rect 12526 18204 12532 18216
rect 12483 18176 12532 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 13906 18204 13912 18216
rect 13867 18176 13912 18204
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 18138 18204 18144 18216
rect 16632 18176 18144 18204
rect 16632 18164 16638 18176
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 11698 18136 11704 18148
rect 11611 18108 11704 18136
rect 11698 18096 11704 18108
rect 11756 18136 11762 18148
rect 14230 18139 14288 18145
rect 14230 18136 14242 18139
rect 11756 18108 14242 18136
rect 11756 18096 11762 18108
rect 10459 18040 10824 18068
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12621 18071 12679 18077
rect 12621 18068 12633 18071
rect 12492 18040 12633 18068
rect 12492 18028 12498 18040
rect 12621 18037 12633 18040
rect 12667 18037 12679 18071
rect 12621 18031 12679 18037
rect 13630 18028 13636 18080
rect 13688 18068 13694 18080
rect 13740 18077 13768 18108
rect 14230 18105 14242 18108
rect 14276 18105 14288 18139
rect 14230 18099 14288 18105
rect 15102 18096 15108 18148
rect 15160 18136 15166 18148
rect 15565 18139 15623 18145
rect 15565 18136 15577 18139
rect 15160 18108 15577 18136
rect 15160 18096 15166 18108
rect 15565 18105 15577 18108
rect 15611 18136 15623 18139
rect 15841 18139 15899 18145
rect 15841 18136 15853 18139
rect 15611 18108 15853 18136
rect 15611 18105 15623 18108
rect 15565 18099 15623 18105
rect 15841 18105 15853 18108
rect 15887 18136 15899 18139
rect 17218 18136 17224 18148
rect 15887 18108 17224 18136
rect 15887 18105 15899 18108
rect 15841 18099 15899 18105
rect 17218 18096 17224 18108
rect 17276 18096 17282 18148
rect 13725 18071 13783 18077
rect 13725 18068 13737 18071
rect 13688 18040 13737 18068
rect 13688 18028 13694 18040
rect 13725 18037 13737 18040
rect 13771 18037 13783 18071
rect 17494 18068 17500 18080
rect 17455 18040 17500 18068
rect 13725 18031 13783 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2774 17864 2780 17876
rect 2735 17836 2780 17864
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 4522 17864 4528 17876
rect 4483 17836 4528 17864
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 7469 17867 7527 17873
rect 7469 17833 7481 17867
rect 7515 17864 7527 17867
rect 7742 17864 7748 17876
rect 7515 17836 7748 17864
rect 7515 17833 7527 17836
rect 7469 17827 7527 17833
rect 7742 17824 7748 17836
rect 7800 17864 7806 17876
rect 7800 17836 8156 17864
rect 7800 17824 7806 17836
rect 1578 17756 1584 17808
rect 1636 17796 1642 17808
rect 1765 17799 1823 17805
rect 1765 17796 1777 17799
rect 1636 17768 1777 17796
rect 1636 17756 1642 17768
rect 1765 17765 1777 17768
rect 1811 17765 1823 17799
rect 1765 17759 1823 17765
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 2406 17796 2412 17808
rect 1912 17768 1957 17796
rect 2367 17768 2412 17796
rect 1912 17756 1918 17768
rect 2406 17756 2412 17768
rect 2464 17756 2470 17808
rect 4706 17756 4712 17808
rect 4764 17796 4770 17808
rect 4982 17796 4988 17808
rect 4764 17768 4988 17796
rect 4764 17756 4770 17768
rect 4982 17756 4988 17768
rect 5040 17796 5046 17808
rect 7926 17805 7932 17808
rect 5214 17799 5272 17805
rect 5214 17796 5226 17799
rect 5040 17768 5226 17796
rect 5040 17756 5046 17768
rect 5214 17765 5226 17768
rect 5260 17765 5272 17799
rect 5214 17759 5272 17765
rect 7923 17759 7932 17805
rect 7984 17796 7990 17808
rect 8128 17796 8156 17836
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 8352 17836 8493 17864
rect 8352 17824 8358 17836
rect 8481 17833 8493 17836
rect 8527 17833 8539 17867
rect 9490 17864 9496 17876
rect 9451 17836 9496 17864
rect 8481 17827 8539 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10321 17867 10379 17873
rect 10321 17864 10333 17867
rect 9732 17836 10333 17864
rect 9732 17824 9738 17836
rect 10321 17833 10333 17836
rect 10367 17833 10379 17867
rect 10686 17864 10692 17876
rect 10647 17836 10692 17864
rect 10321 17827 10379 17833
rect 10686 17824 10692 17836
rect 10744 17864 10750 17876
rect 11330 17864 11336 17876
rect 10744 17836 11192 17864
rect 11291 17836 11336 17864
rect 10744 17824 10750 17836
rect 9508 17796 9536 17824
rect 7984 17768 8023 17796
rect 8128 17768 9536 17796
rect 11164 17796 11192 17836
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 12158 17864 12164 17876
rect 12119 17836 12164 17864
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12434 17864 12440 17876
rect 12360 17836 12440 17864
rect 11238 17796 11244 17808
rect 11164 17768 11244 17796
rect 7926 17756 7932 17759
rect 7984 17756 7990 17768
rect 11238 17756 11244 17768
rect 11296 17796 11302 17808
rect 12360 17796 12388 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 13170 17864 13176 17876
rect 13131 17836 13176 17864
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 15102 17864 15108 17876
rect 14415 17836 15108 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 16209 17867 16267 17873
rect 16209 17833 16221 17867
rect 16255 17864 16267 17867
rect 16482 17864 16488 17876
rect 16255 17836 16488 17864
rect 16255 17833 16267 17836
rect 16209 17827 16267 17833
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 17494 17864 17500 17876
rect 17455 17836 17500 17864
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 18138 17864 18144 17876
rect 18099 17836 18144 17864
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 11296 17768 12388 17796
rect 11296 17756 11302 17768
rect 13630 17756 13636 17808
rect 13688 17796 13694 17808
rect 15654 17805 15660 17808
rect 13811 17799 13869 17805
rect 13811 17796 13823 17799
rect 13688 17768 13823 17796
rect 13688 17756 13694 17768
rect 13811 17765 13823 17768
rect 13857 17796 13869 17799
rect 15651 17796 15660 17805
rect 13857 17768 15660 17796
rect 13857 17765 13869 17768
rect 13811 17759 13869 17765
rect 15651 17759 15660 17768
rect 15654 17756 15660 17759
rect 15712 17756 15718 17808
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 10686 17728 10692 17740
rect 9723 17700 10692 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 11882 17728 11888 17740
rect 11843 17700 11888 17728
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 13170 17728 13176 17740
rect 12483 17700 13176 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 17310 17728 17316 17740
rect 17271 17700 17316 17728
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18690 17737 18696 17740
rect 18668 17731 18696 17737
rect 18668 17697 18680 17731
rect 18668 17691 18696 17697
rect 18690 17688 18696 17691
rect 18748 17688 18754 17740
rect 4890 17660 4896 17672
rect 4851 17632 4896 17660
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 7558 17660 7564 17672
rect 7519 17632 7564 17660
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10134 17660 10140 17672
rect 10091 17632 10140 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 13320 17632 13461 17660
rect 13320 17620 13326 17632
rect 13449 17629 13461 17632
rect 13495 17660 13507 17663
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 13495 17632 14657 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 15470 17660 15476 17672
rect 15335 17632 15476 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 9784 17592 9812 17620
rect 9953 17595 10011 17601
rect 9953 17592 9965 17595
rect 9784 17564 9965 17592
rect 9953 17561 9965 17564
rect 9999 17561 10011 17595
rect 9953 17555 10011 17561
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5592 17496 5825 17524
rect 5592 17484 5598 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 7098 17524 7104 17536
rect 7059 17496 7104 17524
rect 5813 17487 5871 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 9122 17524 9128 17536
rect 9083 17496 9128 17524
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 9842 17527 9900 17533
rect 9842 17493 9854 17527
rect 9888 17524 9900 17527
rect 10042 17524 10048 17536
rect 9888 17496 10048 17524
rect 9888 17493 9900 17496
rect 9842 17487 9900 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 11793 17527 11851 17533
rect 11793 17524 11805 17527
rect 11204 17496 11805 17524
rect 11204 17484 11210 17496
rect 11793 17493 11805 17496
rect 11839 17524 11851 17527
rect 12894 17524 12900 17536
rect 11839 17496 12900 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 18739 17527 18797 17533
rect 18739 17524 18751 17527
rect 18196 17496 18751 17524
rect 18196 17484 18202 17496
rect 18739 17493 18751 17496
rect 18785 17493 18797 17527
rect 18739 17487 18797 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1765 17323 1823 17329
rect 1765 17289 1777 17323
rect 1811 17320 1823 17323
rect 1854 17320 1860 17332
rect 1811 17292 1860 17320
rect 1811 17289 1823 17292
rect 1765 17283 1823 17289
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 3568 17292 3709 17320
rect 3568 17280 3574 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 3697 17283 3755 17289
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17320 6699 17323
rect 7558 17320 7564 17332
rect 6687 17292 7564 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 8478 17320 8484 17332
rect 8439 17292 8484 17320
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 8849 17323 8907 17329
rect 8849 17289 8861 17323
rect 8895 17320 8907 17323
rect 10042 17320 10048 17332
rect 8895 17292 10048 17320
rect 8895 17289 8907 17292
rect 8849 17283 8907 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10686 17320 10692 17332
rect 10647 17292 10692 17320
rect 10686 17280 10692 17292
rect 10744 17320 10750 17332
rect 10870 17320 10876 17332
rect 10744 17292 10876 17320
rect 10744 17280 10750 17292
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11146 17320 11152 17332
rect 11103 17292 11152 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 12069 17323 12127 17329
rect 12069 17320 12081 17323
rect 11940 17292 12081 17320
rect 11940 17280 11946 17292
rect 12069 17289 12081 17292
rect 12115 17320 12127 17323
rect 12434 17320 12440 17332
rect 12115 17292 12440 17320
rect 12115 17289 12127 17292
rect 12069 17283 12127 17289
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13630 17320 13636 17332
rect 13591 17292 13636 17320
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 16669 17323 16727 17329
rect 16669 17289 16681 17323
rect 16715 17320 16727 17323
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16715 17292 17141 17320
rect 16715 17289 16727 17292
rect 16669 17283 16727 17289
rect 17129 17289 17141 17292
rect 17175 17320 17187 17323
rect 17310 17320 17316 17332
rect 17175 17292 17316 17320
rect 17175 17289 17187 17292
rect 17129 17283 17187 17289
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 18233 17323 18291 17329
rect 18233 17289 18245 17323
rect 18279 17320 18291 17323
rect 19058 17320 19064 17332
rect 18279 17292 19064 17320
rect 18279 17289 18291 17292
rect 18233 17283 18291 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 2961 17255 3019 17261
rect 2961 17221 2973 17255
rect 3007 17252 3019 17255
rect 5905 17255 5963 17261
rect 5905 17252 5917 17255
rect 3007 17224 5917 17252
rect 3007 17221 3019 17224
rect 2961 17215 3019 17221
rect 5905 17221 5917 17224
rect 5951 17221 5963 17255
rect 5905 17215 5963 17221
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17184 2007 17187
rect 2038 17184 2044 17196
rect 1995 17156 2044 17184
rect 1995 17153 2007 17156
rect 1949 17147 2007 17153
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 2590 17184 2596 17196
rect 2551 17156 2596 17184
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 2041 17051 2099 17057
rect 2041 17017 2053 17051
rect 2087 17048 2099 17051
rect 2222 17048 2228 17060
rect 2087 17020 2228 17048
rect 2087 17017 2099 17020
rect 2041 17011 2099 17017
rect 2222 17008 2228 17020
rect 2280 17048 2286 17060
rect 2976 17048 3004 17215
rect 17678 17212 17684 17264
rect 17736 17252 17742 17264
rect 18690 17252 18696 17264
rect 17736 17224 18696 17252
rect 17736 17212 17742 17224
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 6181 17187 6239 17193
rect 6181 17184 6193 17187
rect 4948 17156 6193 17184
rect 4948 17144 4954 17156
rect 6181 17153 6193 17156
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 7098 17144 7104 17196
rect 7156 17184 7162 17196
rect 7558 17184 7564 17196
rect 7156 17156 7564 17184
rect 7156 17144 7162 17156
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 9858 17184 9864 17196
rect 9819 17156 9864 17184
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 13262 17184 13268 17196
rect 13223 17156 13268 17184
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 3326 17116 3332 17128
rect 3239 17088 3332 17116
rect 3326 17076 3332 17088
rect 3384 17116 3390 17128
rect 4062 17116 4068 17128
rect 3384 17088 4068 17116
rect 3384 17076 3390 17088
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4571 17088 4997 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 4985 17085 4997 17088
rect 5031 17116 5043 17119
rect 5534 17116 5540 17128
rect 5031 17088 5540 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 9306 17116 9312 17128
rect 9267 17088 9312 17116
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9456 17088 9781 17116
rect 9456 17076 9462 17088
rect 9769 17085 9781 17088
rect 9815 17085 9827 17119
rect 9769 17079 9827 17085
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10008 17088 10885 17116
rect 10008 17076 10014 17088
rect 10873 17085 10885 17088
rect 10919 17116 10931 17119
rect 11333 17119 11391 17125
rect 11333 17116 11345 17119
rect 10919 17088 11345 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 11333 17085 11345 17088
rect 11379 17085 11391 17119
rect 11333 17079 11391 17085
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17116 12863 17119
rect 12894 17116 12900 17128
rect 12851 17088 12900 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13170 17116 13176 17128
rect 13127 17088 13176 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13170 17076 13176 17088
rect 13228 17076 13234 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13924 17088 14105 17116
rect 7926 17057 7932 17060
rect 5347 17051 5405 17057
rect 5347 17048 5359 17051
rect 2280 17020 3004 17048
rect 5000 17020 5359 17048
rect 2280 17008 2286 17020
rect 5000 16992 5028 17020
rect 5347 17017 5359 17020
rect 5393 17048 5405 17051
rect 7101 17051 7159 17057
rect 7101 17048 7113 17051
rect 5393 17020 7113 17048
rect 5393 17017 5405 17020
rect 5347 17011 5405 17017
rect 7101 17017 7113 17020
rect 7147 17048 7159 17051
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 7147 17020 7481 17048
rect 7147 17017 7159 17020
rect 7101 17011 7159 17017
rect 7469 17017 7481 17020
rect 7515 17048 7527 17051
rect 7923 17048 7932 17057
rect 7515 17020 7932 17048
rect 7515 17017 7527 17020
rect 7469 17011 7527 17017
rect 7923 17011 7932 17020
rect 7926 17008 7932 17011
rect 7984 17008 7990 17060
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 9217 17051 9275 17057
rect 9217 17048 9229 17051
rect 9180 17020 9229 17048
rect 9180 17008 9186 17020
rect 9217 17017 9229 17020
rect 9263 17048 9275 17051
rect 9582 17048 9588 17060
rect 9263 17020 9588 17048
rect 9263 17017 9275 17020
rect 9217 17011 9275 17017
rect 9582 17008 9588 17020
rect 9640 17008 9646 17060
rect 13924 16992 13952 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14642 17116 14648 17128
rect 14603 17088 14648 17116
rect 14093 17079 14151 17085
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 14875 17088 15761 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 15749 17085 15761 17088
rect 15795 17116 15807 17119
rect 15838 17116 15844 17128
rect 15795 17088 15844 17116
rect 15795 17085 15807 17088
rect 15749 17079 15807 17085
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17116 17923 17119
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17911 17088 18061 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 18049 17085 18061 17088
rect 18095 17116 18107 17119
rect 18138 17116 18144 17128
rect 18095 17088 18144 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 15289 17051 15347 17057
rect 15289 17017 15301 17051
rect 15335 17048 15347 17051
rect 16070 17051 16128 17057
rect 16070 17048 16082 17051
rect 15335 17020 16082 17048
rect 15335 17017 15347 17020
rect 15289 17011 15347 17017
rect 15672 16992 15700 17020
rect 16070 17017 16082 17020
rect 16116 17017 16128 17051
rect 16070 17011 16128 17017
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 4982 16980 4988 16992
rect 4939 16952 4988 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10192 16952 10333 16980
rect 10192 16940 10198 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 11790 16980 11796 16992
rect 11751 16952 11796 16980
rect 10321 16943 10379 16949
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 13906 16980 13912 16992
rect 13867 16952 13912 16980
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 15654 16980 15660 16992
rect 15615 16952 15660 16980
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 1673 16779 1731 16785
rect 1673 16776 1685 16779
rect 1636 16748 1685 16776
rect 1636 16736 1642 16748
rect 1673 16745 1685 16748
rect 1719 16745 1731 16779
rect 1673 16739 1731 16745
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2682 16776 2688 16788
rect 2547 16748 2688 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 4948 16748 5273 16776
rect 4948 16736 4954 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 9306 16776 9312 16788
rect 9267 16748 9312 16776
rect 5261 16739 5319 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9858 16776 9864 16788
rect 9819 16748 9864 16776
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12575 16748 12909 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 12897 16739 12955 16745
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 13136 16748 13553 16776
rect 13136 16736 13142 16748
rect 13541 16745 13553 16748
rect 13587 16776 13599 16779
rect 14642 16776 14648 16788
rect 13587 16748 14648 16776
rect 13587 16745 13599 16748
rect 13541 16739 13599 16745
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 15838 16776 15844 16788
rect 15799 16748 15844 16776
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 2096 16680 2360 16708
rect 2096 16668 2102 16680
rect 2222 16640 2228 16652
rect 2183 16612 2228 16640
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 2332 16640 2360 16680
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 3234 16708 3240 16720
rect 2648 16680 3240 16708
rect 2648 16668 2654 16680
rect 3234 16668 3240 16680
rect 3292 16708 3298 16720
rect 3421 16711 3479 16717
rect 3421 16708 3433 16711
rect 3292 16680 3433 16708
rect 3292 16668 3298 16680
rect 3421 16677 3433 16680
rect 3467 16677 3479 16711
rect 3421 16671 3479 16677
rect 4709 16711 4767 16717
rect 4709 16677 4721 16711
rect 4755 16708 4767 16711
rect 4755 16680 6224 16708
rect 4755 16677 4767 16680
rect 4709 16671 4767 16677
rect 3053 16643 3111 16649
rect 3053 16640 3065 16643
rect 2332 16612 3065 16640
rect 3053 16609 3065 16612
rect 3099 16609 3111 16643
rect 4062 16640 4068 16652
rect 4023 16612 4068 16640
rect 3053 16603 3111 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 4985 16643 5043 16649
rect 4985 16640 4997 16643
rect 4948 16612 4997 16640
rect 4948 16600 4954 16612
rect 4985 16609 4997 16612
rect 5031 16609 5043 16643
rect 5350 16640 5356 16652
rect 5311 16612 5356 16640
rect 4985 16603 5043 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 6196 16649 6224 16680
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 11057 16711 11115 16717
rect 6972 16680 7512 16708
rect 6972 16668 6978 16680
rect 7484 16652 7512 16680
rect 11057 16677 11069 16711
rect 11103 16708 11115 16711
rect 11238 16708 11244 16720
rect 11103 16680 11244 16708
rect 11103 16677 11115 16680
rect 11057 16671 11115 16677
rect 11238 16668 11244 16680
rect 11296 16708 11302 16720
rect 11606 16708 11612 16720
rect 11296 16680 11612 16708
rect 11296 16668 11302 16680
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 11793 16711 11851 16717
rect 11793 16677 11805 16711
rect 11839 16708 11851 16711
rect 13096 16708 13124 16736
rect 13814 16708 13820 16720
rect 11839 16680 13124 16708
rect 13775 16680 13820 16708
rect 11839 16677 11851 16680
rect 11793 16671 11851 16677
rect 13814 16668 13820 16680
rect 13872 16668 13878 16720
rect 15470 16708 15476 16720
rect 15431 16680 15476 16708
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 15746 16668 15752 16720
rect 15804 16708 15810 16720
rect 16393 16711 16451 16717
rect 16393 16708 16405 16711
rect 15804 16680 16405 16708
rect 15804 16668 15810 16680
rect 16393 16677 16405 16680
rect 16439 16677 16451 16711
rect 17954 16708 17960 16720
rect 17915 16680 17960 16708
rect 16393 16671 16451 16677
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 5997 16643 6055 16649
rect 5997 16640 6009 16643
rect 5552 16612 6009 16640
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 5552 16572 5580 16612
rect 5997 16609 6009 16612
rect 6043 16640 6055 16643
rect 6181 16643 6239 16649
rect 6043 16612 6132 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 4396 16544 5580 16572
rect 6104 16572 6132 16612
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6362 16640 6368 16652
rect 6227 16612 6368 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6638 16640 6644 16652
rect 6472 16612 6644 16640
rect 6472 16572 6500 16612
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 7742 16640 7748 16652
rect 7524 16612 7748 16640
rect 7524 16600 7530 16612
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8386 16640 8392 16652
rect 7883 16612 8392 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8386 16600 8392 16612
rect 8444 16640 8450 16652
rect 9674 16640 9680 16652
rect 8444 16612 9680 16640
rect 8444 16600 8450 16612
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 12158 16600 12164 16652
rect 12216 16640 12222 16652
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12216 16612 12633 16640
rect 12216 16600 12222 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16640 12955 16643
rect 13170 16640 13176 16652
rect 12943 16612 13176 16640
rect 12943 16609 12955 16612
rect 12897 16603 12955 16609
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13538 16600 13544 16652
rect 13596 16600 13602 16652
rect 19334 16640 19340 16652
rect 15120 16612 16160 16640
rect 19295 16612 19340 16640
rect 6104 16544 6500 16572
rect 4396 16532 4402 16544
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 9766 16572 9772 16584
rect 9640 16544 9772 16572
rect 9640 16532 9646 16544
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16572 11483 16575
rect 11514 16572 11520 16584
rect 11471 16544 11520 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 11514 16532 11520 16544
rect 11572 16572 11578 16584
rect 11790 16572 11796 16584
rect 11572 16544 11796 16572
rect 11572 16532 11578 16544
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 13556 16572 13584 16600
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 13556 16544 13737 16572
rect 13725 16541 13737 16544
rect 13771 16572 13783 16575
rect 14182 16572 14188 16584
rect 13771 16544 14188 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16572 14427 16575
rect 15120 16572 15148 16612
rect 14415 16544 15148 16572
rect 16132 16572 16160 16612
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 16301 16575 16359 16581
rect 16301 16572 16313 16575
rect 16132 16544 16313 16572
rect 14415 16541 14427 16544
rect 14369 16535 14427 16541
rect 16301 16541 16313 16544
rect 16347 16572 16359 16575
rect 16666 16572 16672 16584
rect 16347 16544 16672 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16945 16575 17003 16581
rect 16945 16541 16957 16575
rect 16991 16572 17003 16575
rect 17034 16572 17040 16584
rect 16991 16544 17040 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 17034 16532 17040 16544
rect 17092 16572 17098 16584
rect 17678 16572 17684 16584
rect 17092 16544 17684 16572
rect 17092 16532 17098 16544
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16572 17923 16575
rect 18598 16572 18604 16584
rect 17911 16544 18604 16572
rect 17911 16541 17923 16544
rect 17865 16535 17923 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 7892 16476 8217 16504
rect 7892 16464 7898 16476
rect 8205 16473 8217 16476
rect 8251 16504 8263 16507
rect 8573 16507 8631 16513
rect 8573 16504 8585 16507
rect 8251 16476 8585 16504
rect 8251 16473 8263 16476
rect 8205 16467 8263 16473
rect 8573 16473 8585 16476
rect 8619 16504 8631 16507
rect 9398 16504 9404 16516
rect 8619 16476 9404 16504
rect 8619 16473 8631 16476
rect 8573 16467 8631 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 16684 16504 16712 16532
rect 18417 16507 18475 16513
rect 18417 16504 18429 16507
rect 16684 16476 18429 16504
rect 18417 16473 18429 16476
rect 18463 16473 18475 16507
rect 18417 16467 18475 16473
rect 8754 16396 8760 16448
rect 8812 16436 8818 16448
rect 8849 16439 8907 16445
rect 8849 16436 8861 16439
rect 8812 16408 8861 16436
rect 8812 16396 8818 16408
rect 8849 16405 8861 16408
rect 8895 16405 8907 16439
rect 8849 16399 8907 16405
rect 10042 16396 10048 16448
rect 10100 16436 10106 16448
rect 10502 16436 10508 16448
rect 10100 16408 10508 16436
rect 10100 16396 10106 16408
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10744 16408 10793 16436
rect 10744 16396 10750 16408
rect 10781 16405 10793 16408
rect 10827 16436 10839 16439
rect 10870 16436 10876 16448
rect 10827 16408 10876 16436
rect 10827 16405 10839 16408
rect 10781 16399 10839 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11238 16445 11244 16448
rect 11222 16439 11244 16445
rect 11222 16405 11234 16439
rect 11222 16399 11244 16405
rect 11238 16396 11244 16399
rect 11296 16396 11302 16448
rect 11330 16396 11336 16448
rect 11388 16436 11394 16448
rect 12069 16439 12127 16445
rect 12069 16436 12081 16439
rect 11388 16408 12081 16436
rect 11388 16396 11394 16408
rect 12069 16405 12081 16408
rect 12115 16436 12127 16439
rect 12805 16439 12863 16445
rect 12805 16436 12817 16439
rect 12115 16408 12817 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 12805 16405 12817 16408
rect 12851 16405 12863 16439
rect 19518 16436 19524 16448
rect 19479 16408 19524 16436
rect 12805 16399 12863 16405
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2222 16192 2228 16244
rect 2280 16232 2286 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 2280 16204 2513 16232
rect 2280 16192 2286 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 4338 16232 4344 16244
rect 4299 16204 4344 16232
rect 2501 16195 2559 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 9398 16232 9404 16244
rect 9355 16204 9404 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9732 16204 9873 16232
rect 9732 16192 9738 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 11020 16204 11069 16232
rect 11020 16192 11026 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 11057 16195 11115 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18598 16232 18604 16244
rect 18559 16204 18604 16232
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 19334 16232 19340 16244
rect 19295 16204 19340 16232
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 3786 16164 3792 16176
rect 3747 16136 3792 16164
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 5534 16164 5540 16176
rect 5495 16136 5540 16164
rect 5534 16124 5540 16136
rect 5592 16124 5598 16176
rect 9122 16164 9128 16176
rect 9083 16136 9128 16164
rect 9122 16124 9128 16136
rect 9180 16164 9186 16176
rect 9582 16164 9588 16176
rect 9180 16136 9588 16164
rect 9180 16124 9186 16136
rect 9582 16124 9588 16136
rect 9640 16124 9646 16176
rect 10689 16167 10747 16173
rect 10689 16133 10701 16167
rect 10735 16164 10747 16167
rect 11330 16164 11336 16176
rect 10735 16136 11336 16164
rect 10735 16133 10747 16136
rect 10689 16127 10747 16133
rect 11072 16108 11100 16136
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 17034 16164 17040 16176
rect 16995 16136 17040 16164
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 1946 16096 1952 16108
rect 1627 16068 1952 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 3234 16096 3240 16108
rect 3195 16068 3240 16096
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 5350 16096 5356 16108
rect 5092 16068 5356 16096
rect 5092 16037 5120 16068
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16096 6699 16099
rect 7650 16096 7656 16108
rect 6687 16068 7656 16096
rect 6687 16065 6699 16068
rect 6641 16059 6699 16065
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 16028 4767 16031
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4755 16000 5089 16028
rect 4755 15997 4767 16000
rect 4709 15991 4767 15997
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5626 16028 5632 16040
rect 5587 16000 5632 16028
rect 5077 15991 5135 15997
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 7576 16037 7604 16068
rect 7650 16056 7656 16068
rect 7708 16096 7714 16108
rect 8662 16096 8668 16108
rect 7708 16068 8668 16096
rect 7708 16056 7714 16068
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16096 8815 16099
rect 8846 16096 8852 16108
rect 8803 16068 8852 16096
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 8846 16056 8852 16068
rect 8904 16096 8910 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 8904 16068 9229 16096
rect 8904 16056 8910 16068
rect 9217 16065 9229 16068
rect 9263 16096 9275 16099
rect 10134 16096 10140 16108
rect 9263 16068 10140 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 10134 16056 10140 16068
rect 10192 16096 10198 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 10192 16068 10793 16096
rect 10192 16056 10198 16068
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 7561 16031 7619 16037
rect 5859 16000 6316 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 1673 15963 1731 15969
rect 1673 15929 1685 15963
rect 1719 15960 1731 15963
rect 1762 15960 1768 15972
rect 1719 15932 1768 15960
rect 1719 15929 1731 15932
rect 1673 15923 1731 15929
rect 1762 15920 1768 15932
rect 1820 15920 1826 15972
rect 2225 15963 2283 15969
rect 2225 15929 2237 15963
rect 2271 15960 2283 15963
rect 2682 15960 2688 15972
rect 2271 15932 2688 15960
rect 2271 15929 2283 15932
rect 2225 15923 2283 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15960 3111 15963
rect 3326 15960 3332 15972
rect 3099 15932 3332 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 6288 15901 6316 16000
rect 7561 15997 7573 16031
rect 7607 15997 7619 16031
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7561 15991 7619 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 8996 16031 9054 16037
rect 8996 16028 9008 16031
rect 8435 16000 9008 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 8996 15997 9008 16000
rect 9042 16028 9054 16031
rect 9042 16000 9260 16028
rect 9042 15997 9054 16000
rect 8996 15991 9054 15997
rect 9232 15972 9260 16000
rect 7006 15920 7012 15972
rect 7064 15960 7070 15972
rect 7374 15960 7380 15972
rect 7064 15932 7380 15960
rect 7064 15920 7070 15932
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 8662 15920 8668 15972
rect 8720 15960 8726 15972
rect 8849 15963 8907 15969
rect 8849 15960 8861 15963
rect 8720 15932 8861 15960
rect 8720 15920 8726 15932
rect 8849 15929 8861 15932
rect 8895 15929 8907 15963
rect 8849 15923 8907 15929
rect 9214 15920 9220 15972
rect 9272 15920 9278 15972
rect 6273 15895 6331 15901
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6362 15892 6368 15904
rect 6319 15864 6368 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 7193 15895 7251 15901
rect 7193 15861 7205 15895
rect 7239 15892 7251 15895
rect 7282 15892 7288 15904
rect 7239 15864 7288 15892
rect 7239 15861 7251 15864
rect 7193 15855 7251 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7558 15892 7564 15904
rect 7519 15864 7564 15892
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10244 15901 10272 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 11054 16056 11060 16108
rect 11112 16056 11118 16108
rect 13262 16096 13268 16108
rect 13223 16068 13268 16096
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16485 16099 16543 16105
rect 16485 16096 16497 16099
rect 15979 16068 16497 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16485 16065 16497 16068
rect 16531 16096 16543 16099
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 16531 16068 18061 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 10502 16028 10508 16040
rect 10470 16000 10508 16028
rect 10502 15988 10508 16000
rect 10560 16037 10566 16040
rect 10560 16031 10618 16037
rect 10560 15997 10572 16031
rect 10606 16028 10618 16031
rect 11698 16028 11704 16040
rect 10606 16000 11704 16028
rect 10606 15997 10618 16000
rect 10560 15991 10618 15997
rect 10560 15988 10566 15991
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 16028 12863 16031
rect 12894 16028 12900 16040
rect 12851 16000 12900 16028
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 13078 16028 13084 16040
rect 13039 16000 13084 16028
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13872 16000 14105 16028
rect 13872 15988 13878 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 10413 15963 10471 15969
rect 10413 15929 10425 15963
rect 10459 15960 10471 15963
rect 10686 15960 10692 15972
rect 10459 15932 10692 15960
rect 10459 15929 10471 15932
rect 10413 15923 10471 15929
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 11238 15920 11244 15972
rect 11296 15960 11302 15972
rect 11517 15963 11575 15969
rect 11517 15960 11529 15963
rect 11296 15932 11529 15960
rect 11296 15920 11302 15932
rect 11517 15929 11529 15932
rect 11563 15960 11575 15963
rect 12618 15960 12624 15972
rect 11563 15932 12624 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 12618 15920 12624 15932
rect 12676 15920 12682 15972
rect 14001 15963 14059 15969
rect 14001 15929 14013 15963
rect 14047 15960 14059 15963
rect 14455 15963 14513 15969
rect 14455 15960 14467 15963
rect 14047 15932 14467 15960
rect 14047 15929 14059 15932
rect 14001 15923 14059 15929
rect 14455 15929 14467 15932
rect 14501 15960 14513 15963
rect 15654 15960 15660 15972
rect 14501 15932 15660 15960
rect 14501 15929 14513 15932
rect 14455 15923 14513 15929
rect 15654 15920 15660 15932
rect 15712 15920 15718 15972
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 16574 15960 16580 15972
rect 16347 15932 16580 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 10100 15864 10241 15892
rect 10100 15852 10106 15864
rect 10229 15861 10241 15864
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 11664 15864 11805 15892
rect 11664 15852 11670 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 11793 15855 11851 15861
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 13630 15892 13636 15904
rect 13591 15864 13636 15892
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 15013 15895 15071 15901
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15102 15892 15108 15904
rect 15059 15864 15108 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 15565 15895 15623 15901
rect 15565 15861 15577 15895
rect 15611 15892 15623 15895
rect 15746 15892 15752 15904
rect 15611 15864 15752 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2332 15660 3249 15688
rect 2332 15632 2360 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3237 15651 3295 15657
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4062 15688 4068 15700
rect 3927 15660 4068 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5350 15688 5356 15700
rect 5307 15660 5356 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5534 15688 5540 15700
rect 5495 15660 5540 15688
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7469 15691 7527 15697
rect 7469 15688 7481 15691
rect 6972 15660 7481 15688
rect 6972 15648 6978 15660
rect 7469 15657 7481 15660
rect 7515 15657 7527 15691
rect 7469 15651 7527 15657
rect 10597 15691 10655 15697
rect 10597 15657 10609 15691
rect 10643 15688 10655 15691
rect 10643 15660 13584 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 2314 15620 2320 15632
rect 2275 15592 2320 15620
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 2409 15623 2467 15629
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 2590 15620 2596 15632
rect 2455 15592 2596 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 8018 15620 8024 15632
rect 7668 15592 8024 15620
rect 3970 15512 3976 15564
rect 4028 15552 4034 15564
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 4028 15524 4077 15552
rect 4028 15512 4034 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 6086 15552 6092 15564
rect 5767 15524 6092 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 7668 15561 7696 15592
rect 8018 15580 8024 15592
rect 8076 15580 8082 15632
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 10744 15592 11529 15620
rect 10744 15580 10750 15592
rect 11517 15589 11529 15592
rect 11563 15620 11575 15623
rect 12253 15623 12311 15629
rect 11563 15592 12204 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 6273 15555 6331 15561
rect 6273 15552 6285 15555
rect 6236 15524 6285 15552
rect 6236 15512 6242 15524
rect 6273 15521 6285 15524
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 7837 15555 7895 15561
rect 7837 15521 7849 15555
rect 7883 15521 7895 15555
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 7837 15515 7895 15521
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 5626 15484 5632 15496
rect 5092 15456 5632 15484
rect 5092 15360 5120 15456
rect 5626 15444 5632 15456
rect 5684 15484 5690 15496
rect 6196 15484 6224 15512
rect 6362 15484 6368 15496
rect 5684 15456 6224 15484
rect 6275 15456 6368 15484
rect 5684 15444 5690 15456
rect 6362 15444 6368 15456
rect 6420 15484 6426 15496
rect 6730 15484 6736 15496
rect 6420 15456 6736 15484
rect 6420 15444 6426 15456
rect 6730 15444 6736 15456
rect 6788 15484 6794 15496
rect 7852 15484 7880 15515
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 9950 15552 9956 15564
rect 9911 15524 9956 15552
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 11698 15561 11704 15564
rect 11664 15555 11704 15561
rect 11664 15552 11676 15555
rect 11611 15524 11676 15552
rect 11664 15521 11676 15524
rect 11756 15552 11762 15564
rect 12066 15552 12072 15564
rect 11756 15524 12072 15552
rect 11664 15515 11704 15521
rect 11698 15512 11704 15515
rect 11756 15512 11762 15524
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 6788 15456 8248 15484
rect 6788 15444 6794 15456
rect 8220 15428 8248 15456
rect 10042 15444 10048 15496
rect 10100 15484 10106 15496
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 10100 15456 10333 15484
rect 10100 15444 10106 15456
rect 10321 15453 10333 15456
rect 10367 15453 10379 15487
rect 10321 15447 10379 15453
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11514 15484 11520 15496
rect 11204 15456 11520 15484
rect 11204 15444 11210 15456
rect 11514 15444 11520 15456
rect 11572 15484 11578 15496
rect 11885 15487 11943 15493
rect 11885 15484 11897 15487
rect 11572 15456 11897 15484
rect 11572 15444 11578 15456
rect 11885 15453 11897 15456
rect 11931 15453 11943 15487
rect 12176 15484 12204 15592
rect 12253 15589 12265 15623
rect 12299 15620 12311 15623
rect 12342 15620 12348 15632
rect 12299 15592 12348 15620
rect 12299 15589 12311 15592
rect 12253 15583 12311 15589
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 13081 15555 13139 15561
rect 13081 15552 13093 15555
rect 12492 15524 13093 15552
rect 12492 15512 12498 15524
rect 13081 15521 13093 15524
rect 13127 15521 13139 15555
rect 13081 15515 13139 15521
rect 12710 15484 12716 15496
rect 12176 15456 12716 15484
rect 11885 15447 11943 15453
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 8202 15376 8208 15428
rect 8260 15376 8266 15428
rect 8941 15419 8999 15425
rect 8941 15385 8953 15419
rect 8987 15416 8999 15419
rect 9122 15416 9128 15428
rect 8987 15388 9128 15416
rect 8987 15385 8999 15388
rect 8941 15379 8999 15385
rect 9122 15376 9128 15388
rect 9180 15416 9186 15428
rect 10229 15419 10287 15425
rect 10229 15416 10241 15419
rect 9180 15388 10241 15416
rect 9180 15376 9186 15388
rect 10229 15385 10241 15388
rect 10275 15416 10287 15419
rect 13096 15416 13124 15515
rect 13446 15512 13452 15564
rect 13504 15552 13510 15564
rect 13556 15561 13584 15660
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 14240 15660 14473 15688
rect 14240 15648 14246 15660
rect 14461 15657 14473 15660
rect 14507 15657 14519 15691
rect 14461 15651 14519 15657
rect 15654 15629 15660 15632
rect 15651 15620 15660 15629
rect 15567 15592 15660 15620
rect 15651 15583 15660 15592
rect 15712 15620 15718 15632
rect 16482 15620 16488 15632
rect 15712 15592 16488 15620
rect 15654 15580 15660 15583
rect 15712 15580 15718 15592
rect 16482 15580 16488 15592
rect 16540 15580 16546 15632
rect 16574 15580 16580 15632
rect 16632 15620 16638 15632
rect 17037 15623 17095 15629
rect 17037 15620 17049 15623
rect 16632 15592 17049 15620
rect 16632 15580 16638 15592
rect 17037 15589 17049 15592
rect 17083 15589 17095 15623
rect 17037 15583 17095 15589
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 13504 15524 13553 15552
rect 13504 15512 13510 15524
rect 13541 15521 13553 15524
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 15804 15524 16221 15552
rect 15804 15512 15810 15524
rect 16209 15521 16221 15524
rect 16255 15552 16267 15555
rect 17494 15552 17500 15564
rect 16255 15524 17500 15552
rect 16255 15521 16267 15524
rect 16209 15515 16267 15521
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 13771 15456 15301 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 15289 15453 15301 15456
rect 15335 15484 15347 15487
rect 16114 15484 16120 15496
rect 15335 15456 16120 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 16666 15484 16672 15496
rect 16623 15456 16672 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 13906 15416 13912 15428
rect 10275 15388 11836 15416
rect 13096 15388 13912 15416
rect 10275 15385 10287 15388
rect 10229 15379 10287 15385
rect 11808 15360 11836 15388
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 1673 15351 1731 15357
rect 1673 15317 1685 15351
rect 1719 15348 1731 15351
rect 1762 15348 1768 15360
rect 1719 15320 1768 15348
rect 1719 15317 1731 15320
rect 1673 15311 1731 15317
rect 1762 15308 1768 15320
rect 1820 15308 1826 15360
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 4893 15351 4951 15357
rect 4893 15317 4905 15351
rect 4939 15348 4951 15351
rect 5074 15348 5080 15360
rect 4939 15320 5080 15348
rect 4939 15317 4951 15320
rect 4893 15311 4951 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 7006 15348 7012 15360
rect 6967 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 9214 15308 9220 15360
rect 9272 15348 9278 15360
rect 9401 15351 9459 15357
rect 9401 15348 9413 15351
rect 9272 15320 9413 15348
rect 9272 15308 9278 15320
rect 9401 15317 9413 15320
rect 9447 15348 9459 15351
rect 10091 15351 10149 15357
rect 10091 15348 10103 15351
rect 9447 15320 10103 15348
rect 9447 15317 9459 15320
rect 9401 15311 9459 15317
rect 10091 15317 10103 15320
rect 10137 15317 10149 15351
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 10091 15311 10149 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11790 15348 11796 15360
rect 11751 15320 11796 15348
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 12621 15351 12679 15357
rect 12621 15317 12633 15351
rect 12667 15348 12679 15351
rect 12894 15348 12900 15360
rect 12667 15320 12900 15348
rect 12667 15317 12679 15320
rect 12621 15311 12679 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 13872 15320 14105 15348
rect 13872 15308 13878 15320
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1762 15144 1768 15156
rect 1723 15116 1768 15144
rect 1762 15104 1768 15116
rect 1820 15104 1826 15156
rect 4890 15144 4896 15156
rect 4851 15116 4896 15144
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 4982 15104 4988 15156
rect 5040 15144 5046 15156
rect 5442 15144 5448 15156
rect 5040 15116 5448 15144
rect 5040 15104 5046 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 6144 15116 6193 15144
rect 6144 15104 6150 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6638 15144 6644 15156
rect 6599 15116 6644 15144
rect 6181 15107 6239 15113
rect 2961 15079 3019 15085
rect 2961 15076 2973 15079
rect 2148 15048 2973 15076
rect 2148 14949 2176 15048
rect 2961 15045 2973 15048
rect 3007 15076 3019 15079
rect 3234 15076 3240 15088
rect 3007 15048 3240 15076
rect 3007 15045 3019 15048
rect 2961 15039 3019 15045
rect 3234 15036 3240 15048
rect 3292 15036 3298 15088
rect 6196 15076 6224 15107
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 8018 15144 8024 15156
rect 6748 15116 8024 15144
rect 6748 15076 6776 15116
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 12066 15144 12072 15156
rect 12027 15116 12072 15144
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 13906 15144 13912 15156
rect 13867 15116 13912 15144
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 15378 15144 15384 15156
rect 15339 15116 15384 15144
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 6196 15048 6776 15076
rect 16577 15079 16635 15085
rect 16577 15045 16589 15079
rect 16623 15076 16635 15079
rect 17862 15076 17868 15088
rect 16623 15048 17868 15076
rect 16623 15045 16635 15048
rect 16577 15039 16635 15045
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 2832 14980 3433 15008
rect 2832 14968 2838 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4571 14980 4997 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4985 14977 4997 14980
rect 5031 15008 5043 15011
rect 5442 15008 5448 15020
rect 5031 14980 5448 15008
rect 5031 14977 5043 14980
rect 4985 14971 5043 14977
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 13633 15011 13691 15017
rect 13633 14977 13645 15011
rect 13679 15008 13691 15011
rect 13722 15008 13728 15020
rect 13679 14980 13728 15008
rect 13679 14977 13691 14980
rect 13633 14971 13691 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 16592 15008 16620 15039
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 15344 14980 16620 15008
rect 15344 14968 15350 14980
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14909 2191 14943
rect 2590 14940 2596 14952
rect 2551 14912 2596 14940
rect 2133 14903 2191 14909
rect 2590 14900 2596 14912
rect 2648 14900 2654 14952
rect 5902 14940 5908 14952
rect 5863 14912 5908 14940
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 7006 14940 7012 14952
rect 6967 14912 7012 14940
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8864 14912 9137 14940
rect 2222 14832 2228 14884
rect 2280 14872 2286 14884
rect 2958 14872 2964 14884
rect 2280 14844 2964 14872
rect 2280 14832 2286 14844
rect 2958 14832 2964 14844
rect 3016 14872 3022 14884
rect 3145 14875 3203 14881
rect 3145 14872 3157 14875
rect 3016 14844 3157 14872
rect 3016 14832 3022 14844
rect 3145 14841 3157 14844
rect 3191 14841 3203 14875
rect 3145 14835 3203 14841
rect 3160 14804 3188 14835
rect 3234 14832 3240 14884
rect 3292 14872 3298 14884
rect 3292 14844 3337 14872
rect 3292 14832 3298 14844
rect 4890 14832 4896 14884
rect 4948 14872 4954 14884
rect 5306 14875 5364 14881
rect 5306 14872 5318 14875
rect 4948 14844 5318 14872
rect 4948 14832 4954 14844
rect 5306 14841 5318 14844
rect 5352 14841 5364 14875
rect 5306 14835 5364 14841
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 3160 14776 4077 14804
rect 4065 14773 4077 14776
rect 4111 14773 4123 14807
rect 4065 14767 4123 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7064 14776 7205 14804
rect 7064 14764 7070 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 8864 14813 8892 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10962 14940 10968 14952
rect 10551 14912 10968 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 12894 14940 12900 14952
rect 12855 14912 12900 14940
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13446 14940 13452 14952
rect 13407 14912 13452 14940
rect 13446 14900 13452 14912
rect 13504 14940 13510 14952
rect 15764 14949 15792 14980
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 13504 14912 14289 14940
rect 13504 14900 13510 14912
rect 14277 14909 14289 14912
rect 14323 14940 14335 14943
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14323 14912 14657 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14909 15807 14943
rect 16666 14940 16672 14952
rect 16627 14912 16672 14940
rect 15749 14903 15807 14909
rect 16666 14900 16672 14912
rect 16724 14940 16730 14952
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 16724 14912 17141 14940
rect 16724 14900 16730 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 9769 14875 9827 14881
rect 9769 14841 9781 14875
rect 9815 14872 9827 14875
rect 9950 14872 9956 14884
rect 9815 14844 9956 14872
rect 9815 14841 9827 14844
rect 9769 14835 9827 14841
rect 9950 14832 9956 14844
rect 10008 14832 10014 14884
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10597 14875 10655 14881
rect 10597 14872 10609 14875
rect 10192 14844 10609 14872
rect 10192 14832 10198 14844
rect 10597 14841 10609 14844
rect 10643 14841 10655 14875
rect 10597 14835 10655 14841
rect 8849 14807 8907 14813
rect 8849 14804 8861 14807
rect 8812 14776 8861 14804
rect 8812 14764 8818 14776
rect 8849 14773 8861 14776
rect 8895 14773 8907 14807
rect 10042 14804 10048 14816
rect 10003 14776 10048 14804
rect 8849 14767 8907 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 11701 14807 11759 14813
rect 11701 14773 11713 14807
rect 11747 14804 11759 14807
rect 11790 14804 11796 14816
rect 11747 14776 11796 14804
rect 11747 14773 11759 14776
rect 11701 14767 11759 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12710 14804 12716 14816
rect 12671 14776 12716 14804
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 16209 14807 16267 14813
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 16482 14804 16488 14816
rect 16255 14776 16488 14804
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16850 14804 16856 14816
rect 16811 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 3200 14572 3249 14600
rect 3200 14560 3206 14572
rect 3237 14569 3249 14572
rect 3283 14569 3295 14603
rect 3237 14563 3295 14569
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 3970 14600 3976 14612
rect 3927 14572 3976 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 5169 14603 5227 14609
rect 5169 14569 5181 14603
rect 5215 14600 5227 14603
rect 5258 14600 5264 14612
rect 5215 14572 5264 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 6638 14600 6644 14612
rect 6599 14572 6644 14600
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7742 14600 7748 14612
rect 7703 14572 7748 14600
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 11790 14600 11796 14612
rect 10827 14572 11796 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 12710 14600 12716 14612
rect 12671 14572 12716 14600
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 13228 14572 13461 14600
rect 13228 14560 13234 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13998 14600 14004 14612
rect 13959 14572 14004 14600
rect 13449 14563 13507 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 16114 14600 16120 14612
rect 16075 14572 16120 14600
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 16850 14600 16856 14612
rect 16811 14572 16856 14600
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 6086 14541 6092 14544
rect 6083 14532 6092 14541
rect 6047 14504 6092 14532
rect 6083 14495 6092 14504
rect 6086 14492 6092 14495
rect 6144 14492 6150 14544
rect 9493 14535 9551 14541
rect 9493 14501 9505 14535
rect 9539 14532 9551 14535
rect 9674 14532 9680 14544
rect 9539 14504 9680 14532
rect 9539 14501 9551 14504
rect 9493 14495 9551 14501
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 12728 14532 12756 14560
rect 12805 14535 12863 14541
rect 12805 14532 12817 14535
rect 12728 14504 12817 14532
rect 12805 14501 12817 14504
rect 12851 14501 12863 14535
rect 15838 14532 15844 14544
rect 12805 14495 12863 14501
rect 15212 14504 15844 14532
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14464 2559 14467
rect 2590 14464 2596 14476
rect 2547 14436 2596 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3234 14464 3240 14476
rect 3007 14436 3240 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 4154 14464 4160 14476
rect 4115 14436 4160 14464
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14464 5779 14467
rect 6178 14464 6184 14476
rect 5767 14436 6184 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 6178 14424 6184 14436
rect 6236 14464 6242 14476
rect 6822 14464 6828 14476
rect 6236 14436 6828 14464
rect 6236 14424 6242 14436
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 7650 14464 7656 14476
rect 7611 14436 7656 14464
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 9950 14473 9956 14476
rect 9907 14467 9956 14473
rect 9907 14433 9919 14467
rect 9953 14433 9956 14467
rect 9907 14427 9956 14433
rect 9950 14424 9956 14427
rect 10008 14424 10014 14476
rect 11517 14467 11575 14473
rect 11517 14433 11529 14467
rect 11563 14433 11575 14467
rect 11974 14464 11980 14476
rect 11935 14436 11980 14464
rect 11517 14427 11575 14433
rect 1670 14396 1676 14408
rect 1583 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14396 1734 14408
rect 1857 14399 1915 14405
rect 1857 14396 1869 14399
rect 1728 14368 1869 14396
rect 1728 14356 1734 14368
rect 1857 14365 1869 14368
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 7561 14399 7619 14405
rect 7561 14396 7573 14399
rect 7239 14368 7573 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 7561 14365 7573 14368
rect 7607 14396 7619 14399
rect 8220 14396 8248 14424
rect 7607 14368 8248 14396
rect 7607 14365 7619 14368
rect 7561 14359 7619 14365
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 9824 14368 10057 14396
rect 9824 14356 9830 14368
rect 10045 14365 10057 14368
rect 10091 14396 10103 14399
rect 10134 14396 10140 14408
rect 10091 14368 10140 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 11532 14396 11560 14427
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 12952 14467 13010 14473
rect 12952 14464 12964 14467
rect 12676 14436 12964 14464
rect 12676 14424 12682 14436
rect 12952 14433 12964 14436
rect 12998 14464 13010 14467
rect 15212 14464 15240 14504
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 12998 14436 15240 14464
rect 15289 14467 15347 14473
rect 12998 14433 13010 14436
rect 12952 14427 13010 14433
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15378 14464 15384 14476
rect 15335 14436 15384 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 11882 14396 11888 14408
rect 11532 14368 11888 14396
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 13173 14399 13231 14405
rect 12860 14368 13124 14396
rect 12860 14356 12866 14368
rect 9122 14328 9128 14340
rect 9083 14300 9128 14328
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 10318 14328 10324 14340
rect 9857 14300 10324 14328
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4341 14263 4399 14269
rect 4341 14260 4353 14263
rect 4120 14232 4353 14260
rect 4120 14220 4126 14232
rect 4341 14229 4353 14232
rect 4387 14229 4399 14263
rect 4341 14223 4399 14229
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5537 14263 5595 14269
rect 5537 14260 5549 14263
rect 5132 14232 5549 14260
rect 5132 14220 5138 14232
rect 5537 14229 5549 14232
rect 5583 14229 5595 14263
rect 5537 14223 5595 14229
rect 8757 14263 8815 14269
rect 8757 14229 8769 14263
rect 8803 14260 8815 14263
rect 8938 14260 8944 14272
rect 8803 14232 8944 14260
rect 8803 14229 8815 14232
rect 8757 14223 8815 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9857 14269 9885 14300
rect 10318 14288 10324 14300
rect 10376 14328 10382 14340
rect 11333 14331 11391 14337
rect 11333 14328 11345 14331
rect 10376 14300 11345 14328
rect 10376 14288 10382 14300
rect 11333 14297 11345 14300
rect 11379 14328 11391 14331
rect 12434 14328 12440 14340
rect 11379 14300 12440 14328
rect 11379 14297 11391 14300
rect 11333 14291 11391 14297
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 13096 14337 13124 14368
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 15488 14396 15516 14427
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16669 14467 16727 14473
rect 16669 14464 16681 14467
rect 16632 14436 16681 14464
rect 16632 14424 16638 14436
rect 16669 14433 16681 14436
rect 16715 14433 16727 14467
rect 16669 14427 16727 14433
rect 13173 14359 13231 14365
rect 15396 14368 15516 14396
rect 13081 14331 13139 14337
rect 12544 14300 13032 14328
rect 9824 14263 9885 14269
rect 9824 14229 9836 14263
rect 9870 14232 9885 14263
rect 9870 14229 9882 14232
rect 9824 14223 9882 14229
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10137 14263 10195 14269
rect 10137 14260 10149 14263
rect 10100 14232 10149 14260
rect 10100 14220 10106 14232
rect 10137 14229 10149 14232
rect 10183 14229 10195 14263
rect 11146 14260 11152 14272
rect 11107 14232 11152 14260
rect 10137 14223 10195 14229
rect 11146 14220 11152 14232
rect 11204 14260 11210 14272
rect 12253 14263 12311 14269
rect 12253 14260 12265 14263
rect 11204 14232 12265 14260
rect 11204 14220 11210 14232
rect 12253 14229 12265 14232
rect 12299 14260 12311 14263
rect 12544 14260 12572 14300
rect 12299 14232 12572 14260
rect 13004 14260 13032 14300
rect 13081 14297 13093 14331
rect 13127 14297 13139 14331
rect 13081 14291 13139 14297
rect 13188 14260 13216 14359
rect 15396 14340 15424 14368
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 13004 14232 13216 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2590 14056 2596 14068
rect 2551 14028 2596 14056
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 4154 14056 4160 14068
rect 4067 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14056 4218 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 4212 14028 5733 14056
rect 4212 14016 4218 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 5721 14019 5779 14025
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 7708 14028 8125 14056
rect 7708 14016 7714 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 8113 14019 8171 14025
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9125 14059 9183 14065
rect 9125 14056 9137 14059
rect 8260 14028 9137 14056
rect 8260 14016 8266 14028
rect 9125 14025 9137 14028
rect 9171 14025 9183 14059
rect 9125 14019 9183 14025
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 10962 14056 10968 14068
rect 9539 14028 10968 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11974 14056 11980 14068
rect 11379 14028 11980 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11974 14016 11980 14028
rect 12032 14056 12038 14068
rect 12032 14028 13584 14056
rect 12032 14016 12038 14028
rect 4709 13991 4767 13997
rect 4709 13957 4721 13991
rect 4755 13988 4767 13991
rect 4890 13988 4896 14000
rect 4755 13960 4896 13988
rect 4755 13957 4767 13960
rect 4709 13951 4767 13957
rect 4890 13948 4896 13960
rect 4948 13988 4954 14000
rect 5997 13991 6055 13997
rect 5997 13988 6009 13991
rect 4948 13960 6009 13988
rect 4948 13948 4954 13960
rect 5997 13957 6009 13960
rect 6043 13988 6055 13991
rect 6086 13988 6092 14000
rect 6043 13960 6092 13988
rect 6043 13957 6055 13960
rect 5997 13951 6055 13957
rect 6086 13948 6092 13960
rect 6144 13988 6150 14000
rect 6822 13988 6828 14000
rect 6144 13960 6828 13988
rect 6144 13948 6150 13960
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 8938 13988 8944 14000
rect 8851 13960 8944 13988
rect 8938 13948 8944 13960
rect 8996 13988 9002 14000
rect 8996 13960 9628 13988
rect 8996 13948 9002 13960
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 3142 13920 3148 13932
rect 3103 13892 3148 13920
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3418 13920 3424 13932
rect 3379 13892 3424 13920
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8619 13892 9045 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 9033 13889 9045 13892
rect 9079 13920 9091 13923
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9079 13892 9505 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13821 3019 13855
rect 2961 13815 3019 13821
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13852 4859 13855
rect 6454 13852 6460 13864
rect 4847 13824 6460 13852
rect 4847 13821 4859 13824
rect 4801 13815 4859 13821
rect 1578 13784 1584 13796
rect 1539 13756 1584 13784
rect 1578 13744 1584 13756
rect 1636 13744 1642 13796
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 2976 13784 3004 13815
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13852 7435 13855
rect 7558 13852 7564 13864
rect 7423 13824 7564 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13852 7711 13855
rect 8202 13852 8208 13864
rect 7699 13824 8208 13852
rect 7699 13821 7711 13824
rect 7653 13815 7711 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8812 13855 8870 13861
rect 8812 13821 8824 13855
rect 8858 13852 8870 13855
rect 9122 13852 9128 13864
rect 8858 13824 9128 13852
rect 8858 13821 8870 13824
rect 8812 13815 8870 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 3234 13784 3240 13796
rect 1728 13756 1773 13784
rect 2976 13756 3240 13784
rect 1728 13744 1734 13756
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 4890 13744 4896 13796
rect 4948 13784 4954 13796
rect 5122 13787 5180 13793
rect 5122 13784 5134 13787
rect 4948 13756 5134 13784
rect 4948 13744 4954 13756
rect 5122 13753 5134 13756
rect 5168 13753 5180 13787
rect 8662 13784 8668 13796
rect 8623 13756 8668 13784
rect 5122 13747 5180 13753
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 9600 13784 9628 13960
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10137 13991 10195 13997
rect 10137 13988 10149 13991
rect 10008 13960 10149 13988
rect 10008 13948 10014 13960
rect 10137 13957 10149 13960
rect 10183 13988 10195 13991
rect 11238 13988 11244 14000
rect 10183 13960 11244 13988
rect 10183 13957 10195 13960
rect 10137 13951 10195 13957
rect 11238 13948 11244 13960
rect 11296 13988 11302 14000
rect 12158 13988 12164 14000
rect 11296 13960 12164 13988
rect 11296 13948 11302 13960
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 13078 13988 13084 14000
rect 12299 13960 13084 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13556 13997 13584 14028
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 13872 14028 14289 14056
rect 13872 14016 13878 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 15746 14056 15752 14068
rect 15707 14028 15752 14056
rect 14277 14019 14335 14025
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16632 14028 16681 14056
rect 16632 14016 16638 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 13541 13991 13599 13997
rect 13541 13957 13553 13991
rect 13587 13988 13599 13991
rect 14166 13991 14224 13997
rect 14166 13988 14178 13991
rect 13587 13960 14178 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 14166 13957 14178 13960
rect 14212 13988 14224 13991
rect 14212 13960 15424 13988
rect 14212 13957 14224 13960
rect 14166 13951 14224 13957
rect 15396 13932 15424 13960
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10318 13920 10324 13932
rect 9732 13892 10324 13920
rect 9732 13880 9738 13892
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 13998 13880 14004 13932
rect 14056 13920 14062 13932
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 14056 13892 14381 13920
rect 14056 13880 14062 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 15378 13920 15384 13932
rect 14516 13892 14561 13920
rect 15339 13892 15384 13920
rect 14516 13880 14522 13892
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 16025 13923 16083 13929
rect 16025 13920 16037 13923
rect 15528 13892 16037 13920
rect 15528 13880 15534 13892
rect 16025 13889 16037 13892
rect 16071 13889 16083 13923
rect 16025 13883 16083 13889
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10686 13852 10692 13864
rect 10284 13824 10329 13852
rect 10647 13824 10692 13852
rect 10284 13812 10290 13824
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 13078 13852 13084 13864
rect 11940 13824 12940 13852
rect 13039 13824 13084 13852
rect 11940 13812 11946 13824
rect 11054 13784 11060 13796
rect 9600 13756 11060 13784
rect 9968 13728 9996 13756
rect 11054 13744 11060 13756
rect 11112 13784 11118 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11112 13756 11805 13784
rect 11112 13744 11118 13756
rect 11793 13753 11805 13756
rect 11839 13784 11851 13787
rect 12802 13784 12808 13796
rect 11839 13756 12808 13784
rect 11839 13753 11851 13756
rect 11793 13747 11851 13753
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 12912 13784 12940 13824
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 15562 13852 15568 13864
rect 13280 13824 14044 13852
rect 15523 13824 15568 13852
rect 13173 13787 13231 13793
rect 13173 13784 13185 13787
rect 12912 13756 13185 13784
rect 13173 13753 13185 13756
rect 13219 13784 13231 13787
rect 13280 13784 13308 13824
rect 14016 13796 14044 13824
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 13998 13784 14004 13796
rect 13219 13756 13308 13784
rect 13959 13756 14004 13784
rect 13219 13753 13231 13756
rect 13173 13747 13231 13753
rect 13998 13744 14004 13756
rect 14056 13744 14062 13796
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9677 13719 9735 13725
rect 9677 13716 9689 13719
rect 9640 13688 9689 13716
rect 9640 13676 9646 13688
rect 9677 13685 9689 13688
rect 9723 13685 9735 13719
rect 9677 13679 9735 13685
rect 9950 13676 9956 13728
rect 10008 13676 10014 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 10192 13688 10333 13716
rect 10192 13676 10198 13688
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 13814 13716 13820 13728
rect 13775 13688 13820 13716
rect 10321 13679 10379 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1397 13515 1455 13521
rect 1397 13481 1409 13515
rect 1443 13512 1455 13515
rect 1946 13512 1952 13524
rect 1443 13484 1952 13512
rect 1443 13481 1455 13484
rect 1397 13475 1455 13481
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13512 6147 13515
rect 6178 13512 6184 13524
rect 6135 13484 6184 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7558 13512 7564 13524
rect 7239 13484 7564 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9582 13512 9588 13524
rect 9171 13484 9588 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 11330 13512 11336 13524
rect 11291 13484 11336 13512
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 11480 13484 12173 13512
rect 11480 13472 11486 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12676 13484 12817 13512
rect 12676 13472 12682 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 13170 13512 13176 13524
rect 13131 13484 13176 13512
rect 12805 13475 12863 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 14056 13484 14105 13512
rect 14056 13472 14062 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 2590 13444 2596 13456
rect 2551 13416 2596 13444
rect 2590 13404 2596 13416
rect 2648 13404 2654 13456
rect 4890 13404 4896 13456
rect 4948 13444 4954 13456
rect 5122 13447 5180 13453
rect 5122 13444 5134 13447
rect 4948 13416 5134 13444
rect 4948 13404 4954 13416
rect 5122 13413 5134 13416
rect 5168 13413 5180 13447
rect 5122 13407 5180 13413
rect 7098 13404 7104 13456
rect 7156 13444 7162 13456
rect 7469 13447 7527 13453
rect 7469 13444 7481 13447
rect 7156 13416 7481 13444
rect 7156 13404 7162 13416
rect 7469 13413 7481 13416
rect 7515 13413 7527 13447
rect 7469 13407 7527 13413
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 15562 13444 15568 13456
rect 12492 13416 15568 13444
rect 12492 13404 12498 13416
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 9582 13376 9588 13388
rect 9539 13348 9588 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9692 13348 9965 13376
rect 9692 13320 9720 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10100 13379 10158 13385
rect 10100 13345 10112 13379
rect 10146 13376 10158 13379
rect 10870 13376 10876 13388
rect 10146 13348 10876 13376
rect 10146 13345 10158 13348
rect 10100 13339 10158 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13376 11575 13379
rect 11606 13376 11612 13388
rect 11563 13348 11612 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 13078 13376 13084 13388
rect 13039 13348 13084 13376
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13630 13376 13636 13388
rect 13591 13348 13636 13376
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2866 13308 2872 13320
rect 2547 13280 2872 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2866 13268 2872 13280
rect 2924 13308 2930 13320
rect 3418 13308 3424 13320
rect 2924 13280 3424 13308
rect 2924 13268 2930 13280
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5258 13308 5264 13320
rect 4847 13280 5264 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 7374 13308 7380 13320
rect 7335 13280 7380 13308
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 7616 13280 7665 13308
rect 7616 13268 7622 13280
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 10318 13308 10324 13320
rect 10231 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13308 10382 13320
rect 10962 13308 10968 13320
rect 10376 13280 10968 13308
rect 10376 13268 10382 13280
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11204 13280 11897 13308
rect 11204 13268 11210 13280
rect 11885 13277 11897 13280
rect 11931 13308 11943 13311
rect 11974 13308 11980 13320
rect 11931 13280 11980 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 3050 13240 3056 13252
rect 3011 13212 3056 13240
rect 3050 13200 3056 13212
rect 3108 13200 3114 13252
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 8404 13212 10425 13240
rect 8404 13184 8432 13212
rect 10413 13209 10425 13212
rect 10459 13240 10471 13243
rect 10686 13240 10692 13252
rect 10459 13212 10692 13240
rect 10459 13209 10471 13212
rect 10413 13203 10471 13209
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 12250 13240 12256 13252
rect 10980 13212 12256 13240
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 1949 13175 2007 13181
rect 1949 13172 1961 13175
rect 1636 13144 1961 13172
rect 1636 13132 1642 13144
rect 1949 13141 1961 13144
rect 1995 13172 2007 13175
rect 2498 13172 2504 13184
rect 1995 13144 2504 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10229 13175 10287 13181
rect 10229 13172 10241 13175
rect 10008 13144 10241 13172
rect 10008 13132 10014 13144
rect 10229 13141 10241 13144
rect 10275 13141 10287 13175
rect 10229 13135 10287 13141
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 10980 13181 11008 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 10965 13175 11023 13181
rect 10965 13172 10977 13175
rect 10652 13144 10977 13172
rect 10652 13132 10658 13144
rect 10965 13141 10977 13144
rect 11011 13141 11023 13175
rect 10965 13135 11023 13141
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 11655 13175 11713 13181
rect 11655 13172 11667 13175
rect 11572 13144 11667 13172
rect 11572 13132 11578 13144
rect 11655 13141 11667 13144
rect 11701 13141 11713 13175
rect 11790 13172 11796 13184
rect 11751 13144 11796 13172
rect 11655 13135 11713 13141
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 2648 12940 3341 12968
rect 2648 12928 2654 12940
rect 3329 12937 3341 12940
rect 3375 12968 3387 12971
rect 4154 12968 4160 12980
rect 3375 12940 4160 12968
rect 3375 12937 3387 12940
rect 3329 12931 3387 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4890 12968 4896 12980
rect 4851 12940 4896 12968
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5534 12968 5540 12980
rect 5495 12940 5540 12968
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7009 12971 7067 12977
rect 7009 12968 7021 12971
rect 6972 12940 7021 12968
rect 6972 12928 6978 12940
rect 7009 12937 7021 12940
rect 7055 12937 7067 12971
rect 7009 12931 7067 12937
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7156 12940 8125 12968
rect 7156 12928 7162 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 8113 12931 8171 12937
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8444 12940 8769 12968
rect 8444 12928 8450 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 8757 12931 8815 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 11698 12968 11704 12980
rect 11572 12940 11704 12968
rect 11572 12928 11578 12940
rect 11698 12928 11704 12940
rect 11756 12968 11762 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11756 12940 11897 12968
rect 11756 12928 11762 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 11885 12931 11943 12937
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12575 12971 12633 12977
rect 12575 12968 12587 12971
rect 12492 12940 12587 12968
rect 12492 12928 12498 12940
rect 12575 12937 12587 12940
rect 12621 12937 12633 12971
rect 13078 12968 13084 12980
rect 12991 12940 13084 12968
rect 12575 12931 12633 12937
rect 13078 12928 13084 12940
rect 13136 12968 13142 12980
rect 13630 12968 13636 12980
rect 13136 12940 13636 12968
rect 13136 12928 13142 12940
rect 13630 12928 13636 12940
rect 13688 12968 13694 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 13688 12940 14841 12968
rect 13688 12928 13694 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 14829 12931 14887 12937
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2866 12900 2872 12912
rect 1811 12872 2872 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10318 12900 10324 12912
rect 10091 12872 10324 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 12713 12903 12771 12909
rect 12713 12900 12725 12903
rect 11296 12872 12725 12900
rect 11296 12860 11302 12872
rect 12713 12869 12725 12872
rect 12759 12900 12771 12903
rect 13170 12900 13176 12912
rect 12759 12872 13176 12900
rect 12759 12869 12771 12872
rect 12713 12863 12771 12869
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 13280 12872 13829 12900
rect 3050 12792 3056 12844
rect 3108 12832 3114 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3108 12804 4169 12832
rect 3108 12792 3114 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7190 12832 7196 12844
rect 6687 12804 7196 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 7432 12804 8401 12832
rect 7432 12792 7438 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 12802 12832 12808 12844
rect 12715 12804 12808 12832
rect 8389 12795 8447 12801
rect 12802 12792 12808 12804
rect 12860 12832 12866 12844
rect 13280 12832 13308 12872
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 14185 12903 14243 12909
rect 14185 12869 14197 12903
rect 14231 12869 14243 12903
rect 14185 12863 14243 12869
rect 14200 12832 14228 12863
rect 12860 12804 13308 12832
rect 13832 12804 14228 12832
rect 12860 12792 12866 12804
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 5350 12724 5356 12736
rect 5408 12764 5414 12776
rect 5905 12767 5963 12773
rect 5905 12764 5917 12767
rect 5408 12736 5917 12764
rect 5408 12724 5414 12736
rect 5905 12733 5917 12736
rect 5951 12733 5963 12767
rect 10594 12764 10600 12776
rect 10555 12736 10600 12764
rect 5905 12727 5963 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10744 12736 10885 12764
rect 10744 12724 10750 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 11609 12767 11667 12773
rect 11609 12733 11621 12767
rect 11655 12764 11667 12767
rect 11790 12764 11796 12776
rect 11655 12736 11796 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 11790 12724 11796 12736
rect 11848 12764 11854 12776
rect 13832 12764 13860 12804
rect 11848 12736 13860 12764
rect 11848 12724 11854 12736
rect 13906 12724 13912 12776
rect 13964 12764 13970 12776
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13964 12736 14013 12764
rect 13964 12724 13970 12736
rect 14001 12733 14013 12736
rect 14047 12764 14059 12767
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 14047 12736 14473 12764
rect 14047 12733 14059 12736
rect 14001 12727 14059 12733
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 2314 12696 2320 12708
rect 2275 12668 2320 12696
rect 2314 12656 2320 12668
rect 2372 12656 2378 12708
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 2682 12696 2688 12708
rect 2455 12668 2688 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2424 12628 2452 12659
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 3878 12696 3884 12708
rect 3839 12668 3884 12696
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4062 12696 4068 12708
rect 4019 12668 4068 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 2179 12600 2452 12628
rect 3697 12631 3755 12637
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 3697 12597 3709 12631
rect 3743 12628 3755 12631
rect 3988 12628 4016 12659
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 7514 12699 7572 12705
rect 7514 12696 7526 12699
rect 6972 12668 7526 12696
rect 6972 12656 6978 12668
rect 7514 12665 7526 12668
rect 7560 12696 7572 12699
rect 7926 12696 7932 12708
rect 7560 12668 7932 12696
rect 7560 12665 7572 12668
rect 7514 12659 7572 12665
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8941 12699 8999 12705
rect 8941 12696 8953 12699
rect 8352 12668 8953 12696
rect 8352 12656 8358 12668
rect 8941 12665 8953 12668
rect 8987 12665 8999 12699
rect 8941 12659 8999 12665
rect 12437 12699 12495 12705
rect 12437 12665 12449 12699
rect 12483 12696 12495 12699
rect 12710 12696 12716 12708
rect 12483 12668 12716 12696
rect 12483 12665 12495 12668
rect 12437 12659 12495 12665
rect 12710 12656 12716 12668
rect 12768 12696 12774 12708
rect 13449 12699 13507 12705
rect 13449 12696 13461 12699
rect 12768 12668 13461 12696
rect 12768 12656 12774 12668
rect 13449 12665 13461 12668
rect 13495 12665 13507 12699
rect 13449 12659 13507 12665
rect 5258 12628 5264 12640
rect 3743 12600 4016 12628
rect 5219 12600 5264 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 10686 12628 10692 12640
rect 10647 12600 10692 12628
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3786 12424 3792 12436
rect 2884 12396 3792 12424
rect 1397 12359 1455 12365
rect 1397 12325 1409 12359
rect 1443 12356 1455 12359
rect 2884 12356 2912 12396
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4614 12424 4620 12436
rect 4527 12396 4620 12424
rect 4614 12384 4620 12396
rect 4672 12424 4678 12436
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 4672 12396 4813 12424
rect 4672 12384 4678 12396
rect 4801 12393 4813 12396
rect 4847 12393 4859 12427
rect 4801 12387 4859 12393
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 6788 12396 6837 12424
rect 6788 12384 6794 12396
rect 6825 12393 6837 12396
rect 6871 12393 6883 12427
rect 6825 12387 6883 12393
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 7156 12396 7297 12424
rect 7156 12384 7162 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 7285 12387 7343 12393
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 9180 12396 9413 12424
rect 9180 12384 9186 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9950 12424 9956 12436
rect 9911 12396 9956 12424
rect 9401 12387 9459 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 11606 12424 11612 12436
rect 11567 12396 11612 12424
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11974 12424 11980 12436
rect 11935 12396 11980 12424
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12434 12424 12440 12436
rect 12395 12396 12440 12424
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 13541 12427 13599 12433
rect 13541 12424 13553 12427
rect 12584 12396 13553 12424
rect 12584 12384 12590 12396
rect 13541 12393 13553 12396
rect 13587 12393 13599 12427
rect 13541 12387 13599 12393
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 13909 12427 13967 12433
rect 13909 12424 13921 12427
rect 13872 12396 13921 12424
rect 13872 12384 13878 12396
rect 13909 12393 13921 12396
rect 13955 12393 13967 12427
rect 13909 12387 13967 12393
rect 1443 12328 2912 12356
rect 2976 12328 5304 12356
rect 1443 12325 1455 12328
rect 1397 12319 1455 12325
rect 2498 12288 2504 12300
rect 2459 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 2976 12297 3004 12328
rect 2961 12291 3019 12297
rect 2961 12288 2973 12291
rect 2924 12260 2973 12288
rect 2924 12248 2930 12260
rect 2961 12257 2973 12260
rect 3007 12257 3019 12291
rect 3878 12288 3884 12300
rect 3839 12260 3884 12288
rect 2961 12251 3019 12257
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4338 12288 4344 12300
rect 4212 12260 4344 12288
rect 4212 12248 4218 12260
rect 4338 12248 4344 12260
rect 4396 12288 4402 12300
rect 5276 12297 5304 12328
rect 7926 12316 7932 12368
rect 7984 12365 7990 12368
rect 7984 12359 8032 12365
rect 7984 12325 7986 12359
rect 8020 12325 8032 12359
rect 7984 12319 8032 12325
rect 10775 12359 10833 12365
rect 10775 12325 10787 12359
rect 10821 12356 10833 12359
rect 10962 12356 10968 12368
rect 10821 12328 10968 12356
rect 10821 12325 10833 12328
rect 10775 12319 10833 12325
rect 7984 12316 7990 12319
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 13170 12356 13176 12368
rect 13131 12328 13176 12356
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4396 12260 4721 12288
rect 4396 12248 4402 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 6086 12288 6092 12300
rect 5307 12260 6092 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6270 12248 6276 12300
rect 6328 12288 6334 12300
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6328 12260 6653 12288
rect 6328 12248 6334 12260
rect 6641 12257 6653 12260
rect 6687 12257 6699 12291
rect 12158 12288 12164 12300
rect 12119 12260 12164 12288
rect 6641 12251 6699 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13078 12288 13084 12300
rect 12759 12260 13084 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7432 12192 7665 12220
rect 7432 12180 7438 12192
rect 7653 12189 7665 12192
rect 7699 12220 7711 12223
rect 7742 12220 7748 12232
rect 7699 12192 7748 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10410 12220 10416 12232
rect 10192 12192 10416 12220
rect 10192 12180 10198 12192
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 1486 12044 1492 12096
rect 1544 12084 1550 12096
rect 1857 12087 1915 12093
rect 1857 12084 1869 12087
rect 1544 12056 1869 12084
rect 1544 12044 1550 12056
rect 1857 12053 1869 12056
rect 1903 12053 1915 12087
rect 1857 12047 1915 12053
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 2222 12084 2228 12096
rect 2004 12056 2228 12084
rect 2004 12044 2010 12056
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6730 12084 6736 12096
rect 6595 12056 6736 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 8570 12084 8576 12096
rect 8531 12056 8576 12084
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 8846 12084 8852 12096
rect 8807 12056 8852 12084
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11204 12056 11345 12084
rect 11204 12044 11210 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 11333 12047 11391 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6086 11880 6092 11892
rect 5951 11852 6092 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 7926 11880 7932 11892
rect 7887 11852 7932 11880
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10410 11880 10416 11892
rect 9815 11852 10416 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12860 11852 12909 11880
rect 12860 11840 12866 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 13078 11840 13084 11892
rect 13136 11880 13142 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 13136 11852 13277 11880
rect 13136 11840 13142 11852
rect 13265 11849 13277 11852
rect 13311 11849 13323 11883
rect 13265 11843 13323 11849
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 12621 11815 12679 11821
rect 12621 11812 12633 11815
rect 12032 11784 12633 11812
rect 12032 11772 12038 11784
rect 12621 11781 12633 11784
rect 12667 11781 12679 11815
rect 12621 11775 12679 11781
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2682 11744 2688 11756
rect 2464 11716 2688 11744
rect 2464 11704 2470 11716
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3326 11744 3332 11756
rect 3287 11716 3332 11744
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 4614 11744 4620 11756
rect 4575 11716 4620 11744
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 7558 11744 7564 11756
rect 7519 11716 7564 11744
rect 7558 11704 7564 11716
rect 7616 11744 7622 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7616 11716 8493 11744
rect 7616 11704 7622 11716
rect 8481 11713 8493 11716
rect 8527 11744 8539 11747
rect 8846 11744 8852 11756
rect 8527 11716 8852 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 10686 11676 10692 11688
rect 10643 11648 10692 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 10686 11636 10692 11648
rect 10744 11676 10750 11688
rect 11238 11676 11244 11688
rect 10744 11648 11244 11676
rect 10744 11636 10750 11648
rect 11238 11636 11244 11648
rect 11296 11636 11302 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12802 11676 12808 11688
rect 12483 11648 12808 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 1486 11608 1492 11620
rect 1447 11580 1492 11608
rect 1486 11568 1492 11580
rect 1544 11568 1550 11620
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11577 1639 11611
rect 1581 11571 1639 11577
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2682 11608 2688 11620
rect 2179 11580 2688 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 1596 11540 1624 11571
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 3145 11611 3203 11617
rect 3145 11608 3157 11611
rect 2976 11580 3157 11608
rect 2976 11552 3004 11580
rect 3145 11577 3157 11580
rect 3191 11577 3203 11611
rect 3145 11571 3203 11577
rect 4525 11611 4583 11617
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 4890 11608 4896 11620
rect 4571 11580 4896 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 4890 11568 4896 11580
rect 4948 11617 4954 11620
rect 4948 11611 4996 11617
rect 4948 11577 4950 11611
rect 4984 11577 4996 11611
rect 4948 11571 4996 11577
rect 4948 11568 4954 11571
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 6917 11611 6975 11617
rect 6917 11608 6929 11611
rect 6788 11580 6929 11608
rect 6788 11568 6794 11580
rect 6917 11577 6929 11580
rect 6963 11577 6975 11611
rect 6917 11571 6975 11577
rect 7006 11568 7012 11620
rect 7064 11608 7070 11620
rect 8570 11608 8576 11620
rect 7064 11580 7109 11608
rect 8483 11580 8576 11608
rect 7064 11568 7070 11580
rect 8570 11568 8576 11580
rect 8628 11568 8634 11620
rect 8754 11568 8760 11620
rect 8812 11608 8818 11620
rect 10962 11617 10968 11620
rect 9125 11611 9183 11617
rect 9125 11608 9137 11611
rect 8812 11580 9137 11608
rect 8812 11568 8818 11580
rect 9125 11577 9137 11580
rect 9171 11577 9183 11611
rect 9125 11571 9183 11577
rect 10137 11611 10195 11617
rect 10137 11577 10149 11611
rect 10183 11608 10195 11611
rect 10505 11611 10563 11617
rect 10505 11608 10517 11611
rect 10183 11580 10517 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10505 11577 10517 11580
rect 10551 11608 10563 11611
rect 10959 11608 10968 11617
rect 10551 11580 10968 11608
rect 10551 11577 10563 11580
rect 10505 11571 10563 11577
rect 10959 11571 10968 11580
rect 11020 11608 11026 11620
rect 16482 11608 16488 11620
rect 11020 11580 16488 11608
rect 10962 11568 10968 11571
rect 11020 11568 11026 11580
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 2498 11540 2504 11552
rect 1452 11512 1624 11540
rect 2459 11512 2504 11540
rect 1452 11500 1458 11512
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 2958 11500 2964 11552
rect 3016 11500 3022 11552
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6641 11543 6699 11549
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 7024 11540 7052 11568
rect 6687 11512 7052 11540
rect 8297 11543 8355 11549
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 8297 11509 8309 11543
rect 8343 11540 8355 11543
rect 8588 11540 8616 11568
rect 9490 11540 9496 11552
rect 8343 11512 9496 11540
rect 8343 11509 8355 11512
rect 8297 11503 8355 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 11514 11540 11520 11552
rect 11475 11512 11520 11540
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 3108 11308 3341 11336
rect 3108 11296 3114 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 3329 11299 3387 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6914 11336 6920 11348
rect 6875 11308 6920 11336
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9122 11336 9128 11348
rect 8987 11308 9128 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 2130 11268 2136 11280
rect 2091 11240 2136 11268
rect 2130 11228 2136 11240
rect 2188 11228 2194 11280
rect 4890 11277 4896 11280
rect 4887 11268 4896 11277
rect 4851 11240 4896 11268
rect 4887 11231 4896 11240
rect 4890 11228 4896 11231
rect 4948 11228 4954 11280
rect 7653 11271 7711 11277
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7926 11268 7932 11280
rect 7699 11240 7932 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 8205 11271 8263 11277
rect 8205 11237 8217 11271
rect 8251 11268 8263 11271
rect 8386 11268 8392 11280
rect 8251 11240 8392 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8386 11228 8392 11240
rect 8444 11268 8450 11280
rect 8754 11268 8760 11280
rect 8444 11240 8760 11268
rect 8444 11228 8450 11240
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 10413 11271 10471 11277
rect 10413 11237 10425 11271
rect 10459 11268 10471 11271
rect 11146 11268 11152 11280
rect 10459 11240 11152 11268
rect 10459 11237 10471 11240
rect 10413 11231 10471 11237
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 11977 11271 12035 11277
rect 11977 11268 11989 11271
rect 11940 11240 11989 11268
rect 11940 11228 11946 11240
rect 11977 11237 11989 11240
rect 12023 11237 12035 11271
rect 11977 11231 12035 11237
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 3200 11172 4537 11200
rect 3200 11160 3206 11172
rect 4525 11169 4537 11172
rect 4571 11200 4583 11203
rect 5534 11200 5540 11212
rect 4571 11172 5540 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 6273 11203 6331 11209
rect 6273 11200 6285 11203
rect 6196 11172 6285 11200
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2498 11132 2504 11144
rect 2087 11104 2504 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2682 11132 2688 11144
rect 2643 11104 2688 11132
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 6196 11076 6224 11172
rect 6273 11169 6285 11172
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 7558 11132 7564 11144
rect 7471 11104 7564 11132
rect 7558 11092 7564 11104
rect 7616 11132 7622 11144
rect 8202 11132 8208 11144
rect 7616 11104 8208 11132
rect 7616 11092 7622 11104
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10778 11132 10784 11144
rect 10367 11104 10784 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 11974 11132 11980 11144
rect 11931 11104 11980 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 1581 11067 1639 11073
rect 1581 11064 1593 11067
rect 1452 11036 1593 11064
rect 1452 11024 1458 11036
rect 1581 11033 1593 11036
rect 1627 11033 1639 11067
rect 2958 11064 2964 11076
rect 2919 11036 2964 11064
rect 1581 11027 1639 11033
rect 2958 11024 2964 11036
rect 3016 11064 3022 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 3016 11036 5457 11064
rect 3016 11024 3022 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 6178 11064 6184 11076
rect 6139 11036 6184 11064
rect 5445 11027 5503 11033
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 10873 11067 10931 11073
rect 10873 11033 10885 11067
rect 10919 11033 10931 11067
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 10873 11027 10931 11033
rect 12268 11036 12449 11064
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8481 10999 8539 11005
rect 8481 10996 8493 10999
rect 8352 10968 8493 10996
rect 8352 10956 8358 10968
rect 8481 10965 8493 10968
rect 8527 10996 8539 10999
rect 8662 10996 8668 11008
rect 8527 10968 8668 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 10134 10996 10140 11008
rect 10095 10968 10140 10996
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10888 10996 10916 11027
rect 11054 10996 11060 11008
rect 10888 10968 11060 10996
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12268 10996 12296 11036
rect 12437 11033 12449 11036
rect 12483 11033 12495 11067
rect 12437 11027 12495 11033
rect 12802 10996 12808 11008
rect 11756 10968 12296 10996
rect 12763 10968 12808 10996
rect 11756 10956 11762 10968
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3326 10792 3332 10804
rect 2516 10764 3332 10792
rect 2516 10736 2544 10764
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 3602 10792 3608 10804
rect 3563 10764 3608 10792
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 4890 10792 4896 10804
rect 4571 10764 4896 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 8662 10801 8668 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5592 10764 6009 10792
rect 5592 10752 5598 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 8646 10795 8668 10801
rect 8646 10792 8658 10795
rect 8575 10764 8658 10792
rect 5997 10755 6055 10761
rect 8646 10761 8658 10764
rect 8720 10792 8726 10804
rect 9122 10792 9128 10804
rect 8720 10764 9128 10792
rect 8646 10755 8668 10761
rect 8662 10752 8668 10755
rect 8720 10752 8726 10764
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 2498 10724 2504 10736
rect 2459 10696 2504 10724
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 5074 10684 5080 10736
rect 5132 10684 5138 10736
rect 8389 10727 8447 10733
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 8754 10724 8760 10736
rect 8435 10696 8760 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 9306 10724 9312 10736
rect 8864 10696 9312 10724
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 1780 10628 2881 10656
rect 1302 10480 1308 10532
rect 1360 10520 1366 10532
rect 1780 10520 1808 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 5092 10656 5120 10684
rect 8864 10665 8892 10696
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 4203 10628 5120 10656
rect 5721 10659 5779 10665
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 3418 10588 3424 10600
rect 3379 10560 3424 10588
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 4908 10597 4936 10628
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 8849 10659 8907 10665
rect 5767 10628 8616 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5169 10591 5227 10597
rect 5169 10588 5181 10591
rect 5132 10560 5181 10588
rect 5132 10548 5138 10560
rect 5169 10557 5181 10560
rect 5215 10588 5227 10591
rect 5736 10588 5764 10619
rect 6914 10588 6920 10600
rect 5215 10560 5764 10588
rect 6875 10560 6920 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 1949 10523 2007 10529
rect 1949 10520 1961 10523
rect 1360 10492 1961 10520
rect 1360 10480 1366 10492
rect 1949 10489 1961 10492
rect 1995 10489 2007 10523
rect 1949 10483 2007 10489
rect 2038 10480 2044 10532
rect 2096 10520 2102 10532
rect 7300 10520 7328 10551
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 8352 10560 8493 10588
rect 8352 10548 8358 10560
rect 8481 10557 8493 10560
rect 8527 10557 8539 10591
rect 8588 10588 8616 10628
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 8956 10588 8984 10619
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 11974 10656 11980 10668
rect 10008 10628 11980 10656
rect 10008 10616 10014 10628
rect 11974 10616 11980 10628
rect 12032 10656 12038 10668
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 12032 10628 12173 10656
rect 12032 10616 12038 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 8588 10560 8984 10588
rect 10781 10591 10839 10597
rect 8481 10551 8539 10557
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 11054 10588 11060 10600
rect 10827 10560 11060 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 12802 10588 12808 10600
rect 11204 10560 12808 10588
rect 11204 10548 11210 10560
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 10134 10520 10140 10532
rect 2096 10492 2141 10520
rect 6564 10492 7328 10520
rect 10095 10492 10140 10520
rect 2096 10480 2102 10492
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 2056 10452 2084 10480
rect 6564 10464 6592 10492
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10520 10287 10523
rect 12437 10523 12495 10529
rect 12437 10520 12449 10523
rect 10275 10492 12449 10520
rect 10275 10489 10287 10492
rect 10229 10483 10287 10489
rect 12437 10489 12449 10492
rect 12483 10489 12495 10523
rect 12437 10483 12495 10489
rect 1811 10424 2084 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 4580 10424 4721 10452
rect 4580 10412 4586 10424
rect 4709 10421 4721 10424
rect 4755 10421 4767 10455
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 4709 10415 4767 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 7006 10452 7012 10464
rect 6963 10424 7012 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7926 10452 7932 10464
rect 7887 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 9953 10455 10011 10461
rect 9953 10421 9965 10455
rect 9999 10452 10011 10455
rect 10244 10452 10272 10483
rect 11882 10452 11888 10464
rect 9999 10424 10272 10452
rect 11843 10424 11888 10452
rect 9999 10421 10011 10424
rect 9953 10415 10011 10421
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2130 10248 2136 10260
rect 2087 10220 2136 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 4430 10248 4436 10260
rect 4343 10220 4436 10248
rect 4430 10208 4436 10220
rect 4488 10248 4494 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4488 10220 4629 10248
rect 4488 10208 4494 10220
rect 4617 10217 4629 10220
rect 4663 10217 4675 10251
rect 7558 10248 7564 10260
rect 7519 10220 7564 10248
rect 4617 10211 4675 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 9306 10248 9312 10260
rect 8803 10220 9312 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9950 10248 9956 10260
rect 9911 10220 9956 10248
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10778 10248 10784 10260
rect 10551 10220 10784 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 7837 10183 7895 10189
rect 7837 10149 7849 10183
rect 7883 10180 7895 10183
rect 8202 10180 8208 10192
rect 7883 10152 8208 10180
rect 7883 10149 7895 10152
rect 7837 10143 7895 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 11149 10183 11207 10189
rect 11149 10149 11161 10183
rect 11195 10180 11207 10183
rect 11514 10180 11520 10192
rect 11195 10152 11520 10180
rect 11195 10149 11207 10152
rect 11149 10143 11207 10149
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 11698 10180 11704 10192
rect 11659 10152 11704 10180
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12529 10183 12587 10189
rect 12529 10180 12541 10183
rect 11940 10152 12541 10180
rect 11940 10140 11946 10152
rect 12529 10149 12541 10152
rect 12575 10149 12587 10183
rect 12529 10143 12587 10149
rect 2866 10112 2872 10124
rect 2827 10084 2872 10112
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 4801 10075 4859 10081
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2130 10044 2136 10056
rect 1443 10016 2136 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4154 10044 4160 10056
rect 4028 10016 4160 10044
rect 4028 10004 4034 10016
rect 4154 10004 4160 10016
rect 4212 10044 4218 10056
rect 4816 10044 4844 10075
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 12618 10112 12624 10124
rect 12579 10084 12624 10112
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 6104 10044 6132 10072
rect 4212 10016 6132 10044
rect 6825 10047 6883 10053
rect 4212 10004 4218 10016
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 6914 10044 6920 10056
rect 6871 10016 6920 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7466 10044 7472 10056
rect 7239 10016 7472 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7466 10004 7472 10016
rect 7524 10044 7530 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7524 10016 7757 10044
rect 7524 10004 7530 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8938 10044 8944 10056
rect 8435 10016 8944 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 3513 9911 3571 9917
rect 3513 9908 3525 9911
rect 3476 9880 3525 9908
rect 3476 9868 3482 9880
rect 3513 9877 3525 9880
rect 3559 9908 3571 9911
rect 4062 9908 4068 9920
rect 3559 9880 4068 9908
rect 3559 9877 3571 9880
rect 3513 9871 3571 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 4890 9704 4896 9716
rect 4387 9676 4896 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5629 9707 5687 9713
rect 5629 9704 5641 9707
rect 5132 9676 5641 9704
rect 5132 9664 5138 9676
rect 5629 9673 5641 9676
rect 5675 9673 5687 9707
rect 6086 9704 6092 9716
rect 6047 9676 6092 9704
rect 5629 9667 5687 9673
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 6546 9704 6552 9716
rect 6507 9676 6552 9704
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 8662 9704 8668 9716
rect 8623 9676 8668 9704
rect 8662 9664 8668 9676
rect 8720 9704 8726 9716
rect 9355 9707 9413 9713
rect 9355 9704 9367 9707
rect 8720 9676 9367 9704
rect 8720 9664 8726 9676
rect 9355 9673 9367 9676
rect 9401 9673 9413 9707
rect 9355 9667 9413 9673
rect 9493 9707 9551 9713
rect 9493 9673 9505 9707
rect 9539 9704 9551 9707
rect 9582 9704 9588 9716
rect 9539 9676 9588 9704
rect 9539 9673 9551 9676
rect 9493 9667 9551 9673
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2866 9636 2872 9648
rect 2455 9608 2872 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1443 9472 2084 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 2056 9373 2084 9472
rect 2792 9441 2820 9608
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 3970 9636 3976 9648
rect 3931 9608 3976 9636
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 8812 9608 9137 9636
rect 8812 9596 8818 9608
rect 9125 9605 9137 9608
rect 9171 9636 9183 9639
rect 9508 9636 9536 9667
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11572 9676 11805 9704
rect 11572 9664 11578 9676
rect 11793 9673 11805 9676
rect 11839 9704 11851 9707
rect 12618 9704 12624 9716
rect 11839 9676 12624 9704
rect 11839 9673 11851 9676
rect 11793 9667 11851 9673
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 9674 9636 9680 9648
rect 9171 9608 9536 9636
rect 9635 9608 9680 9636
rect 9171 9605 9183 9608
rect 9125 9599 9183 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 11238 9636 11244 9648
rect 11199 9608 11244 9636
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3050 9568 3056 9580
rect 3007 9540 3056 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3326 9568 3332 9580
rect 3287 9540 3332 9568
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 4430 9568 4436 9580
rect 4391 9540 4436 9568
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 6972 9540 7297 9568
rect 6972 9528 6978 9540
rect 7285 9537 7297 9540
rect 7331 9568 7343 9571
rect 8018 9568 8024 9580
rect 7331 9540 8024 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9364 9540 9597 9568
rect 9364 9528 9370 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 5353 9503 5411 9509
rect 5353 9500 5365 9503
rect 3620 9472 5365 9500
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 3053 9435 3111 9441
rect 3053 9432 3065 9435
rect 2823 9404 3065 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 3053 9401 3065 9404
rect 3099 9432 3111 9435
rect 3620 9432 3648 9472
rect 5353 9469 5365 9472
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 10689 9503 10747 9509
rect 10689 9500 10701 9503
rect 9548 9472 10701 9500
rect 9548 9460 9554 9472
rect 10689 9469 10701 9472
rect 10735 9500 10747 9503
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10735 9472 10885 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 3099 9404 3648 9432
rect 4795 9435 4853 9441
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 4795 9401 4807 9435
rect 4841 9432 4853 9435
rect 4890 9432 4896 9444
rect 4841 9404 4896 9432
rect 4841 9401 4853 9404
rect 4795 9395 4853 9401
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 7606 9435 7664 9441
rect 7606 9432 7618 9435
rect 7116 9404 7618 9432
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2222 9364 2228 9376
rect 2087 9336 2228 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 7116 9373 7144 9404
rect 7606 9401 7618 9404
rect 7652 9401 7664 9435
rect 7606 9395 7664 9401
rect 9122 9392 9128 9444
rect 9180 9432 9186 9444
rect 9217 9435 9275 9441
rect 9217 9432 9229 9435
rect 9180 9404 9229 9432
rect 9180 9392 9186 9404
rect 9217 9401 9229 9404
rect 9263 9432 9275 9435
rect 9398 9432 9404 9444
rect 9263 9404 9404 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 7101 9367 7159 9373
rect 7101 9364 7113 9367
rect 6512 9336 7113 9364
rect 6512 9324 6518 9336
rect 7101 9333 7113 9336
rect 7147 9333 7159 9367
rect 8202 9364 8208 9376
rect 8163 9336 8208 9364
rect 7101 9327 7159 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 4304 9132 4353 9160
rect 4304 9120 4310 9132
rect 4341 9129 4353 9132
rect 4387 9160 4399 9163
rect 5166 9160 5172 9172
rect 4387 9132 5172 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 6052 9132 6285 9160
rect 6052 9120 6058 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 8018 9160 8024 9172
rect 7979 9132 8024 9160
rect 6273 9123 6331 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 2406 9092 2412 9104
rect 2367 9064 2412 9092
rect 2406 9052 2412 9064
rect 2464 9052 2470 9104
rect 2961 9095 3019 9101
rect 2961 9061 2973 9095
rect 3007 9092 3019 9095
rect 3326 9092 3332 9104
rect 3007 9064 3332 9092
rect 3007 9061 3019 9064
rect 2961 9055 3019 9061
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 4795 9095 4853 9101
rect 4795 9061 4807 9095
rect 4841 9092 4853 9095
rect 4890 9092 4896 9104
rect 4841 9064 4896 9092
rect 4841 9061 4853 9064
rect 4795 9055 4853 9061
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 6454 9052 6460 9104
rect 6512 9092 6518 9104
rect 6778 9095 6836 9101
rect 6778 9092 6790 9095
rect 6512 9064 6790 9092
rect 6512 9052 6518 9064
rect 6778 9061 6790 9064
rect 6824 9061 6836 9095
rect 6778 9055 6836 9061
rect 7745 9095 7803 9101
rect 7745 9061 7757 9095
rect 7791 9092 7803 9095
rect 8202 9092 8208 9104
rect 7791 9064 8208 9092
rect 7791 9061 7803 9064
rect 7745 9055 7803 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4522 9024 4528 9036
rect 4479 8996 4528 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 11330 9033 11336 9036
rect 11308 9027 11336 9033
rect 11308 9024 11320 9027
rect 11243 8996 11320 9024
rect 11308 8993 11320 8996
rect 11388 9024 11394 9036
rect 11698 9024 11704 9036
rect 11388 8996 11704 9024
rect 11308 8987 11336 8993
rect 11330 8984 11336 8987
rect 11388 8984 11394 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2188 8928 2329 8956
rect 2188 8916 2194 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6546 8956 6552 8968
rect 6503 8928 6552 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6546 8916 6552 8928
rect 6604 8956 6610 8968
rect 6822 8956 6828 8968
rect 6604 8928 6828 8956
rect 6604 8916 6610 8928
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 8202 8956 8208 8968
rect 8163 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 8812 8928 9689 8956
rect 8812 8916 8818 8928
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 3697 8891 3755 8897
rect 3697 8857 3709 8891
rect 3743 8888 3755 8891
rect 4522 8888 4528 8900
rect 3743 8860 4528 8888
rect 3743 8857 3755 8860
rect 3697 8851 3755 8857
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3016 8792 3249 8820
rect 3016 8780 3022 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 5353 8823 5411 8829
rect 5353 8820 5365 8823
rect 4396 8792 5365 8820
rect 4396 8780 4402 8792
rect 5353 8789 5365 8792
rect 5399 8789 5411 8823
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 5353 8783 5411 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9122 8820 9128 8832
rect 8720 8792 9128 8820
rect 8720 8780 8726 8792
rect 9122 8780 9128 8792
rect 9180 8820 9186 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 9180 8792 9229 8820
rect 9180 8780 9186 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 11379 8823 11437 8829
rect 11379 8820 11391 8823
rect 11112 8792 11391 8820
rect 11112 8780 11118 8792
rect 11379 8789 11391 8792
rect 11425 8789 11437 8823
rect 11379 8783 11437 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2406 8616 2412 8628
rect 2179 8588 2412 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 4430 8616 4436 8628
rect 3743 8588 4436 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 4948 8588 5181 8616
rect 4948 8576 4954 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 3050 8508 3056 8560
rect 3108 8548 3114 8560
rect 3237 8551 3295 8557
rect 3237 8548 3249 8551
rect 3108 8520 3249 8548
rect 3108 8508 3114 8520
rect 3237 8517 3249 8520
rect 3283 8548 3295 8551
rect 5184 8548 5212 8579
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5859 8619 5917 8625
rect 5859 8616 5871 8619
rect 5592 8588 5871 8616
rect 5592 8576 5598 8588
rect 5859 8585 5871 8588
rect 5905 8585 5917 8619
rect 5859 8579 5917 8585
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8202 8616 8208 8628
rect 8159 8588 8208 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9766 8616 9772 8628
rect 9727 8588 9772 8616
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 11330 8616 11336 8628
rect 11291 8588 11336 8616
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 6454 8548 6460 8560
rect 3283 8520 4568 8548
rect 5184 8520 6460 8548
rect 3283 8517 3295 8520
rect 3237 8511 3295 8517
rect 4540 8492 4568 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1578 8480 1584 8492
rect 1360 8452 1584 8480
rect 1360 8440 1366 8452
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2332 8452 2697 8480
rect 2332 8424 2360 8452
rect 2685 8449 2697 8452
rect 2731 8480 2743 8483
rect 2958 8480 2964 8492
rect 2731 8452 2964 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4338 8480 4344 8492
rect 4111 8452 4344 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4522 8480 4528 8492
rect 4483 8452 4528 8480
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6052 8452 7113 8480
rect 6052 8440 6058 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7101 8443 7159 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8220 8480 8248 8576
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8220 8452 8677 8480
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8938 8480 8944 8492
rect 8899 8452 8944 8480
rect 8665 8443 8723 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1670 8412 1676 8424
rect 1443 8384 1676 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 2314 8372 2320 8424
rect 2372 8372 2378 8424
rect 5626 8412 5632 8424
rect 5587 8384 5632 8412
rect 5626 8372 5632 8384
rect 5684 8412 5690 8424
rect 5756 8415 5814 8421
rect 5756 8412 5768 8415
rect 5684 8384 5768 8412
rect 5684 8372 5690 8384
rect 5756 8381 5768 8384
rect 5802 8381 5814 8415
rect 5756 8375 5814 8381
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 2777 8347 2835 8353
rect 2547 8316 2636 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 2608 8276 2636 8316
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 4246 8344 4252 8356
rect 2823 8316 4016 8344
rect 4207 8316 4252 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 2792 8276 2820 8307
rect 2608 8248 2820 8276
rect 3988 8276 4016 8316
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 7193 8347 7251 8353
rect 4396 8316 4441 8344
rect 4396 8304 4402 8316
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 7374 8344 7380 8356
rect 7239 8316 7380 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 8481 8347 8539 8353
rect 8481 8313 8493 8347
rect 8527 8344 8539 8347
rect 8754 8344 8760 8356
rect 8527 8316 8760 8344
rect 8527 8313 8539 8316
rect 8481 8307 8539 8313
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 4154 8276 4160 8288
rect 3988 8248 4160 8276
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1486 8072 1492 8084
rect 1443 8044 1492 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2869 8075 2927 8081
rect 2869 8072 2881 8075
rect 2832 8044 2881 8072
rect 2832 8032 2838 8044
rect 2869 8041 2881 8044
rect 2915 8041 2927 8075
rect 2869 8035 2927 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4212 8044 4353 8072
rect 4212 8032 4218 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 6546 8072 6552 8084
rect 6507 8044 6552 8072
rect 4341 8035 4399 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7432 8044 7665 8072
rect 7432 8032 7438 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 8294 8032 8300 8084
rect 8352 8081 8358 8084
rect 8352 8075 8401 8081
rect 8352 8041 8355 8075
rect 8389 8041 8401 8075
rect 8352 8035 8401 8041
rect 8352 8032 8358 8035
rect 6822 8004 6828 8016
rect 6783 7976 6828 8004
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3510 7936 3516 7948
rect 3099 7908 3516 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 4338 7936 4344 7948
rect 4299 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 7466 7936 7472 7948
rect 7423 7908 7472 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 8272 7939 8330 7945
rect 8272 7905 8284 7939
rect 8318 7936 8330 7939
rect 8386 7936 8392 7948
rect 8318 7908 8392 7936
rect 8318 7905 8330 7908
rect 8272 7899 8330 7905
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6236 7840 6745 7868
rect 6236 7828 6242 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 3237 7531 3295 7537
rect 3237 7497 3249 7531
rect 3283 7528 3295 7531
rect 3510 7528 3516 7540
rect 3283 7500 3516 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 3878 7528 3884 7540
rect 3660 7500 3705 7528
rect 3839 7500 3884 7528
rect 3660 7488 3666 7500
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 4338 7528 4344 7540
rect 4299 7500 4344 7528
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 8386 7528 8392 7540
rect 8343 7500 8392 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 2038 7420 2044 7472
rect 2096 7460 2102 7472
rect 2096 7432 2176 7460
rect 2096 7420 2102 7432
rect 2148 7401 2176 7432
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 4939 7463 4997 7469
rect 4939 7460 4951 7463
rect 4120 7432 4951 7460
rect 4120 7420 4126 7432
rect 4939 7429 4951 7432
rect 4985 7429 4997 7463
rect 4939 7423 4997 7429
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 6822 7392 6828 7404
rect 6687 7364 6828 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 2682 7324 2688 7336
rect 2087 7296 2688 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3660 7296 3709 7324
rect 3660 7284 3666 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 3697 7287 3755 7293
rect 4798 7284 4804 7336
rect 4856 7333 4862 7336
rect 4856 7327 4894 7333
rect 4882 7324 4894 7327
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 4882 7296 5273 7324
rect 4882 7293 4894 7296
rect 4856 7287 4894 7293
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 7374 7324 7380 7336
rect 7335 7296 7380 7324
rect 5261 7287 5319 7293
rect 4856 7284 4862 7287
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 6917 6987 6975 6993
rect 6917 6953 6929 6987
rect 6963 6984 6975 6987
rect 7374 6984 7380 6996
rect 6963 6956 7380 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2038 6848 2044 6860
rect 1951 6820 2044 6848
rect 2038 6808 2044 6820
rect 2096 6848 2102 6860
rect 2406 6848 2412 6860
rect 2096 6820 2412 6848
rect 2096 6808 2102 6820
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 3028 6851 3086 6857
rect 3028 6817 3040 6851
rect 3074 6848 3086 6851
rect 3326 6848 3332 6860
rect 3074 6820 3332 6848
rect 3074 6817 3086 6820
rect 3028 6811 3086 6817
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 3099 6715 3157 6721
rect 3099 6681 3111 6715
rect 3145 6712 3157 6715
rect 4062 6712 4068 6724
rect 3145 6684 4068 6712
rect 3145 6681 3157 6684
rect 3099 6675 3157 6681
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7616 6616 7757 6644
rect 7616 6604 7622 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2590 6400 2596 6452
rect 2648 6449 2654 6452
rect 2648 6443 2697 6449
rect 2648 6409 2651 6443
rect 2685 6409 2697 6443
rect 3326 6440 3332 6452
rect 3287 6412 3332 6440
rect 2648 6403 2697 6409
rect 2648 6400 2654 6403
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 8110 6304 8116 6316
rect 8071 6276 8116 6304
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 1412 6168 1440 6199
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2536 6239 2594 6245
rect 2536 6236 2548 6239
rect 1820 6208 2548 6236
rect 1820 6196 1826 6208
rect 2536 6205 2548 6208
rect 2582 6236 2594 6239
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 2582 6208 2973 6236
rect 2582 6205 2594 6208
rect 2536 6199 2594 6205
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7616 6208 7757 6236
rect 7616 6196 7622 6208
rect 7745 6205 7757 6208
rect 7791 6205 7803 6239
rect 8386 6236 8392 6248
rect 8347 6208 8392 6236
rect 7745 6199 7803 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 2406 6168 2412 6180
rect 1412 6140 2412 6168
rect 2406 6128 2412 6140
rect 2464 6128 2470 6180
rect 7653 6171 7711 6177
rect 7653 6137 7665 6171
rect 7699 6168 7711 6171
rect 8404 6168 8432 6196
rect 7699 6140 8432 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1535 5899 1593 5905
rect 1535 5865 1547 5899
rect 1581 5896 1593 5899
rect 1854 5896 1860 5908
rect 1581 5868 1860 5896
rect 1581 5865 1593 5868
rect 1535 5859 1593 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2590 5905 2596 5908
rect 2547 5899 2596 5905
rect 2547 5865 2559 5899
rect 2593 5865 2596 5899
rect 2547 5859 2596 5865
rect 2590 5856 2596 5859
rect 2648 5856 2654 5908
rect 1486 5769 1492 5772
rect 1464 5763 1492 5769
rect 1464 5729 1476 5763
rect 1464 5723 1492 5729
rect 1486 5720 1492 5723
rect 1544 5720 1550 5772
rect 2498 5769 2504 5772
rect 2476 5763 2504 5769
rect 2476 5729 2488 5763
rect 2476 5723 2504 5729
rect 2498 5720 2504 5723
rect 2556 5720 2562 5772
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7616 5732 7665 5760
rect 7616 5720 7622 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 8018 5556 8024 5568
rect 7979 5528 8024 5556
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1486 5312 1492 5364
rect 1544 5352 1550 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 1544 5324 2237 5352
rect 1544 5312 1550 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2556 5324 2605 5352
rect 2556 5312 2562 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 8018 5352 8024 5364
rect 7979 5324 8024 5352
rect 2593 5315 2651 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 1535 5219 1593 5225
rect 1535 5185 1547 5219
rect 1581 5216 1593 5219
rect 1946 5216 1952 5228
rect 1581 5188 1952 5216
rect 1581 5185 1593 5188
rect 1535 5179 1593 5185
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 8662 5216 8668 5228
rect 8623 5188 8668 5216
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 1394 5108 1400 5160
rect 1452 5157 1458 5160
rect 1452 5151 1490 5157
rect 1478 5148 1490 5151
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1478 5120 1869 5148
rect 1478 5117 1490 5120
rect 1452 5111 1490 5117
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 1452 5108 1458 5111
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 8076 5120 8125 5148
rect 8076 5108 8082 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 8386 5148 8392 5160
rect 8343 5120 8392 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8386 5108 8392 5120
rect 8444 5148 8450 5160
rect 8444 5120 8800 5148
rect 8444 5108 8450 5120
rect 8772 5024 8800 5120
rect 7558 5012 7564 5024
rect 7519 4984 7564 5012
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8812 4984 8953 5012
rect 8812 4972 8818 4984
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 8941 4975 8999 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1578 4817 1584 4820
rect 1535 4811 1584 4817
rect 1535 4777 1547 4811
rect 1581 4777 1584 4811
rect 1535 4771 1584 4777
rect 1578 4768 1584 4771
rect 1636 4768 1642 4820
rect 1394 4632 1400 4684
rect 1452 4681 1458 4684
rect 1452 4675 1490 4681
rect 1478 4641 1490 4675
rect 1452 4635 1490 4641
rect 1452 4632 1458 4635
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1452 4236 1593 4264
rect 1452 4224 1458 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1581 4227 1639 4233
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1535 3723 1593 3729
rect 1535 3689 1547 3723
rect 1581 3720 1593 3723
rect 2314 3720 2320 3732
rect 1581 3692 2320 3720
rect 1581 3689 1593 3692
rect 1535 3683 1593 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 1394 3544 1400 3596
rect 1452 3593 1458 3596
rect 1452 3587 1490 3593
rect 1478 3553 1490 3587
rect 1452 3547 1490 3553
rect 1452 3544 1458 3547
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 19242 3516 19248 3528
rect 18012 3488 19248 3516
rect 18012 3476 18018 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1578 3185 1584 3188
rect 1535 3179 1584 3185
rect 1535 3145 1547 3179
rect 1581 3145 1584 3179
rect 1535 3139 1584 3145
rect 1578 3136 1584 3139
rect 1636 3136 1642 3188
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 2225 3111 2283 3117
rect 2225 3108 2237 3111
rect 1452 3080 2237 3108
rect 1452 3068 1458 3080
rect 2225 3077 2237 3080
rect 2271 3077 2283 3111
rect 2225 3071 2283 3077
rect 1486 2981 1492 2984
rect 1464 2975 1492 2981
rect 1464 2972 1476 2975
rect 1399 2944 1476 2972
rect 1464 2941 1476 2944
rect 1544 2972 1550 2984
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1544 2944 1869 2972
rect 1464 2935 1492 2941
rect 1486 2932 1492 2935
rect 1544 2932 1550 2944
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2641 1584 2644
rect 1535 2635 1584 2641
rect 1535 2601 1547 2635
rect 1581 2601 1584 2635
rect 1535 2595 1584 2601
rect 1578 2592 1584 2595
rect 1636 2592 1642 2644
rect 1394 2456 1400 2508
rect 1452 2505 1458 2508
rect 1452 2499 1490 2505
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1452 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 2476 2499 2534 2505
rect 2476 2465 2488 2499
rect 2522 2496 2534 2499
rect 2866 2496 2872 2508
rect 2522 2468 2872 2496
rect 2522 2465 2534 2468
rect 2476 2459 2534 2465
rect 1452 2456 1458 2459
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 2547 2363 2605 2369
rect 2547 2329 2559 2363
rect 2593 2360 2605 2363
rect 2682 2360 2688 2372
rect 2593 2332 2688 2360
rect 2593 2329 2605 2332
rect 2547 2323 2605 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 4068 26256 4120 26308
rect 6552 26256 6604 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 12900 25440 12952 25492
rect 13912 25483 13964 25492
rect 13912 25449 13921 25483
rect 13921 25449 13955 25483
rect 13955 25449 13964 25483
rect 13912 25440 13964 25449
rect 4068 25304 4120 25356
rect 9220 25304 9272 25356
rect 9772 25347 9824 25356
rect 9772 25313 9816 25347
rect 9816 25313 9824 25347
rect 11612 25347 11664 25356
rect 9772 25304 9824 25313
rect 11612 25313 11621 25347
rect 11621 25313 11655 25347
rect 11655 25313 11664 25347
rect 11612 25304 11664 25313
rect 12624 25347 12676 25356
rect 12624 25313 12633 25347
rect 12633 25313 12667 25347
rect 12667 25313 12676 25347
rect 12624 25304 12676 25313
rect 13820 25304 13872 25356
rect 16304 25304 16356 25356
rect 9680 25100 9732 25152
rect 10692 25100 10744 25152
rect 11428 25143 11480 25152
rect 11428 25109 11437 25143
rect 11437 25109 11471 25143
rect 11471 25109 11480 25143
rect 11428 25100 11480 25109
rect 14280 25143 14332 25152
rect 14280 25109 14289 25143
rect 14289 25109 14323 25143
rect 14323 25109 14332 25143
rect 14280 25100 14332 25109
rect 15752 25100 15804 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 9220 24939 9272 24948
rect 9220 24905 9229 24939
rect 9229 24905 9263 24939
rect 9263 24905 9272 24939
rect 9220 24896 9272 24905
rect 9772 24939 9824 24948
rect 9772 24905 9781 24939
rect 9781 24905 9815 24939
rect 9815 24905 9824 24939
rect 9772 24896 9824 24905
rect 16304 24939 16356 24948
rect 16304 24905 16313 24939
rect 16313 24905 16347 24939
rect 16347 24905 16356 24939
rect 16304 24896 16356 24905
rect 8760 24760 8812 24812
rect 14372 24760 14424 24812
rect 14740 24760 14792 24812
rect 7012 24556 7064 24608
rect 8300 24556 8352 24608
rect 9864 24692 9916 24744
rect 11612 24667 11664 24676
rect 11612 24633 11621 24667
rect 11621 24633 11655 24667
rect 11655 24633 11664 24667
rect 11612 24624 11664 24633
rect 12164 24624 12216 24676
rect 12440 24667 12492 24676
rect 12440 24633 12449 24667
rect 12449 24633 12483 24667
rect 12483 24633 12492 24667
rect 12440 24624 12492 24633
rect 8852 24599 8904 24608
rect 8852 24565 8861 24599
rect 8861 24565 8895 24599
rect 8895 24565 8904 24599
rect 8852 24556 8904 24565
rect 10968 24599 11020 24608
rect 10968 24565 10977 24599
rect 10977 24565 11011 24599
rect 11011 24565 11020 24599
rect 10968 24556 11020 24565
rect 12256 24599 12308 24608
rect 12256 24565 12265 24599
rect 12265 24565 12299 24599
rect 12299 24565 12308 24599
rect 12624 24692 12676 24744
rect 14280 24667 14332 24676
rect 14280 24633 14289 24667
rect 14289 24633 14323 24667
rect 14323 24633 14332 24667
rect 14280 24624 14332 24633
rect 12256 24556 12308 24565
rect 13636 24556 13688 24608
rect 14832 24556 14884 24608
rect 16856 24599 16908 24608
rect 16856 24565 16865 24599
rect 16865 24565 16899 24599
rect 16899 24565 16908 24599
rect 16856 24556 16908 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 14556 24395 14608 24404
rect 14556 24361 14565 24395
rect 14565 24361 14599 24395
rect 14599 24361 14608 24395
rect 14556 24352 14608 24361
rect 15936 24352 15988 24404
rect 11428 24327 11480 24336
rect 11428 24293 11437 24327
rect 11437 24293 11471 24327
rect 11471 24293 11480 24327
rect 11428 24284 11480 24293
rect 12256 24284 12308 24336
rect 4160 24259 4212 24268
rect 4160 24225 4178 24259
rect 4178 24225 4212 24259
rect 4160 24216 4212 24225
rect 5448 24216 5500 24268
rect 6552 24259 6604 24268
rect 6552 24225 6596 24259
rect 6596 24225 6604 24259
rect 8116 24259 8168 24268
rect 6552 24216 6604 24225
rect 8116 24225 8125 24259
rect 8125 24225 8159 24259
rect 8159 24225 8168 24259
rect 8116 24216 8168 24225
rect 9772 24259 9824 24268
rect 9772 24225 9781 24259
rect 9781 24225 9815 24259
rect 9815 24225 9824 24259
rect 9772 24216 9824 24225
rect 15384 24259 15436 24268
rect 15384 24225 15393 24259
rect 15393 24225 15427 24259
rect 15427 24225 15436 24259
rect 15384 24216 15436 24225
rect 16580 24216 16632 24268
rect 18236 24259 18288 24268
rect 18236 24225 18254 24259
rect 18254 24225 18288 24259
rect 18236 24216 18288 24225
rect 25136 24216 25188 24268
rect 11612 24148 11664 24200
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 13176 24191 13228 24200
rect 13176 24157 13185 24191
rect 13185 24157 13219 24191
rect 13219 24157 13228 24191
rect 13176 24148 13228 24157
rect 14648 24148 14700 24200
rect 12348 24080 12400 24132
rect 13820 24123 13872 24132
rect 13820 24089 13829 24123
rect 13829 24089 13863 24123
rect 13863 24089 13872 24123
rect 13820 24080 13872 24089
rect 17960 24080 18012 24132
rect 4896 24012 4948 24064
rect 6828 24012 6880 24064
rect 8024 24055 8076 24064
rect 8024 24021 8033 24055
rect 8033 24021 8067 24055
rect 8067 24021 8076 24055
rect 8024 24012 8076 24021
rect 8852 24055 8904 24064
rect 8852 24021 8861 24055
rect 8861 24021 8895 24055
rect 8895 24021 8904 24055
rect 8852 24012 8904 24021
rect 9956 24055 10008 24064
rect 9956 24021 9965 24055
rect 9965 24021 9999 24055
rect 9999 24021 10008 24055
rect 9956 24012 10008 24021
rect 12532 24055 12584 24064
rect 12532 24021 12541 24055
rect 12541 24021 12575 24055
rect 12575 24021 12584 24055
rect 12532 24012 12584 24021
rect 23572 24012 23624 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1400 23647 1452 23656
rect 1400 23613 1444 23647
rect 1444 23613 1452 23647
rect 1400 23604 1452 23613
rect 4620 23808 4672 23860
rect 5264 23851 5316 23860
rect 5264 23817 5273 23851
rect 5273 23817 5307 23851
rect 5307 23817 5316 23851
rect 5264 23808 5316 23817
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 7748 23808 7800 23860
rect 9772 23808 9824 23860
rect 11060 23808 11112 23860
rect 11428 23808 11480 23860
rect 13820 23808 13872 23860
rect 4160 23783 4212 23792
rect 4160 23749 4169 23783
rect 4169 23749 4203 23783
rect 4203 23749 4212 23783
rect 4160 23740 4212 23749
rect 8852 23740 8904 23792
rect 9128 23715 9180 23724
rect 9128 23681 9137 23715
rect 9137 23681 9171 23715
rect 9171 23681 9180 23715
rect 9128 23672 9180 23681
rect 12164 23672 12216 23724
rect 12624 23672 12676 23724
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 14556 23672 14608 23681
rect 14832 23715 14884 23724
rect 14832 23681 14841 23715
rect 14841 23681 14875 23715
rect 14875 23681 14884 23715
rect 14832 23672 14884 23681
rect 8116 23647 8168 23656
rect 2688 23536 2740 23588
rect 5264 23536 5316 23588
rect 8116 23613 8125 23647
rect 8125 23613 8159 23647
rect 8159 23613 8168 23647
rect 8116 23604 8168 23613
rect 8484 23604 8536 23656
rect 11612 23647 11664 23656
rect 11612 23613 11621 23647
rect 11621 23613 11655 23647
rect 11655 23613 11664 23647
rect 11612 23604 11664 23613
rect 18236 23808 18288 23860
rect 18972 23851 19024 23860
rect 18972 23817 18981 23851
rect 18981 23817 19015 23851
rect 19015 23817 19024 23851
rect 18972 23808 19024 23817
rect 18972 23604 19024 23656
rect 21180 23808 21232 23860
rect 21272 23808 21324 23860
rect 21916 23851 21968 23860
rect 21916 23817 21925 23851
rect 21925 23817 21959 23851
rect 21959 23817 21968 23851
rect 21916 23808 21968 23817
rect 25504 23851 25556 23860
rect 25504 23817 25513 23851
rect 25513 23817 25547 23851
rect 25547 23817 25556 23851
rect 25504 23808 25556 23817
rect 22008 23740 22060 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 26148 23740 26200 23792
rect 21916 23604 21968 23656
rect 25504 23604 25556 23656
rect 8392 23536 8444 23588
rect 3148 23468 3200 23520
rect 8576 23468 8628 23520
rect 9864 23468 9916 23520
rect 10140 23468 10192 23520
rect 10324 23579 10376 23588
rect 10324 23545 10333 23579
rect 10333 23545 10367 23579
rect 10367 23545 10376 23579
rect 12532 23579 12584 23588
rect 10324 23536 10376 23545
rect 12532 23545 12541 23579
rect 12541 23545 12575 23579
rect 12575 23545 12584 23579
rect 12532 23536 12584 23545
rect 12624 23579 12676 23588
rect 12624 23545 12633 23579
rect 12633 23545 12667 23579
rect 12667 23545 12676 23579
rect 12624 23536 12676 23545
rect 14648 23579 14700 23588
rect 14648 23545 14657 23579
rect 14657 23545 14691 23579
rect 14691 23545 14700 23579
rect 14648 23536 14700 23545
rect 15200 23536 15252 23588
rect 10784 23468 10836 23520
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 12256 23468 12308 23520
rect 15384 23468 15436 23520
rect 16580 23468 16632 23520
rect 17960 23468 18012 23520
rect 19340 23468 19392 23520
rect 19524 23468 19576 23520
rect 23480 23468 23532 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 9680 23264 9732 23316
rect 10784 23307 10836 23316
rect 10784 23273 10793 23307
rect 10793 23273 10827 23307
rect 10827 23273 10836 23307
rect 10784 23264 10836 23273
rect 12900 23307 12952 23316
rect 12900 23273 12909 23307
rect 12909 23273 12943 23307
rect 12943 23273 12952 23307
rect 12900 23264 12952 23273
rect 6920 23196 6972 23248
rect 7748 23239 7800 23248
rect 7748 23205 7757 23239
rect 7757 23205 7791 23239
rect 7791 23205 7800 23239
rect 7748 23196 7800 23205
rect 8024 23196 8076 23248
rect 8852 23196 8904 23248
rect 9956 23196 10008 23248
rect 11060 23196 11112 23248
rect 11796 23196 11848 23248
rect 13728 23196 13780 23248
rect 15108 23264 15160 23316
rect 17040 23264 17092 23316
rect 14372 23239 14424 23248
rect 14372 23205 14381 23239
rect 14381 23205 14415 23239
rect 14415 23205 14424 23239
rect 14372 23196 14424 23205
rect 15292 23196 15344 23248
rect 2044 23128 2096 23180
rect 2780 23128 2832 23180
rect 5632 23171 5684 23180
rect 5632 23137 5641 23171
rect 5641 23137 5675 23171
rect 5675 23137 5684 23171
rect 5632 23128 5684 23137
rect 7104 23128 7156 23180
rect 7564 23128 7616 23180
rect 12532 23171 12584 23180
rect 12532 23137 12541 23171
rect 12541 23137 12575 23171
rect 12575 23137 12584 23171
rect 12532 23128 12584 23137
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 10876 22992 10928 23044
rect 13544 23060 13596 23112
rect 16304 23103 16356 23112
rect 15568 22992 15620 23044
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 18512 23128 18564 23180
rect 17224 23060 17276 23112
rect 1584 22924 1636 22976
rect 1676 22924 1728 22976
rect 6092 22924 6144 22976
rect 8668 22967 8720 22976
rect 8668 22933 8677 22967
rect 8677 22933 8711 22967
rect 8711 22933 8720 22967
rect 8668 22924 8720 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2780 22720 2832 22772
rect 7104 22763 7156 22772
rect 7104 22729 7113 22763
rect 7113 22729 7147 22763
rect 7147 22729 7156 22763
rect 7104 22720 7156 22729
rect 8024 22763 8076 22772
rect 8024 22729 8033 22763
rect 8033 22729 8067 22763
rect 8067 22729 8076 22763
rect 8024 22720 8076 22729
rect 9956 22720 10008 22772
rect 11796 22763 11848 22772
rect 11796 22729 11805 22763
rect 11805 22729 11839 22763
rect 11839 22729 11848 22763
rect 11796 22720 11848 22729
rect 12440 22720 12492 22772
rect 13728 22763 13780 22772
rect 13728 22729 13737 22763
rect 13737 22729 13771 22763
rect 13771 22729 13780 22763
rect 13728 22720 13780 22729
rect 17224 22763 17276 22772
rect 17224 22729 17233 22763
rect 17233 22729 17267 22763
rect 17267 22729 17276 22763
rect 17224 22720 17276 22729
rect 9128 22695 9180 22704
rect 9128 22661 9137 22695
rect 9137 22661 9171 22695
rect 9171 22661 9180 22695
rect 9128 22652 9180 22661
rect 9680 22652 9732 22704
rect 2872 22584 2924 22636
rect 8668 22584 8720 22636
rect 9772 22584 9824 22636
rect 10876 22627 10928 22636
rect 1400 22559 1452 22568
rect 1400 22525 1444 22559
rect 1444 22525 1452 22559
rect 1400 22516 1452 22525
rect 2688 22448 2740 22500
rect 2044 22380 2096 22432
rect 2412 22380 2464 22432
rect 3332 22516 3384 22568
rect 10876 22593 10885 22627
rect 10885 22593 10919 22627
rect 10919 22593 10928 22627
rect 10876 22584 10928 22593
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 12624 22584 12676 22636
rect 13176 22627 13228 22636
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 14832 22627 14884 22636
rect 14832 22593 14841 22627
rect 14841 22593 14875 22627
rect 14875 22593 14884 22627
rect 14832 22584 14884 22593
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 16304 22584 16356 22636
rect 3516 22380 3568 22432
rect 8300 22423 8352 22432
rect 8300 22389 8309 22423
rect 8309 22389 8343 22423
rect 8343 22389 8352 22423
rect 10876 22448 10928 22500
rect 11612 22448 11664 22500
rect 14464 22491 14516 22500
rect 8300 22380 8352 22389
rect 12440 22380 12492 22432
rect 14464 22457 14473 22491
rect 14473 22457 14507 22491
rect 14507 22457 14516 22491
rect 14464 22448 14516 22457
rect 15660 22448 15712 22500
rect 13912 22380 13964 22432
rect 15292 22380 15344 22432
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 7748 22219 7800 22228
rect 7748 22185 7757 22219
rect 7757 22185 7791 22219
rect 7791 22185 7800 22219
rect 7748 22176 7800 22185
rect 8300 22219 8352 22228
rect 8300 22185 8309 22219
rect 8309 22185 8343 22219
rect 8343 22185 8352 22219
rect 8300 22176 8352 22185
rect 11336 22176 11388 22228
rect 11888 22219 11940 22228
rect 11888 22185 11897 22219
rect 11897 22185 11931 22219
rect 11931 22185 11940 22219
rect 11888 22176 11940 22185
rect 13544 22176 13596 22228
rect 14372 22176 14424 22228
rect 16212 22219 16264 22228
rect 16212 22185 16221 22219
rect 16221 22185 16255 22219
rect 16255 22185 16264 22219
rect 16212 22176 16264 22185
rect 11060 22151 11112 22160
rect 11060 22117 11069 22151
rect 11069 22117 11103 22151
rect 11103 22117 11112 22151
rect 11060 22108 11112 22117
rect 11612 22151 11664 22160
rect 11612 22117 11621 22151
rect 11621 22117 11655 22151
rect 11655 22117 11664 22151
rect 11612 22108 11664 22117
rect 13820 22108 13872 22160
rect 16488 22151 16540 22160
rect 16488 22117 16497 22151
rect 16497 22117 16531 22151
rect 16531 22117 16540 22151
rect 16488 22108 16540 22117
rect 2320 22040 2372 22092
rect 3056 22083 3108 22092
rect 3056 22049 3074 22083
rect 3074 22049 3108 22083
rect 3056 22040 3108 22049
rect 6552 22040 6604 22092
rect 7472 22040 7524 22092
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 8208 21904 8260 21956
rect 10048 21904 10100 21956
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12992 22083 13044 22092
rect 12440 22040 12492 22049
rect 12992 22049 13001 22083
rect 13001 22049 13035 22083
rect 13035 22049 13044 22083
rect 12992 22040 13044 22049
rect 14188 22083 14240 22092
rect 14188 22049 14232 22083
rect 14232 22049 14240 22083
rect 14188 22040 14240 22049
rect 14740 22040 14792 22092
rect 10784 21972 10836 22024
rect 15476 22040 15528 22092
rect 18236 22083 18288 22092
rect 18236 22049 18245 22083
rect 18245 22049 18279 22083
rect 18279 22049 18288 22083
rect 18236 22040 18288 22049
rect 16028 21972 16080 22024
rect 16396 22015 16448 22024
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16396 21972 16448 21981
rect 16672 22015 16724 22024
rect 16672 21981 16681 22015
rect 16681 21981 16715 22015
rect 16715 21981 16724 22015
rect 16672 21972 16724 21981
rect 11612 21904 11664 21956
rect 15384 21904 15436 21956
rect 2136 21836 2188 21888
rect 3976 21836 4028 21888
rect 6184 21879 6236 21888
rect 6184 21845 6193 21879
rect 6193 21845 6227 21879
rect 6227 21845 6236 21879
rect 6184 21836 6236 21845
rect 15568 21836 15620 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 6552 21675 6604 21684
rect 6552 21641 6561 21675
rect 6561 21641 6595 21675
rect 6595 21641 6604 21675
rect 6552 21632 6604 21641
rect 8576 21632 8628 21684
rect 9128 21632 9180 21684
rect 1952 21564 2004 21616
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 1400 21471 1452 21480
rect 1400 21437 1444 21471
rect 1444 21437 1452 21471
rect 1400 21428 1452 21437
rect 2504 21471 2556 21480
rect 2504 21437 2522 21471
rect 2522 21437 2556 21471
rect 2504 21428 2556 21437
rect 3424 21471 3476 21480
rect 3424 21437 3468 21471
rect 3468 21437 3476 21471
rect 3424 21428 3476 21437
rect 4344 21428 4396 21480
rect 2688 21360 2740 21412
rect 4160 21360 4212 21412
rect 8208 21471 8260 21480
rect 8208 21437 8217 21471
rect 8217 21437 8251 21471
rect 8251 21437 8260 21471
rect 8208 21428 8260 21437
rect 8760 21428 8812 21480
rect 10968 21632 11020 21684
rect 12072 21632 12124 21684
rect 12440 21632 12492 21684
rect 12992 21632 13044 21684
rect 14188 21675 14240 21684
rect 14188 21641 14197 21675
rect 14197 21641 14231 21675
rect 14231 21641 14240 21675
rect 14188 21632 14240 21641
rect 14832 21632 14884 21684
rect 15292 21632 15344 21684
rect 16028 21632 16080 21684
rect 16488 21632 16540 21684
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 10048 21428 10100 21480
rect 12808 21564 12860 21616
rect 15384 21564 15436 21616
rect 16672 21564 16724 21616
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 11428 21428 11480 21480
rect 12808 21428 12860 21480
rect 11520 21403 11572 21412
rect 11520 21369 11529 21403
rect 11529 21369 11563 21403
rect 11563 21369 11572 21403
rect 11520 21360 11572 21369
rect 12624 21360 12676 21412
rect 14648 21428 14700 21480
rect 15660 21428 15712 21480
rect 2320 21335 2372 21344
rect 2320 21301 2329 21335
rect 2329 21301 2363 21335
rect 2363 21301 2372 21335
rect 2320 21292 2372 21301
rect 3056 21292 3108 21344
rect 5448 21292 5500 21344
rect 6000 21292 6052 21344
rect 8024 21335 8076 21344
rect 8024 21301 8033 21335
rect 8033 21301 8067 21335
rect 8067 21301 8076 21335
rect 8024 21292 8076 21301
rect 8392 21292 8444 21344
rect 12716 21335 12768 21344
rect 12716 21301 12725 21335
rect 12725 21301 12759 21335
rect 12759 21301 12768 21335
rect 12716 21292 12768 21301
rect 16580 21292 16632 21344
rect 18236 21292 18288 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 8576 21088 8628 21140
rect 10876 21131 10928 21140
rect 10876 21097 10885 21131
rect 10885 21097 10919 21131
rect 10919 21097 10928 21131
rect 10876 21088 10928 21097
rect 12348 21088 12400 21140
rect 13636 21088 13688 21140
rect 14004 21131 14056 21140
rect 14004 21097 14013 21131
rect 14013 21097 14047 21131
rect 14047 21097 14056 21131
rect 14004 21088 14056 21097
rect 15384 21088 15436 21140
rect 16580 21131 16632 21140
rect 16580 21097 16589 21131
rect 16589 21097 16623 21131
rect 16623 21097 16632 21131
rect 16580 21088 16632 21097
rect 17868 21088 17920 21140
rect 6460 21063 6512 21072
rect 6460 21029 6469 21063
rect 6469 21029 6503 21063
rect 6503 21029 6512 21063
rect 6460 21020 6512 21029
rect 8116 21020 8168 21072
rect 10600 21020 10652 21072
rect 10784 21020 10836 21072
rect 13268 21020 13320 21072
rect 15476 21020 15528 21072
rect 1400 20995 1452 21004
rect 1400 20961 1444 20995
rect 1444 20961 1452 20995
rect 4712 20995 4764 21004
rect 1400 20952 1452 20961
rect 4712 20961 4721 20995
rect 4721 20961 4755 20995
rect 4755 20961 4764 20995
rect 4712 20952 4764 20961
rect 11888 20995 11940 21004
rect 11888 20961 11906 20995
rect 11906 20961 11940 20995
rect 11888 20952 11940 20961
rect 12348 20952 12400 21004
rect 12716 20952 12768 21004
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 1584 20884 1636 20936
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 9956 20927 10008 20936
rect 2504 20748 2556 20800
rect 4620 20748 4672 20800
rect 7472 20748 7524 20800
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 8208 20748 8260 20800
rect 11428 20748 11480 20800
rect 12808 20748 12860 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20544 1452 20596
rect 4712 20544 4764 20596
rect 8484 20544 8536 20596
rect 10968 20544 11020 20596
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 13820 20544 13872 20596
rect 15292 20544 15344 20596
rect 17408 20587 17460 20596
rect 17408 20553 17417 20587
rect 17417 20553 17451 20587
rect 17451 20553 17460 20587
rect 17408 20544 17460 20553
rect 14648 20519 14700 20528
rect 14648 20485 14657 20519
rect 14657 20485 14691 20519
rect 14691 20485 14700 20519
rect 14648 20476 14700 20485
rect 16120 20519 16172 20528
rect 16120 20485 16129 20519
rect 16129 20485 16163 20519
rect 16163 20485 16172 20519
rect 16120 20476 16172 20485
rect 2688 20408 2740 20460
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 8024 20408 8076 20417
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 2320 20340 2372 20392
rect 9772 20383 9824 20392
rect 2228 20272 2280 20324
rect 5908 20315 5960 20324
rect 5908 20281 5917 20315
rect 5917 20281 5951 20315
rect 5951 20281 5960 20315
rect 5908 20272 5960 20281
rect 2688 20204 2740 20256
rect 3424 20247 3476 20256
rect 3424 20213 3433 20247
rect 3433 20213 3467 20247
rect 3467 20213 3476 20247
rect 3424 20204 3476 20213
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 18144 20383 18196 20392
rect 18144 20349 18162 20383
rect 18162 20349 18196 20383
rect 18144 20340 18196 20349
rect 8116 20272 8168 20324
rect 10692 20272 10744 20324
rect 6460 20204 6512 20256
rect 6828 20247 6880 20256
rect 6828 20213 6837 20247
rect 6837 20213 6871 20247
rect 6871 20213 6880 20247
rect 6828 20204 6880 20213
rect 13084 20204 13136 20256
rect 13268 20247 13320 20256
rect 13268 20213 13277 20247
rect 13277 20213 13311 20247
rect 13311 20213 13320 20247
rect 13636 20247 13688 20256
rect 13268 20204 13320 20213
rect 13636 20213 13645 20247
rect 13645 20213 13679 20247
rect 13679 20213 13688 20247
rect 14832 20272 14884 20324
rect 18788 20272 18840 20324
rect 13636 20204 13688 20213
rect 15476 20204 15528 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2872 20000 2924 20052
rect 4160 20000 4212 20052
rect 6368 20043 6420 20052
rect 2596 19932 2648 19984
rect 4804 19975 4856 19984
rect 4804 19941 4813 19975
rect 4813 19941 4847 19975
rect 4847 19941 4856 19975
rect 4804 19932 4856 19941
rect 5080 19932 5132 19984
rect 6368 20009 6377 20043
rect 6377 20009 6411 20043
rect 6411 20009 6420 20043
rect 6368 20000 6420 20009
rect 6736 20000 6788 20052
rect 8116 20043 8168 20052
rect 8116 20009 8125 20043
rect 8125 20009 8159 20043
rect 8159 20009 8168 20043
rect 8116 20000 8168 20009
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 9956 20043 10008 20052
rect 9956 20009 9965 20043
rect 9965 20009 9999 20043
rect 9999 20009 10008 20043
rect 9956 20000 10008 20009
rect 11336 20043 11388 20052
rect 11336 20009 11345 20043
rect 11345 20009 11379 20043
rect 11379 20009 11388 20043
rect 11336 20000 11388 20009
rect 12716 20000 12768 20052
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 5908 19932 5960 19984
rect 7472 19975 7524 19984
rect 7472 19941 7481 19975
rect 7481 19941 7515 19975
rect 7515 19941 7524 19975
rect 7472 19932 7524 19941
rect 6276 19796 6328 19848
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 2320 19771 2372 19780
rect 2320 19737 2329 19771
rect 2329 19737 2363 19771
rect 2363 19737 2372 19771
rect 2320 19728 2372 19737
rect 6552 19728 6604 19780
rect 8392 19864 8444 19916
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 12072 19932 12124 19984
rect 13636 19932 13688 19984
rect 15660 19932 15712 19984
rect 17316 19975 17368 19984
rect 17316 19941 17325 19975
rect 17325 19941 17359 19975
rect 17359 19941 17368 19975
rect 17316 19932 17368 19941
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 18788 19907 18840 19916
rect 18788 19873 18797 19907
rect 18797 19873 18831 19907
rect 18831 19873 18840 19907
rect 18788 19864 18840 19873
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 15476 19796 15528 19848
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 14372 19771 14424 19780
rect 14372 19737 14381 19771
rect 14381 19737 14415 19771
rect 14415 19737 14424 19771
rect 14372 19728 14424 19737
rect 17132 19728 17184 19780
rect 18144 19796 18196 19848
rect 6368 19660 6420 19712
rect 8668 19660 8720 19712
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 12348 19660 12400 19712
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 16580 19703 16632 19712
rect 12440 19660 12492 19669
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 4804 19456 4856 19508
rect 6276 19499 6328 19508
rect 6276 19465 6285 19499
rect 6285 19465 6319 19499
rect 6319 19465 6328 19499
rect 6276 19456 6328 19465
rect 1860 19320 1912 19372
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 2596 19252 2648 19304
rect 3792 19295 3844 19304
rect 3792 19261 3801 19295
rect 3801 19261 3835 19295
rect 3835 19261 3844 19295
rect 3792 19252 3844 19261
rect 4988 19252 5040 19304
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 8576 19252 8628 19304
rect 8760 19252 8812 19304
rect 9956 19456 10008 19508
rect 12072 19456 12124 19508
rect 15660 19499 15712 19508
rect 11152 19320 11204 19372
rect 15660 19465 15669 19499
rect 15669 19465 15703 19499
rect 15703 19465 15712 19499
rect 15660 19456 15712 19465
rect 17316 19456 17368 19508
rect 18788 19456 18840 19508
rect 14372 19388 14424 19440
rect 15476 19388 15528 19440
rect 12164 19252 12216 19304
rect 15568 19320 15620 19372
rect 12532 19252 12584 19304
rect 12992 19252 13044 19304
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 1676 19227 1728 19236
rect 1676 19193 1685 19227
rect 1685 19193 1719 19227
rect 1719 19193 1728 19227
rect 1676 19184 1728 19193
rect 1768 19227 1820 19236
rect 1768 19193 1777 19227
rect 1777 19193 1811 19227
rect 1811 19193 1820 19227
rect 1768 19184 1820 19193
rect 8116 19184 8168 19236
rect 8208 19184 8260 19236
rect 1952 19116 2004 19168
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 4804 19116 4856 19168
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 10692 19184 10744 19236
rect 11704 19184 11756 19236
rect 14556 19227 14608 19236
rect 14556 19193 14565 19227
rect 14565 19193 14599 19227
rect 14599 19193 14608 19227
rect 14556 19184 14608 19193
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 13636 19116 13688 19168
rect 16580 19227 16632 19236
rect 16580 19193 16589 19227
rect 16589 19193 16623 19227
rect 16623 19193 16632 19227
rect 17132 19227 17184 19236
rect 16580 19184 16632 19193
rect 17132 19193 17141 19227
rect 17141 19193 17175 19227
rect 17175 19193 17184 19227
rect 17132 19184 17184 19193
rect 17224 19184 17276 19236
rect 16948 19116 17000 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1768 18912 1820 18964
rect 1952 18912 2004 18964
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 6828 18912 6880 18964
rect 8576 18955 8628 18964
rect 8576 18921 8585 18955
rect 8585 18921 8619 18955
rect 8619 18921 8628 18955
rect 8576 18912 8628 18921
rect 9772 18955 9824 18964
rect 9772 18921 9781 18955
rect 9781 18921 9815 18955
rect 9815 18921 9824 18955
rect 9772 18912 9824 18921
rect 12256 18955 12308 18964
rect 12256 18921 12265 18955
rect 12265 18921 12299 18955
rect 12299 18921 12308 18955
rect 12256 18912 12308 18921
rect 12348 18912 12400 18964
rect 15752 18955 15804 18964
rect 15752 18921 15761 18955
rect 15761 18921 15795 18955
rect 15795 18921 15804 18955
rect 15752 18912 15804 18921
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 2688 18844 2740 18896
rect 4620 18887 4672 18896
rect 4620 18853 4629 18887
rect 4629 18853 4663 18887
rect 4663 18853 4672 18887
rect 4620 18844 4672 18853
rect 11704 18887 11756 18896
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 6184 18776 6236 18828
rect 7380 18776 7432 18828
rect 11704 18853 11707 18887
rect 11707 18853 11741 18887
rect 11741 18853 11756 18887
rect 11704 18844 11756 18853
rect 16028 18887 16080 18896
rect 16028 18853 16037 18887
rect 16037 18853 16071 18887
rect 16071 18853 16080 18887
rect 16028 18844 16080 18853
rect 17132 18844 17184 18896
rect 17500 18844 17552 18896
rect 18144 18887 18196 18896
rect 18144 18853 18153 18887
rect 18153 18853 18187 18887
rect 18187 18853 18196 18887
rect 18144 18844 18196 18853
rect 8024 18819 8076 18828
rect 8024 18785 8033 18819
rect 8033 18785 8067 18819
rect 8067 18785 8076 18819
rect 8024 18776 8076 18785
rect 9496 18776 9548 18828
rect 10048 18776 10100 18828
rect 10140 18776 10192 18828
rect 10876 18776 10928 18828
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 12808 18776 12860 18828
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 13176 18776 13228 18828
rect 1768 18708 1820 18760
rect 4528 18751 4580 18760
rect 4528 18717 4537 18751
rect 4537 18717 4571 18751
rect 4571 18717 4580 18751
rect 4528 18708 4580 18717
rect 15292 18708 15344 18760
rect 17868 18708 17920 18760
rect 2596 18683 2648 18692
rect 2596 18649 2605 18683
rect 2605 18649 2639 18683
rect 2639 18649 2648 18683
rect 2596 18640 2648 18649
rect 5080 18683 5132 18692
rect 5080 18649 5089 18683
rect 5089 18649 5123 18683
rect 5123 18649 5132 18683
rect 5080 18640 5132 18649
rect 9036 18640 9088 18692
rect 5540 18615 5592 18624
rect 5540 18581 5549 18615
rect 5549 18581 5583 18615
rect 5583 18581 5592 18615
rect 5540 18572 5592 18581
rect 6184 18615 6236 18624
rect 6184 18581 6193 18615
rect 6193 18581 6227 18615
rect 6227 18581 6236 18615
rect 6184 18572 6236 18581
rect 9220 18572 9272 18624
rect 11060 18572 11112 18624
rect 11244 18615 11296 18624
rect 11244 18581 11253 18615
rect 11253 18581 11287 18615
rect 11287 18581 11296 18615
rect 11244 18572 11296 18581
rect 13912 18572 13964 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 4620 18368 4672 18420
rect 7380 18411 7432 18420
rect 7380 18377 7389 18411
rect 7389 18377 7423 18411
rect 7423 18377 7432 18411
rect 7380 18368 7432 18377
rect 8760 18368 8812 18420
rect 13084 18411 13136 18420
rect 13084 18377 13093 18411
rect 13093 18377 13127 18411
rect 13127 18377 13136 18411
rect 13084 18368 13136 18377
rect 14832 18411 14884 18420
rect 14832 18377 14841 18411
rect 14841 18377 14875 18411
rect 14875 18377 14884 18411
rect 14832 18368 14884 18377
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 2412 18343 2464 18352
rect 2412 18309 2421 18343
rect 2421 18309 2455 18343
rect 2455 18309 2464 18343
rect 2412 18300 2464 18309
rect 9220 18343 9272 18352
rect 9220 18309 9244 18343
rect 9244 18309 9272 18343
rect 9220 18300 9272 18309
rect 10048 18300 10100 18352
rect 11060 18300 11112 18352
rect 15200 18343 15252 18352
rect 15200 18309 15209 18343
rect 15209 18309 15243 18343
rect 15243 18309 15252 18343
rect 15200 18300 15252 18309
rect 15568 18300 15620 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 2780 18232 2832 18284
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 3792 18275 3844 18284
rect 3792 18241 3801 18275
rect 3801 18241 3835 18275
rect 3835 18241 3844 18275
rect 3792 18232 3844 18241
rect 4068 18232 4120 18284
rect 8852 18232 8904 18284
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 7748 18207 7800 18216
rect 7748 18173 7757 18207
rect 7757 18173 7791 18207
rect 7791 18173 7800 18207
rect 7748 18164 7800 18173
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 9128 18164 9180 18216
rect 1952 18139 2004 18148
rect 1952 18105 1961 18139
rect 1961 18105 1995 18139
rect 1995 18105 2004 18139
rect 1952 18096 2004 18105
rect 3516 18139 3568 18148
rect 3516 18105 3525 18139
rect 3525 18105 3559 18139
rect 3559 18105 3568 18139
rect 3516 18096 3568 18105
rect 4896 18139 4948 18148
rect 4896 18105 4905 18139
rect 4905 18105 4939 18139
rect 4939 18105 4948 18139
rect 4896 18096 4948 18105
rect 6368 18096 6420 18148
rect 2688 18028 2740 18080
rect 6000 18028 6052 18080
rect 6920 18028 6972 18080
rect 8852 18071 8904 18080
rect 8852 18037 8861 18071
rect 8861 18037 8895 18071
rect 8895 18037 8904 18071
rect 8852 18028 8904 18037
rect 9036 18139 9088 18148
rect 9036 18105 9045 18139
rect 9045 18105 9079 18139
rect 9079 18105 9088 18139
rect 9036 18096 9088 18105
rect 10692 18096 10744 18148
rect 9588 18028 9640 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 10140 18028 10192 18080
rect 11244 18232 11296 18284
rect 11796 18232 11848 18284
rect 13176 18232 13228 18284
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 16028 18232 16080 18284
rect 12532 18164 12584 18216
rect 13912 18207 13964 18216
rect 13912 18173 13921 18207
rect 13921 18173 13955 18207
rect 13955 18173 13964 18207
rect 13912 18164 13964 18173
rect 16580 18164 16632 18216
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 11704 18139 11756 18148
rect 11704 18105 11713 18139
rect 11713 18105 11747 18139
rect 11747 18105 11756 18139
rect 11704 18096 11756 18105
rect 12440 18028 12492 18080
rect 13636 18028 13688 18080
rect 15108 18096 15160 18148
rect 17224 18096 17276 18148
rect 17500 18071 17552 18080
rect 17500 18037 17509 18071
rect 17509 18037 17543 18071
rect 17543 18037 17552 18071
rect 17500 18028 17552 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 4528 17867 4580 17876
rect 4528 17833 4537 17867
rect 4537 17833 4571 17867
rect 4571 17833 4580 17867
rect 4528 17824 4580 17833
rect 7748 17824 7800 17876
rect 1584 17756 1636 17808
rect 1860 17799 1912 17808
rect 1860 17765 1869 17799
rect 1869 17765 1903 17799
rect 1903 17765 1912 17799
rect 2412 17799 2464 17808
rect 1860 17756 1912 17765
rect 2412 17765 2421 17799
rect 2421 17765 2455 17799
rect 2455 17765 2464 17799
rect 2412 17756 2464 17765
rect 4712 17756 4764 17808
rect 4988 17756 5040 17808
rect 7932 17799 7984 17808
rect 7932 17765 7935 17799
rect 7935 17765 7969 17799
rect 7969 17765 7984 17799
rect 8300 17824 8352 17876
rect 9496 17867 9548 17876
rect 9496 17833 9505 17867
rect 9505 17833 9539 17867
rect 9539 17833 9548 17867
rect 9496 17824 9548 17833
rect 9680 17824 9732 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 11336 17867 11388 17876
rect 10692 17824 10744 17833
rect 11336 17833 11345 17867
rect 11345 17833 11379 17867
rect 11379 17833 11388 17867
rect 11336 17824 11388 17833
rect 12164 17867 12216 17876
rect 12164 17833 12173 17867
rect 12173 17833 12207 17867
rect 12207 17833 12216 17867
rect 12164 17824 12216 17833
rect 7932 17756 7984 17765
rect 11244 17756 11296 17808
rect 12440 17824 12492 17876
rect 13176 17867 13228 17876
rect 13176 17833 13185 17867
rect 13185 17833 13219 17867
rect 13219 17833 13228 17867
rect 13176 17824 13228 17833
rect 15108 17824 15160 17876
rect 16488 17824 16540 17876
rect 17500 17867 17552 17876
rect 17500 17833 17509 17867
rect 17509 17833 17543 17867
rect 17543 17833 17552 17867
rect 17500 17824 17552 17833
rect 18144 17867 18196 17876
rect 18144 17833 18153 17867
rect 18153 17833 18187 17867
rect 18187 17833 18196 17867
rect 18144 17824 18196 17833
rect 13636 17756 13688 17808
rect 15660 17799 15712 17808
rect 15660 17765 15663 17799
rect 15663 17765 15697 17799
rect 15697 17765 15712 17799
rect 15660 17756 15712 17765
rect 10692 17688 10744 17740
rect 11888 17731 11940 17740
rect 11888 17697 11897 17731
rect 11897 17697 11931 17731
rect 11931 17697 11940 17731
rect 11888 17688 11940 17697
rect 13176 17688 13228 17740
rect 17316 17731 17368 17740
rect 17316 17697 17325 17731
rect 17325 17697 17359 17731
rect 17359 17697 17368 17731
rect 17316 17688 17368 17697
rect 18696 17731 18748 17740
rect 18696 17697 18714 17731
rect 18714 17697 18748 17731
rect 18696 17688 18748 17697
rect 4896 17663 4948 17672
rect 4896 17629 4905 17663
rect 4905 17629 4939 17663
rect 4939 17629 4948 17663
rect 4896 17620 4948 17629
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 9772 17620 9824 17672
rect 10140 17620 10192 17672
rect 13268 17620 13320 17672
rect 15476 17620 15528 17672
rect 5540 17484 5592 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 10048 17484 10100 17536
rect 11152 17484 11204 17536
rect 12900 17484 12952 17536
rect 18144 17484 18196 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1860 17280 1912 17332
rect 3516 17280 3568 17332
rect 7564 17280 7616 17332
rect 8484 17323 8536 17332
rect 8484 17289 8493 17323
rect 8493 17289 8527 17323
rect 8527 17289 8536 17323
rect 8484 17280 8536 17289
rect 10048 17280 10100 17332
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 10876 17280 10928 17332
rect 11152 17280 11204 17332
rect 11888 17280 11940 17332
rect 12440 17280 12492 17332
rect 13636 17323 13688 17332
rect 13636 17289 13645 17323
rect 13645 17289 13679 17323
rect 13679 17289 13688 17323
rect 13636 17280 13688 17289
rect 17316 17280 17368 17332
rect 19064 17280 19116 17332
rect 2044 17144 2096 17196
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 2228 17008 2280 17060
rect 17684 17212 17736 17264
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 4896 17144 4948 17196
rect 7104 17144 7156 17196
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 3332 17119 3384 17128
rect 3332 17085 3341 17119
rect 3341 17085 3375 17119
rect 3375 17085 3384 17119
rect 4068 17119 4120 17128
rect 3332 17076 3384 17085
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 5540 17076 5592 17128
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 9404 17076 9456 17128
rect 9956 17076 10008 17128
rect 12900 17076 12952 17128
rect 13176 17076 13228 17128
rect 7932 17051 7984 17060
rect 7932 17017 7935 17051
rect 7935 17017 7969 17051
rect 7969 17017 7984 17051
rect 7932 17008 7984 17017
rect 9128 17008 9180 17060
rect 9588 17008 9640 17060
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 14648 17076 14700 17085
rect 15844 17076 15896 17128
rect 18144 17076 18196 17128
rect 4988 16940 5040 16992
rect 10140 16940 10192 16992
rect 11796 16983 11848 16992
rect 11796 16949 11805 16983
rect 11805 16949 11839 16983
rect 11839 16949 11848 16983
rect 11796 16940 11848 16949
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 15660 16983 15712 16992
rect 15660 16949 15669 16983
rect 15669 16949 15703 16983
rect 15703 16949 15712 16983
rect 15660 16940 15712 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16736 1636 16788
rect 2688 16736 2740 16788
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 4896 16736 4948 16788
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 9864 16779 9916 16788
rect 9864 16745 9873 16779
rect 9873 16745 9907 16779
rect 9907 16745 9916 16779
rect 9864 16736 9916 16745
rect 13084 16736 13136 16788
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 15844 16779 15896 16788
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 2044 16668 2096 16720
rect 2228 16643 2280 16652
rect 2228 16609 2237 16643
rect 2237 16609 2271 16643
rect 2271 16609 2280 16643
rect 2228 16600 2280 16609
rect 2596 16668 2648 16720
rect 3240 16668 3292 16720
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 4896 16600 4948 16652
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 6920 16668 6972 16720
rect 11244 16668 11296 16720
rect 11612 16668 11664 16720
rect 13820 16711 13872 16720
rect 13820 16677 13829 16711
rect 13829 16677 13863 16711
rect 13863 16677 13872 16711
rect 13820 16668 13872 16677
rect 15476 16711 15528 16720
rect 15476 16677 15485 16711
rect 15485 16677 15519 16711
rect 15519 16677 15528 16711
rect 15476 16668 15528 16677
rect 15752 16668 15804 16720
rect 17960 16711 18012 16720
rect 17960 16677 17969 16711
rect 17969 16677 18003 16711
rect 18003 16677 18012 16711
rect 17960 16668 18012 16677
rect 4344 16532 4396 16584
rect 6368 16600 6420 16652
rect 6644 16600 6696 16652
rect 7472 16600 7524 16652
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 8392 16600 8444 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 12164 16600 12216 16652
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 13544 16600 13596 16652
rect 19340 16643 19392 16652
rect 9588 16532 9640 16584
rect 9772 16532 9824 16584
rect 11520 16532 11572 16584
rect 11796 16532 11848 16584
rect 14188 16532 14240 16584
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 16672 16532 16724 16584
rect 17040 16532 17092 16584
rect 17684 16532 17736 16584
rect 18604 16532 18656 16584
rect 7840 16464 7892 16516
rect 9404 16464 9456 16516
rect 8760 16396 8812 16448
rect 10048 16396 10100 16448
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 10692 16396 10744 16448
rect 10876 16396 10928 16448
rect 11244 16439 11296 16448
rect 11244 16405 11268 16439
rect 11268 16405 11296 16439
rect 11244 16396 11296 16405
rect 11336 16439 11388 16448
rect 11336 16405 11345 16439
rect 11345 16405 11379 16439
rect 11379 16405 11388 16439
rect 11336 16396 11388 16405
rect 19524 16439 19576 16448
rect 19524 16405 19533 16439
rect 19533 16405 19567 16439
rect 19567 16405 19576 16439
rect 19524 16396 19576 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2228 16192 2280 16244
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 9404 16192 9456 16244
rect 9680 16192 9732 16244
rect 10968 16192 11020 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 19340 16235 19392 16244
rect 19340 16201 19349 16235
rect 19349 16201 19383 16235
rect 19383 16201 19392 16235
rect 19340 16192 19392 16201
rect 3792 16167 3844 16176
rect 3792 16133 3801 16167
rect 3801 16133 3835 16167
rect 3835 16133 3844 16167
rect 3792 16124 3844 16133
rect 5540 16167 5592 16176
rect 5540 16133 5549 16167
rect 5549 16133 5583 16167
rect 5583 16133 5592 16167
rect 5540 16124 5592 16133
rect 9128 16167 9180 16176
rect 9128 16133 9137 16167
rect 9137 16133 9171 16167
rect 9171 16133 9180 16167
rect 9128 16124 9180 16133
rect 9588 16124 9640 16176
rect 11336 16124 11388 16176
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 1952 16056 2004 16108
rect 3240 16099 3292 16108
rect 3240 16065 3249 16099
rect 3249 16065 3283 16099
rect 3283 16065 3292 16099
rect 3240 16056 3292 16065
rect 5356 16056 5408 16108
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 7656 16056 7708 16108
rect 8668 16056 8720 16108
rect 8852 16056 8904 16108
rect 10140 16056 10192 16108
rect 1768 15920 1820 15972
rect 2688 15920 2740 15972
rect 3332 15963 3384 15972
rect 3332 15929 3341 15963
rect 3341 15929 3375 15963
rect 3375 15929 3384 15963
rect 3332 15920 3384 15929
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 7012 15920 7064 15972
rect 7380 15920 7432 15972
rect 8668 15920 8720 15972
rect 9220 15920 9272 15972
rect 6368 15852 6420 15904
rect 7288 15852 7340 15904
rect 7564 15895 7616 15904
rect 7564 15861 7573 15895
rect 7573 15861 7607 15895
rect 7607 15861 7616 15895
rect 7564 15852 7616 15861
rect 10048 15852 10100 15904
rect 11060 16056 11112 16108
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 10508 15988 10560 16040
rect 11704 15988 11756 16040
rect 12900 15988 12952 16040
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 13820 15988 13872 16040
rect 10692 15920 10744 15972
rect 11244 15920 11296 15972
rect 12624 15920 12676 15972
rect 15660 15920 15712 15972
rect 16580 15963 16632 15972
rect 16580 15929 16589 15963
rect 16589 15929 16623 15963
rect 16623 15929 16632 15963
rect 16580 15920 16632 15929
rect 11612 15852 11664 15904
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 15108 15852 15160 15904
rect 15752 15852 15804 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 4068 15648 4120 15700
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 5356 15648 5408 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 6920 15648 6972 15700
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 2596 15580 2648 15632
rect 3976 15512 4028 15564
rect 6092 15512 6144 15564
rect 6184 15512 6236 15564
rect 8024 15580 8076 15632
rect 10692 15580 10744 15632
rect 8208 15555 8260 15564
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 5632 15444 5684 15496
rect 6368 15487 6420 15496
rect 6368 15453 6377 15487
rect 6377 15453 6411 15487
rect 6411 15453 6420 15487
rect 6368 15444 6420 15453
rect 6736 15444 6788 15496
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 11704 15555 11756 15564
rect 11704 15521 11710 15555
rect 11710 15521 11756 15555
rect 11704 15512 11756 15521
rect 12072 15512 12124 15564
rect 10048 15444 10100 15496
rect 11152 15444 11204 15496
rect 11520 15444 11572 15496
rect 12348 15580 12400 15632
rect 12440 15512 12492 15564
rect 12716 15444 12768 15496
rect 8208 15376 8260 15428
rect 9128 15376 9180 15428
rect 13452 15512 13504 15564
rect 14188 15648 14240 15700
rect 15660 15623 15712 15632
rect 15660 15589 15663 15623
rect 15663 15589 15697 15623
rect 15697 15589 15712 15623
rect 15660 15580 15712 15589
rect 16488 15580 16540 15632
rect 16580 15580 16632 15632
rect 15752 15512 15804 15564
rect 17500 15555 17552 15564
rect 17500 15521 17509 15555
rect 17509 15521 17543 15555
rect 17543 15521 17552 15555
rect 17500 15512 17552 15521
rect 16120 15444 16172 15496
rect 16672 15444 16724 15496
rect 13912 15376 13964 15428
rect 1768 15308 1820 15360
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 5080 15308 5132 15360
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 9220 15308 9272 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 13820 15308 13872 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 4896 15147 4948 15156
rect 4896 15113 4905 15147
rect 4905 15113 4939 15147
rect 4939 15113 4948 15147
rect 4896 15104 4948 15113
rect 4988 15104 5040 15156
rect 5448 15104 5500 15156
rect 6092 15104 6144 15156
rect 6644 15147 6696 15156
rect 3240 15036 3292 15088
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 12072 15147 12124 15156
rect 12072 15113 12081 15147
rect 12081 15113 12115 15147
rect 12115 15113 12124 15147
rect 12072 15104 12124 15113
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 2780 14968 2832 15020
rect 5448 14968 5500 15020
rect 13728 14968 13780 15020
rect 15292 14968 15344 15020
rect 17868 15036 17920 15088
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 2596 14900 2648 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7012 14900 7064 14909
rect 2228 14832 2280 14884
rect 2964 14832 3016 14884
rect 3240 14875 3292 14884
rect 3240 14841 3249 14875
rect 3249 14841 3283 14875
rect 3283 14841 3292 14875
rect 3240 14832 3292 14841
rect 4896 14832 4948 14884
rect 7012 14764 7064 14816
rect 8760 14764 8812 14816
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 16672 14943 16724 14952
rect 16672 14909 16681 14943
rect 16681 14909 16715 14943
rect 16715 14909 16724 14943
rect 16672 14900 16724 14909
rect 9956 14832 10008 14884
rect 10140 14832 10192 14884
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 11796 14764 11848 14816
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 16488 14764 16540 14816
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 3148 14560 3200 14612
rect 3976 14560 4028 14612
rect 5264 14560 5316 14612
rect 6644 14603 6696 14612
rect 6644 14569 6653 14603
rect 6653 14569 6687 14603
rect 6687 14569 6696 14603
rect 6644 14560 6696 14569
rect 7748 14603 7800 14612
rect 7748 14569 7757 14603
rect 7757 14569 7791 14603
rect 7791 14569 7800 14603
rect 7748 14560 7800 14569
rect 11796 14560 11848 14612
rect 12716 14603 12768 14612
rect 12716 14569 12725 14603
rect 12725 14569 12759 14603
rect 12759 14569 12768 14603
rect 12716 14560 12768 14569
rect 13176 14560 13228 14612
rect 14004 14603 14056 14612
rect 14004 14569 14013 14603
rect 14013 14569 14047 14603
rect 14047 14569 14056 14603
rect 14004 14560 14056 14569
rect 16120 14603 16172 14612
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 16856 14603 16908 14612
rect 16856 14569 16865 14603
rect 16865 14569 16899 14603
rect 16899 14569 16908 14603
rect 16856 14560 16908 14569
rect 6092 14535 6144 14544
rect 6092 14501 6095 14535
rect 6095 14501 6129 14535
rect 6129 14501 6144 14535
rect 6092 14492 6144 14501
rect 9680 14535 9732 14544
rect 9680 14501 9689 14535
rect 9689 14501 9723 14535
rect 9723 14501 9732 14535
rect 9680 14492 9732 14501
rect 15844 14535 15896 14544
rect 2596 14424 2648 14476
rect 3240 14424 3292 14476
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 6184 14424 6236 14476
rect 6828 14424 6880 14476
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 9956 14424 10008 14476
rect 11980 14467 12032 14476
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 9772 14356 9824 14408
rect 10140 14356 10192 14408
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 12624 14424 12676 14476
rect 15844 14501 15853 14535
rect 15853 14501 15887 14535
rect 15887 14501 15896 14535
rect 15844 14492 15896 14501
rect 15384 14424 15436 14476
rect 11888 14356 11940 14408
rect 12808 14356 12860 14408
rect 9128 14331 9180 14340
rect 9128 14297 9137 14331
rect 9137 14297 9171 14331
rect 9171 14297 9180 14331
rect 9128 14288 9180 14297
rect 4068 14220 4120 14272
rect 5080 14220 5132 14272
rect 8944 14220 8996 14272
rect 10324 14288 10376 14340
rect 12440 14288 12492 14340
rect 16580 14424 16632 14476
rect 10048 14220 10100 14272
rect 11152 14263 11204 14272
rect 11152 14229 11161 14263
rect 11161 14229 11195 14263
rect 11195 14229 11204 14263
rect 11152 14220 11204 14229
rect 15384 14288 15436 14340
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2596 14059 2648 14068
rect 2596 14025 2605 14059
rect 2605 14025 2639 14059
rect 2639 14025 2648 14059
rect 2596 14016 2648 14025
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 7656 14016 7708 14068
rect 8208 14016 8260 14068
rect 10968 14016 11020 14068
rect 11980 14016 12032 14068
rect 4896 13948 4948 14000
rect 6092 13948 6144 14000
rect 6828 13948 6880 14000
rect 8944 13991 8996 14000
rect 8944 13957 8953 13991
rect 8953 13957 8987 13991
rect 8987 13957 8996 13991
rect 8944 13948 8996 13957
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 6460 13855 6512 13864
rect 1584 13787 1636 13796
rect 1584 13753 1593 13787
rect 1593 13753 1627 13787
rect 1627 13753 1636 13787
rect 1584 13744 1636 13753
rect 1676 13787 1728 13796
rect 1676 13753 1685 13787
rect 1685 13753 1719 13787
rect 1719 13753 1728 13787
rect 6460 13821 6469 13855
rect 6469 13821 6503 13855
rect 6503 13821 6512 13855
rect 6460 13812 6512 13821
rect 7564 13812 7616 13864
rect 8208 13812 8260 13864
rect 9128 13812 9180 13864
rect 3240 13787 3292 13796
rect 1676 13744 1728 13753
rect 3240 13753 3249 13787
rect 3249 13753 3283 13787
rect 3283 13753 3292 13787
rect 3240 13744 3292 13753
rect 4896 13744 4948 13796
rect 8668 13787 8720 13796
rect 8668 13753 8677 13787
rect 8677 13753 8711 13787
rect 8711 13753 8720 13787
rect 8668 13744 8720 13753
rect 9956 13948 10008 14000
rect 11244 13948 11296 14000
rect 12164 13948 12216 14000
rect 13084 13948 13136 14000
rect 13820 14016 13872 14068
rect 15752 14059 15804 14068
rect 15752 14025 15761 14059
rect 15761 14025 15795 14059
rect 15795 14025 15804 14059
rect 15752 14016 15804 14025
rect 16580 14016 16632 14068
rect 9680 13880 9732 13932
rect 10324 13880 10376 13932
rect 14004 13880 14056 13932
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 15384 13923 15436 13932
rect 14464 13880 14516 13889
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 15476 13880 15528 13932
rect 10232 13855 10284 13864
rect 10232 13821 10241 13855
rect 10241 13821 10275 13855
rect 10275 13821 10284 13855
rect 10692 13855 10744 13864
rect 10232 13812 10284 13821
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 11888 13812 11940 13864
rect 13084 13855 13136 13864
rect 11060 13744 11112 13796
rect 12808 13744 12860 13796
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 14004 13787 14056 13796
rect 14004 13753 14013 13787
rect 14013 13753 14047 13787
rect 14047 13753 14056 13787
rect 14004 13744 14056 13753
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 9588 13676 9640 13728
rect 9956 13676 10008 13728
rect 10140 13676 10192 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1952 13472 2004 13524
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 6184 13472 6236 13524
rect 7564 13472 7616 13524
rect 9588 13472 9640 13524
rect 11336 13515 11388 13524
rect 11336 13481 11345 13515
rect 11345 13481 11379 13515
rect 11379 13481 11388 13515
rect 11336 13472 11388 13481
rect 11428 13472 11480 13524
rect 12624 13472 12676 13524
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 14004 13472 14056 13524
rect 2596 13447 2648 13456
rect 2596 13413 2605 13447
rect 2605 13413 2639 13447
rect 2639 13413 2648 13447
rect 2596 13404 2648 13413
rect 4896 13404 4948 13456
rect 7104 13404 7156 13456
rect 12440 13404 12492 13456
rect 15568 13447 15620 13456
rect 15568 13413 15577 13447
rect 15577 13413 15611 13447
rect 15611 13413 15620 13447
rect 15568 13404 15620 13413
rect 9588 13336 9640 13388
rect 10876 13336 10928 13388
rect 11612 13336 11664 13388
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 2872 13268 2924 13320
rect 3424 13268 3476 13320
rect 5264 13268 5316 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 7564 13268 7616 13320
rect 9680 13268 9732 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10968 13268 11020 13320
rect 11152 13268 11204 13320
rect 11980 13268 12032 13320
rect 3056 13243 3108 13252
rect 3056 13209 3065 13243
rect 3065 13209 3099 13243
rect 3099 13209 3108 13243
rect 3056 13200 3108 13209
rect 10692 13200 10744 13252
rect 1584 13132 1636 13184
rect 2504 13132 2556 13184
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 9956 13132 10008 13184
rect 10600 13132 10652 13184
rect 12256 13200 12308 13252
rect 11520 13132 11572 13184
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2596 12928 2648 12980
rect 4160 12928 4212 12980
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 5540 12971 5592 12980
rect 5540 12937 5549 12971
rect 5549 12937 5583 12971
rect 5583 12937 5592 12971
rect 5540 12928 5592 12937
rect 6920 12928 6972 12980
rect 7104 12928 7156 12980
rect 8392 12928 8444 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 11520 12928 11572 12980
rect 11704 12928 11756 12980
rect 12440 12928 12492 12980
rect 13084 12971 13136 12980
rect 13084 12937 13093 12971
rect 13093 12937 13127 12971
rect 13127 12937 13136 12971
rect 13084 12928 13136 12937
rect 13636 12928 13688 12980
rect 2872 12903 2924 12912
rect 2872 12869 2881 12903
rect 2881 12869 2915 12903
rect 2915 12869 2924 12903
rect 2872 12860 2924 12869
rect 10324 12860 10376 12912
rect 11244 12860 11296 12912
rect 13176 12860 13228 12912
rect 3056 12792 3108 12844
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7380 12792 7432 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 10692 12724 10744 12776
rect 11796 12724 11848 12776
rect 13912 12724 13964 12776
rect 2320 12699 2372 12708
rect 2320 12665 2329 12699
rect 2329 12665 2363 12699
rect 2363 12665 2372 12699
rect 2320 12656 2372 12665
rect 2688 12656 2740 12708
rect 3884 12699 3936 12708
rect 3884 12665 3893 12699
rect 3893 12665 3927 12699
rect 3927 12665 3936 12699
rect 3884 12656 3936 12665
rect 4068 12656 4120 12708
rect 6920 12656 6972 12708
rect 7932 12656 7984 12708
rect 8300 12656 8352 12708
rect 12716 12656 12768 12708
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 10692 12588 10744 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3792 12384 3844 12436
rect 4620 12427 4672 12436
rect 4620 12393 4629 12427
rect 4629 12393 4663 12427
rect 4663 12393 4672 12427
rect 4620 12384 4672 12393
rect 6736 12384 6788 12436
rect 7104 12384 7156 12436
rect 9128 12384 9180 12436
rect 9956 12427 10008 12436
rect 9956 12393 9965 12427
rect 9965 12393 9999 12427
rect 9999 12393 10008 12427
rect 9956 12384 10008 12393
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 12532 12384 12584 12436
rect 13820 12384 13872 12436
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 2872 12248 2924 12300
rect 3884 12291 3936 12300
rect 3884 12257 3893 12291
rect 3893 12257 3927 12291
rect 3927 12257 3936 12291
rect 3884 12248 3936 12257
rect 4160 12248 4212 12300
rect 4344 12248 4396 12300
rect 7932 12316 7984 12368
rect 10968 12316 11020 12368
rect 13176 12359 13228 12368
rect 13176 12325 13185 12359
rect 13185 12325 13219 12359
rect 13219 12325 13228 12359
rect 13176 12316 13228 12325
rect 6092 12248 6144 12300
rect 6276 12248 6328 12300
rect 12164 12291 12216 12300
rect 12164 12257 12173 12291
rect 12173 12257 12207 12291
rect 12207 12257 12216 12291
rect 12164 12248 12216 12257
rect 13084 12248 13136 12300
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 7380 12180 7432 12232
rect 7748 12180 7800 12232
rect 10140 12180 10192 12232
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 1492 12044 1544 12096
rect 1952 12044 2004 12096
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 6736 12044 6788 12096
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 8852 12087 8904 12096
rect 8852 12053 8861 12087
rect 8861 12053 8895 12087
rect 8895 12053 8904 12087
rect 8852 12044 8904 12053
rect 11152 12044 11204 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 6092 11840 6144 11892
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 10416 11840 10468 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 12808 11840 12860 11892
rect 13084 11840 13136 11892
rect 11980 11772 12032 11824
rect 2412 11704 2464 11756
rect 2688 11704 2740 11756
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 4620 11704 4672 11713
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 8852 11704 8904 11756
rect 10692 11636 10744 11688
rect 11244 11636 11296 11688
rect 12808 11636 12860 11688
rect 1492 11611 1544 11620
rect 1492 11577 1501 11611
rect 1501 11577 1535 11611
rect 1535 11577 1544 11611
rect 1492 11568 1544 11577
rect 1400 11500 1452 11552
rect 2688 11568 2740 11620
rect 4896 11568 4948 11620
rect 6736 11568 6788 11620
rect 7012 11611 7064 11620
rect 7012 11577 7021 11611
rect 7021 11577 7055 11611
rect 7055 11577 7064 11611
rect 8576 11611 8628 11620
rect 7012 11568 7064 11577
rect 8576 11577 8585 11611
rect 8585 11577 8619 11611
rect 8619 11577 8628 11611
rect 8576 11568 8628 11577
rect 8760 11568 8812 11620
rect 10968 11611 11020 11620
rect 10968 11577 10971 11611
rect 10971 11577 11005 11611
rect 11005 11577 11020 11611
rect 10968 11568 11020 11577
rect 16488 11568 16540 11620
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 2964 11500 3016 11552
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 9496 11500 9548 11552
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3056 11296 3108 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 9128 11296 9180 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 2136 11271 2188 11280
rect 2136 11237 2145 11271
rect 2145 11237 2179 11271
rect 2179 11237 2188 11271
rect 2136 11228 2188 11237
rect 4896 11271 4948 11280
rect 4896 11237 4899 11271
rect 4899 11237 4933 11271
rect 4933 11237 4948 11271
rect 4896 11228 4948 11237
rect 7932 11228 7984 11280
rect 8392 11228 8444 11280
rect 8760 11228 8812 11280
rect 11152 11228 11204 11280
rect 11888 11228 11940 11280
rect 3148 11160 3200 11212
rect 5540 11160 5592 11212
rect 2504 11092 2556 11144
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 8208 11092 8260 11144
rect 10784 11092 10836 11144
rect 11980 11092 12032 11144
rect 1400 11024 1452 11076
rect 2964 11067 3016 11076
rect 2964 11033 2973 11067
rect 2973 11033 3007 11067
rect 3007 11033 3016 11067
rect 2964 11024 3016 11033
rect 6184 11067 6236 11076
rect 6184 11033 6193 11067
rect 6193 11033 6227 11067
rect 6227 11033 6236 11067
rect 6184 11024 6236 11033
rect 8300 10956 8352 11008
rect 8668 10956 8720 11008
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 11060 10956 11112 11008
rect 11704 10956 11756 11008
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 3608 10795 3660 10804
rect 3608 10761 3617 10795
rect 3617 10761 3651 10795
rect 3651 10761 3660 10795
rect 3608 10752 3660 10761
rect 4896 10752 4948 10804
rect 5540 10752 5592 10804
rect 8668 10795 8720 10804
rect 8668 10761 8692 10795
rect 8692 10761 8720 10795
rect 8668 10752 8720 10761
rect 9128 10752 9180 10804
rect 2504 10727 2556 10736
rect 2504 10693 2513 10727
rect 2513 10693 2547 10727
rect 2547 10693 2556 10727
rect 2504 10684 2556 10693
rect 5080 10684 5132 10736
rect 8760 10727 8812 10736
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 1308 10480 1360 10532
rect 9312 10684 9364 10736
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 5080 10548 5132 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 8300 10548 8352 10600
rect 9956 10616 10008 10668
rect 11980 10616 12032 10668
rect 11060 10548 11112 10600
rect 11152 10591 11204 10600
rect 11152 10557 11161 10591
rect 11161 10557 11195 10591
rect 11195 10557 11204 10591
rect 12808 10591 12860 10600
rect 11152 10548 11204 10557
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 10140 10523 10192 10532
rect 2044 10480 2096 10489
rect 10140 10489 10149 10523
rect 10149 10489 10183 10523
rect 10183 10489 10192 10523
rect 10140 10480 10192 10489
rect 4528 10412 4580 10464
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 7012 10412 7064 10464
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2136 10208 2188 10260
rect 4436 10251 4488 10260
rect 4436 10217 4445 10251
rect 4445 10217 4479 10251
rect 4479 10217 4488 10251
rect 4436 10208 4488 10217
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 10784 10208 10836 10260
rect 8208 10140 8260 10192
rect 11520 10140 11572 10192
rect 11704 10183 11756 10192
rect 11704 10149 11713 10183
rect 11713 10149 11747 10183
rect 11747 10149 11756 10183
rect 11704 10140 11756 10149
rect 11888 10140 11940 10192
rect 2872 10115 2924 10124
rect 2872 10081 2881 10115
rect 2881 10081 2915 10115
rect 2915 10081 2924 10115
rect 2872 10072 2924 10081
rect 5080 10115 5132 10124
rect 2136 10004 2188 10056
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 3976 10004 4028 10056
rect 4160 10004 4212 10056
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 6920 10004 6972 10056
rect 7472 10004 7524 10056
rect 8944 10004 8996 10056
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 3424 9868 3476 9920
rect 4068 9868 4120 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 4896 9664 4948 9716
rect 5080 9664 5132 9716
rect 6092 9707 6144 9716
rect 6092 9673 6101 9707
rect 6101 9673 6135 9707
rect 6135 9673 6144 9707
rect 6092 9664 6144 9673
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 8668 9707 8720 9716
rect 8668 9673 8677 9707
rect 8677 9673 8711 9707
rect 8711 9673 8720 9707
rect 8668 9664 8720 9673
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 2872 9596 2924 9648
rect 3976 9639 4028 9648
rect 3976 9605 3985 9639
rect 3985 9605 4019 9639
rect 4019 9605 4028 9639
rect 3976 9596 4028 9605
rect 8760 9596 8812 9648
rect 9588 9664 9640 9716
rect 11520 9664 11572 9716
rect 12624 9707 12676 9716
rect 12624 9673 12633 9707
rect 12633 9673 12667 9707
rect 12667 9673 12676 9707
rect 12624 9664 12676 9673
rect 9680 9639 9732 9648
rect 9680 9605 9689 9639
rect 9689 9605 9723 9639
rect 9723 9605 9732 9639
rect 9680 9596 9732 9605
rect 11244 9639 11296 9648
rect 11244 9605 11253 9639
rect 11253 9605 11287 9639
rect 11287 9605 11296 9639
rect 11244 9596 11296 9605
rect 3056 9528 3108 9580
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 6920 9528 6972 9580
rect 8024 9528 8076 9580
rect 9312 9528 9364 9580
rect 9496 9460 9548 9512
rect 4896 9392 4948 9444
rect 2228 9324 2280 9376
rect 6460 9324 6512 9376
rect 9128 9392 9180 9444
rect 9404 9392 9456 9444
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 4252 9120 4304 9172
rect 5172 9120 5224 9172
rect 6000 9120 6052 9172
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 2412 9095 2464 9104
rect 2412 9061 2421 9095
rect 2421 9061 2455 9095
rect 2455 9061 2464 9095
rect 2412 9052 2464 9061
rect 3332 9052 3384 9104
rect 4896 9052 4948 9104
rect 6460 9052 6512 9104
rect 8208 9052 8260 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 4528 8984 4580 9036
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 11336 9027 11388 9036
rect 11336 8993 11354 9027
rect 11354 8993 11388 9027
rect 11336 8984 11388 8993
rect 11704 8984 11756 9036
rect 2136 8916 2188 8968
rect 6552 8916 6604 8968
rect 6828 8916 6880 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8760 8916 8812 8968
rect 4528 8848 4580 8900
rect 2964 8780 3016 8832
rect 4344 8780 4396 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 8668 8780 8720 8832
rect 9128 8780 9180 8832
rect 11060 8780 11112 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2412 8576 2464 8628
rect 4436 8576 4488 8628
rect 4896 8576 4948 8628
rect 3056 8508 3108 8560
rect 5540 8576 5592 8628
rect 8208 8576 8260 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 6460 8551 6512 8560
rect 6460 8517 6469 8551
rect 6469 8517 6503 8551
rect 6503 8517 6512 8551
rect 6460 8508 6512 8517
rect 1308 8440 1360 8492
rect 1584 8440 1636 8492
rect 2964 8440 3016 8492
rect 4344 8440 4396 8492
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 6000 8440 6052 8492
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 1676 8372 1728 8424
rect 2320 8372 2372 8424
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 4252 8347 4304 8356
rect 4252 8313 4261 8347
rect 4261 8313 4295 8347
rect 4295 8313 4304 8347
rect 4252 8304 4304 8313
rect 4344 8347 4396 8356
rect 4344 8313 4353 8347
rect 4353 8313 4387 8347
rect 4387 8313 4396 8347
rect 4344 8304 4396 8313
rect 7380 8304 7432 8356
rect 8760 8347 8812 8356
rect 8760 8313 8769 8347
rect 8769 8313 8803 8347
rect 8803 8313 8812 8347
rect 8760 8304 8812 8313
rect 4160 8236 4212 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1492 8032 1544 8084
rect 2136 8032 2188 8084
rect 2780 8032 2832 8084
rect 4160 8032 4212 8084
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 7380 8032 7432 8084
rect 8300 8032 8352 8084
rect 6828 8007 6880 8016
rect 6828 7973 6837 8007
rect 6837 7973 6871 8007
rect 6871 7973 6880 8007
rect 6828 7964 6880 7973
rect 3516 7896 3568 7948
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 7472 7896 7524 7948
rect 8392 7896 8444 7948
rect 6184 7828 6236 7880
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 3516 7488 3568 7540
rect 3608 7531 3660 7540
rect 3608 7497 3617 7531
rect 3617 7497 3651 7531
rect 3651 7497 3660 7531
rect 3884 7531 3936 7540
rect 3608 7488 3660 7497
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 8392 7488 8444 7540
rect 2044 7420 2096 7472
rect 4068 7420 4120 7472
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 2688 7327 2740 7336
rect 2688 7293 2697 7327
rect 2697 7293 2731 7327
rect 2731 7293 2740 7327
rect 2688 7284 2740 7293
rect 3608 7284 3660 7336
rect 4804 7327 4856 7336
rect 4804 7293 4848 7327
rect 4848 7293 4856 7327
rect 4804 7284 4856 7293
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 7380 6944 7432 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 2412 6808 2464 6860
rect 3332 6808 3384 6860
rect 4068 6672 4120 6724
rect 7564 6604 7616 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1676 6400 1728 6452
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2596 6400 2648 6452
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 3332 6400 3384 6409
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 1768 6196 1820 6248
rect 7564 6196 7616 6248
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 2412 6171 2464 6180
rect 2412 6137 2421 6171
rect 2421 6137 2455 6171
rect 2455 6137 2464 6171
rect 2412 6128 2464 6137
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1860 5856 1912 5908
rect 2596 5856 2648 5908
rect 1492 5763 1544 5772
rect 1492 5729 1510 5763
rect 1510 5729 1544 5763
rect 1492 5720 1544 5729
rect 2504 5763 2556 5772
rect 2504 5729 2522 5763
rect 2522 5729 2556 5763
rect 2504 5720 2556 5729
rect 7564 5720 7616 5772
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1492 5312 1544 5364
rect 2504 5312 2556 5364
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 1952 5176 2004 5228
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 1400 5151 1452 5160
rect 1400 5117 1444 5151
rect 1444 5117 1452 5151
rect 1400 5108 1452 5117
rect 8024 5108 8076 5160
rect 8392 5108 8444 5160
rect 7564 5015 7616 5024
rect 7564 4981 7573 5015
rect 7573 4981 7607 5015
rect 7607 4981 7616 5015
rect 7564 4972 7616 4981
rect 8760 4972 8812 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1584 4768 1636 4820
rect 1400 4675 1452 4684
rect 1400 4641 1444 4675
rect 1444 4641 1452 4675
rect 1400 4632 1452 4641
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1400 4224 1452 4276
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2320 3680 2372 3732
rect 1400 3587 1452 3596
rect 1400 3553 1444 3587
rect 1444 3553 1452 3587
rect 1400 3544 1452 3553
rect 17960 3476 18012 3528
rect 19248 3476 19300 3528
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1584 3136 1636 3188
rect 1400 3068 1452 3120
rect 1492 2975 1544 2984
rect 1492 2941 1510 2975
rect 1510 2941 1544 2975
rect 1492 2932 1544 2941
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2592 1636 2644
rect 1400 2499 1452 2508
rect 1400 2465 1444 2499
rect 1444 2465 1452 2499
rect 1400 2456 1452 2465
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 2688 2320 2740 2372
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 478 27520 534 28000
rect 1490 27520 1546 28000
rect 2502 27520 2558 28000
rect 3514 27520 3570 28000
rect 4618 27520 4674 28000
rect 5630 27520 5686 28000
rect 6642 27520 6698 28000
rect 7654 27520 7710 28000
rect 8758 27520 8814 28000
rect 9770 27520 9826 28000
rect 10782 27520 10838 28000
rect 11794 27520 11850 28000
rect 12898 27520 12954 28000
rect 13910 27520 13966 28000
rect 14922 27520 14978 28000
rect 15934 27520 15990 28000
rect 17038 27520 17094 28000
rect 18050 27520 18106 28000
rect 19062 27520 19118 28000
rect 20074 27520 20130 28000
rect 21178 27520 21234 28000
rect 22190 27520 22246 28000
rect 23202 27520 23258 28000
rect 24214 27520 24270 28000
rect 25318 27520 25374 28000
rect 26330 27520 26386 28000
rect 27342 27520 27398 28000
rect 492 21593 520 27520
rect 1398 24304 1454 24313
rect 1398 24239 1454 24248
rect 1412 23662 1440 24239
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1504 23497 1532 27520
rect 1490 23488 1546 23497
rect 1490 23423 1546 23432
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 2044 23180 2096 23186
rect 1412 22574 1440 23151
rect 2044 23122 2096 23128
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1398 22264 1454 22273
rect 1398 22199 1454 22208
rect 478 21584 534 21593
rect 478 21519 534 21528
rect 1412 21486 1440 22199
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1596 21185 1624 22918
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1412 21010 1440 21111
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 20602 1440 20946
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1400 20596 1452 20602
rect 1400 20538 1452 20544
rect 1596 17814 1624 20878
rect 1688 19242 1716 22918
rect 2056 22438 2084 23122
rect 2044 22432 2096 22438
rect 2044 22374 2096 22380
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 1952 21616 2004 21622
rect 1952 21558 2004 21564
rect 1872 19378 1900 19417
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1676 19236 1728 19242
rect 1676 19178 1728 19184
rect 1768 19236 1820 19242
rect 1768 19178 1820 19184
rect 1780 18970 1808 19178
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1584 17808 1636 17814
rect 1584 17750 1636 17756
rect 1596 16794 1624 17750
rect 1780 17218 1808 18702
rect 1872 18290 1900 19314
rect 1964 19258 1992 21558
rect 2056 19961 2084 22374
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2042 19952 2098 19961
rect 2042 19887 2098 19896
rect 1964 19230 2084 19258
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1964 18970 1992 19110
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1950 18320 2006 18329
rect 1860 18284 1912 18290
rect 1950 18255 2006 18264
rect 1860 18226 1912 18232
rect 1964 18154 1992 18255
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1858 18048 1914 18057
rect 1858 17983 1914 17992
rect 1872 17814 1900 17983
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1872 17338 1900 17750
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1780 17190 1900 17218
rect 2056 17202 2084 19230
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1780 15366 1808 15914
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 15162 1808 15302
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13802 1716 14350
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1596 13190 1624 13738
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11626 1532 12038
rect 1674 11792 1730 11801
rect 1674 11727 1730 11736
rect 1492 11620 1544 11626
rect 1492 11562 1544 11568
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 11082 1440 11494
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1308 10532 1360 10538
rect 1308 10474 1360 10480
rect 1320 8498 1348 10474
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1412 6866 1440 11018
rect 1504 8090 1532 11562
rect 1582 10840 1638 10849
rect 1582 10775 1638 10784
rect 1596 9654 1624 10775
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1688 9194 1716 11727
rect 1766 9752 1822 9761
rect 1766 9687 1822 9696
rect 1596 9166 1716 9194
rect 1596 8634 1624 9166
rect 1674 9072 1730 9081
rect 1674 9007 1676 9016
rect 1728 9007 1730 9016
rect 1676 8978 1728 8984
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1490 7712 1546 7721
rect 1490 7647 1546 7656
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1504 5778 1532 7647
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1398 5672 1454 5681
rect 1398 5607 1454 5616
rect 1412 5166 1440 5607
rect 1504 5370 1532 5714
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1596 4826 1624 8434
rect 1688 8430 1716 8978
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1780 6746 1808 9687
rect 1688 6718 1808 6746
rect 1688 6458 1716 6718
rect 1766 6624 1822 6633
rect 1766 6559 1822 6568
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 6254 1808 6559
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1872 5914 1900 17190
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16726 2084 17138
rect 2044 16720 2096 16726
rect 2148 16697 2176 21830
rect 2332 21350 2360 22034
rect 2320 21344 2372 21350
rect 2318 21312 2320 21321
rect 2372 21312 2374 21321
rect 2318 21247 2374 21256
rect 2320 20392 2372 20398
rect 2226 20360 2282 20369
rect 2320 20334 2372 20340
rect 2226 20295 2228 20304
rect 2280 20295 2282 20304
rect 2228 20266 2280 20272
rect 2332 20097 2360 20334
rect 2318 20088 2374 20097
rect 2318 20023 2374 20032
rect 2320 19780 2372 19786
rect 2320 19722 2372 19728
rect 2332 19378 2360 19722
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2424 18578 2452 22374
rect 2516 21486 2544 27520
rect 2778 27432 2834 27441
rect 2778 27367 2834 27376
rect 2686 23624 2742 23633
rect 2686 23559 2688 23568
rect 2740 23559 2742 23568
rect 2688 23530 2740 23536
rect 2792 23186 2820 27367
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 3330 23488 3386 23497
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 22778 2820 23122
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2686 22536 2742 22545
rect 2686 22471 2688 22480
rect 2740 22471 2742 22480
rect 2688 22442 2740 22448
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2686 21448 2742 21457
rect 2686 21383 2688 21392
rect 2740 21383 2742 21392
rect 2688 21354 2740 21360
rect 2504 20800 2556 20806
rect 2504 20742 2556 20748
rect 2516 19825 2544 20742
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2700 20346 2728 20402
rect 2700 20318 2820 20346
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2502 19816 2558 19825
rect 2502 19751 2558 19760
rect 2608 19310 2636 19926
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2700 18986 2728 20198
rect 2792 19145 2820 20318
rect 2884 20058 2912 22578
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3068 21350 3096 22034
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2870 19952 2926 19961
rect 2870 19887 2926 19896
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2516 18958 2728 18986
rect 2516 18601 2544 18958
rect 2688 18896 2740 18902
rect 2688 18838 2740 18844
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2332 18550 2452 18578
rect 2502 18592 2558 18601
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 2044 16662 2096 16668
rect 2134 16688 2190 16697
rect 2240 16658 2268 17002
rect 2134 16623 2190 16632
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2240 16250 2268 16594
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1964 15366 1992 16050
rect 2332 15638 2360 18550
rect 2502 18527 2558 18536
rect 2410 18456 2466 18465
rect 2410 18391 2466 18400
rect 2424 18358 2452 18391
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2424 17814 2452 18294
rect 2412 17808 2464 17814
rect 2412 17750 2464 17756
rect 2608 17202 2636 18634
rect 2700 18086 2728 18838
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16726 2636 17138
rect 2700 16794 2728 18022
rect 2792 17882 2820 18226
rect 2884 18193 2912 19887
rect 2870 18184 2926 18193
rect 2870 18119 2926 18128
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15858 2728 15914
rect 3068 15858 3096 21286
rect 2700 15830 3096 15858
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 13530 1992 15302
rect 2608 14958 2636 15574
rect 2792 15026 2820 15830
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2596 14952 2648 14958
rect 2594 14920 2596 14929
rect 2648 14920 2650 14929
rect 2228 14884 2280 14890
rect 2976 14890 3004 15438
rect 2594 14855 2650 14864
rect 2964 14884 3016 14890
rect 2228 14826 2280 14832
rect 2240 13938 2268 14826
rect 2608 14482 2636 14855
rect 2964 14826 3016 14832
rect 3160 14618 3188 23462
rect 3330 23423 3386 23432
rect 3344 22574 3372 23423
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3528 22438 3556 27520
rect 4066 26344 4122 26353
rect 4066 26279 4068 26288
rect 4120 26279 4122 26288
rect 4068 26250 4120 26256
rect 4066 25392 4122 25401
rect 4066 25327 4068 25336
rect 4120 25327 4122 25336
rect 4068 25298 4120 25304
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 4172 23798 4200 24210
rect 4632 23866 4660 27520
rect 5644 25242 5672 27520
rect 6552 26308 6604 26314
rect 6552 26250 6604 26256
rect 5552 25214 5672 25242
rect 5552 24290 5580 25214
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5460 24274 5580 24290
rect 6564 24274 6592 26250
rect 5448 24268 5580 24274
rect 5500 24262 5580 24268
rect 6552 24268 6604 24274
rect 5448 24210 5500 24216
rect 6552 24210 6604 24216
rect 5262 24168 5318 24177
rect 5262 24103 5318 24112
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3422 21584 3478 21593
rect 3422 21519 3478 21528
rect 3436 21486 3464 21519
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3436 18290 3464 20198
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3804 19145 3832 19246
rect 3790 19136 3846 19145
rect 3790 19071 3846 19080
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 3436 17882 3464 18226
rect 3516 18148 3568 18154
rect 3516 18090 3568 18096
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3528 17338 3556 18090
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3252 16114 3280 16662
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3344 15978 3372 17070
rect 3804 16182 3832 18226
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3988 15570 4016 21830
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4160 21412 4212 21418
rect 4160 21354 4212 21360
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 18290 4108 21247
rect 4172 20058 4200 21354
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4356 18465 4384 21422
rect 4526 21176 4582 21185
rect 4526 21111 4582 21120
rect 4540 18766 4568 21111
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4632 18902 4660 20742
rect 4724 20602 4752 20946
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4724 20074 4752 20538
rect 4724 20046 4844 20074
rect 4816 19990 4844 20046
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4816 19514 4844 19926
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4816 19174 4844 19450
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4342 18456 4398 18465
rect 4342 18391 4398 18400
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4540 17882 4568 18702
rect 4632 18426 4660 18838
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4724 17814 4752 19110
rect 4908 18306 4936 24006
rect 5276 23866 5304 24103
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6564 23866 6592 24210
rect 6656 24177 6684 27520
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 6642 24168 6698 24177
rect 6642 24103 6698 24112
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 4988 19304 5040 19310
rect 4986 19272 4988 19281
rect 5040 19272 5042 19281
rect 4986 19207 5042 19216
rect 5092 18698 5120 19926
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 4816 18278 4936 18306
rect 4712 17808 4764 17814
rect 4712 17750 4764 17756
rect 4066 17232 4122 17241
rect 4066 17167 4122 17176
rect 4080 17134 4108 17167
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4250 17096 4306 17105
rect 4250 17031 4306 17040
rect 4264 16794 4292 17031
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4066 16688 4122 16697
rect 4066 16623 4068 16632
rect 4120 16623 4122 16632
rect 4068 16594 4120 16600
rect 4080 15706 4108 16594
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16250 4384 16526
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4250 16008 4306 16017
rect 4250 15943 4306 15952
rect 4264 15706 4292 15943
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3252 14890 3280 15030
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3252 14793 3280 14826
rect 3238 14784 3294 14793
rect 3238 14719 3294 14728
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2608 14074 2636 14418
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 3160 13938 3188 14554
rect 3252 14482 3280 14719
rect 3988 14618 4016 15506
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3606 13968 3662 13977
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3424 13932 3476 13938
rect 3606 13903 3662 13912
rect 3424 13874 3476 13880
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3252 13705 3280 13738
rect 3238 13696 3294 13705
rect 3238 13631 3294 13640
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2516 12866 2544 13126
rect 2608 12986 2636 13398
rect 3436 13326 3464 13874
rect 3514 13696 3570 13705
rect 3514 13631 3570 13640
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2884 12918 2912 13262
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 2872 12912 2924 12918
rect 2516 12838 2636 12866
rect 2872 12854 2924 12860
rect 3068 12850 3096 13194
rect 2320 12708 2372 12714
rect 2240 12668 2320 12696
rect 2240 12102 2268 12668
rect 2320 12650 2372 12656
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1964 5234 1992 12038
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2134 11384 2190 11393
rect 2134 11319 2190 11328
rect 2148 11286 2176 11319
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 2056 7478 2084 10474
rect 2148 10266 2176 11222
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2148 10146 2176 10202
rect 2424 10146 2452 11698
rect 2516 11558 2544 12242
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11257 2544 11494
rect 2502 11248 2558 11257
rect 2502 11183 2558 11192
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2516 10742 2544 11086
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2148 10118 2360 10146
rect 2424 10118 2544 10146
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 8974 2176 9998
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8090 2176 8910
rect 2240 8265 2268 9318
rect 2332 8514 2360 10118
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2424 9110 2452 9998
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2424 8634 2452 9046
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2332 8486 2452 8514
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2226 8256 2282 8265
rect 2226 8191 2282 8200
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 6458 2084 6802
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1766 4720 1822 4729
rect 1400 4684 1452 4690
rect 1766 4655 1822 4664
rect 1400 4626 1452 4632
rect 1412 4593 1440 4626
rect 1398 4584 1454 4593
rect 1398 4519 1454 4528
rect 1412 4282 1440 4519
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 3505 1440 3538
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 1412 3126 1440 3431
rect 1596 3194 1624 3431
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1398 2544 1454 2553
rect 1398 2479 1400 2488
rect 1452 2479 1454 2488
rect 1400 2450 1452 2456
rect 1504 1465 1532 2926
rect 1582 2680 1638 2689
rect 1582 2615 1584 2624
rect 1636 2615 1638 2624
rect 1584 2586 1636 2592
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 1780 480 1808 4655
rect 2332 3738 2360 8366
rect 2424 6866 2452 8486
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2410 6216 2466 6225
rect 2410 6151 2412 6160
rect 2464 6151 2466 6160
rect 2412 6122 2464 6128
rect 2516 5778 2544 10118
rect 2608 6458 2636 12838
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2688 12708 2740 12714
rect 2740 12668 2820 12696
rect 2688 12650 2740 12656
rect 2686 12608 2742 12617
rect 2686 12543 2742 12552
rect 2700 11762 2728 12543
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2700 11150 2728 11562
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 9761 2728 11086
rect 2686 9752 2742 9761
rect 2686 9687 2742 9696
rect 2792 8090 2820 12668
rect 3068 12617 3096 12786
rect 3054 12608 3110 12617
rect 3054 12543 3110 12552
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2884 11898 2912 12242
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 3054 11792 3110 11801
rect 3054 11727 3056 11736
rect 3108 11727 3110 11736
rect 3056 11698 3108 11704
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11082 3004 11494
rect 3068 11354 3096 11698
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3160 11218 3188 12174
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 9654 2912 10066
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2976 9330 3004 11018
rect 3344 10810 3372 11698
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3436 9926 3464 10542
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 2884 9302 3004 9330
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 7970 2912 9302
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8498 3004 8774
rect 3068 8566 3096 9522
rect 3344 9110 3372 9522
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2700 7942 2912 7970
rect 2700 7342 2728 7942
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 3344 6866 3372 9046
rect 3528 7954 3556 13631
rect 3620 10810 3648 13903
rect 4080 12714 4108 14214
rect 4172 14074 4200 14418
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4172 12986 4200 14010
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3792 12436 3844 12442
rect 3896 12424 3924 12650
rect 3844 12396 3924 12424
rect 3792 12378 3844 12384
rect 3896 12306 3924 12396
rect 4356 12306 4384 16186
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4172 11558 4200 12242
rect 4632 11762 4660 12378
rect 4816 11801 4844 18278
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4908 18057 4936 18090
rect 4894 18048 4950 18057
rect 4894 17983 4950 17992
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4908 17202 4936 17614
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4908 16794 4936 17138
rect 5000 16998 5028 17750
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5000 16674 5028 16934
rect 4908 16658 5028 16674
rect 4896 16652 5028 16658
rect 4948 16646 5028 16652
rect 4896 16594 4948 16600
rect 4908 15162 4936 16594
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4908 14890 4936 15098
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4908 14006 4936 14826
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4908 13802 4936 13942
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4908 13462 4936 13738
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4908 12986 4936 13398
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4802 11792 4858 11801
rect 4620 11756 4672 11762
rect 4802 11727 4858 11736
rect 4620 11698 4672 11704
rect 4908 11626 4936 12922
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 4172 10062 4200 11494
rect 4908 11286 4936 11562
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4908 10810 4936 11222
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3988 9654 4016 9998
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3882 8800 3938 8809
rect 3882 8735 3938 8744
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3528 7546 3556 7890
rect 3606 7576 3662 7585
rect 3516 7540 3568 7546
rect 3896 7546 3924 8735
rect 3606 7511 3608 7520
rect 3516 7482 3568 7488
rect 3660 7511 3662 7520
rect 3884 7540 3936 7546
rect 3608 7482 3660 7488
rect 3884 7482 3936 7488
rect 3620 7342 3648 7482
rect 4080 7478 4108 9862
rect 4448 9586 4476 10202
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4264 8362 4292 9114
rect 4540 9058 4568 10406
rect 4802 9752 4858 9761
rect 4908 9722 4936 10746
rect 4802 9687 4858 9696
rect 4896 9716 4948 9722
rect 4448 9042 4568 9058
rect 4448 9036 4580 9042
rect 4448 9030 4528 9036
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8498 4384 8774
rect 4448 8634 4476 9030
rect 4528 8978 4580 8984
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4540 8498 4568 8842
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4356 8362 4384 8434
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 8090 4200 8230
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4356 7954 4384 8298
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4356 7546 4384 7890
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4816 7342 4844 9687
rect 4896 9658 4948 9664
rect 4908 9450 4936 9658
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4908 9110 4936 9386
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4908 8634 4936 9046
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 7585 5028 15098
rect 5092 14278 5120 15302
rect 5276 14770 5304 23530
rect 6840 23338 6868 24006
rect 6840 23310 6960 23338
rect 6932 23254 6960 23310
rect 6920 23248 6972 23254
rect 5630 23216 5686 23225
rect 6920 23190 6972 23196
rect 5630 23151 5632 23160
rect 5684 23151 5686 23160
rect 5632 23122 5684 23128
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5354 17912 5410 17921
rect 5354 17847 5410 17856
rect 5368 16658 5396 17847
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 16114 5396 16594
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5368 15706 5396 16050
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5460 15162 5488 21286
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 5920 19990 5948 20266
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 18834 6040 21286
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5552 18222 5580 18566
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18216 5592 18222
rect 5538 18184 5540 18193
rect 5592 18184 5594 18193
rect 5538 18119 5594 18128
rect 6012 18086 6040 18770
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5552 17241 5580 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5538 17232 5594 17241
rect 5538 17167 5594 17176
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 16182 5580 17070
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5552 15042 5580 15642
rect 5644 15502 5672 15982
rect 6104 15688 6132 22918
rect 6552 22092 6604 22098
rect 6552 22034 6604 22040
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 18834 6224 21830
rect 6564 21690 6592 22034
rect 6918 21992 6974 22001
rect 6918 21927 6974 21936
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6460 21072 6512 21078
rect 6460 21014 6512 21020
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6380 20058 6408 20878
rect 6472 20262 6500 21014
rect 6460 20256 6512 20262
rect 6458 20224 6460 20233
rect 6512 20224 6514 20233
rect 6458 20159 6514 20168
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6288 19514 6316 19790
rect 6564 19786 6592 21626
rect 6932 21554 6960 21927
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6564 19657 6592 19722
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6380 19281 6408 19654
rect 6366 19272 6422 19281
rect 6366 19207 6422 19216
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6012 15660 6132 15688
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5460 15026 5580 15042
rect 5448 15020 5580 15026
rect 5500 15014 5580 15020
rect 5448 14962 5500 14968
rect 5908 14952 5960 14958
rect 5906 14920 5908 14929
rect 5960 14920 5962 14929
rect 5906 14855 5962 14864
rect 5184 14742 5304 14770
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 11801 5120 14214
rect 5078 11792 5134 11801
rect 5078 11727 5134 11736
rect 5092 11257 5120 11727
rect 5078 11248 5134 11257
rect 5078 11183 5134 11192
rect 5092 10742 5120 11183
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10130 5120 10542
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9722 5120 10066
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5184 9178 5212 14742
rect 5262 14648 5318 14657
rect 5262 14583 5264 14592
rect 5316 14583 5318 14592
rect 5264 14554 5316 14560
rect 5538 14512 5594 14521
rect 5538 14447 5594 14456
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12646 5304 13262
rect 5552 12986 5580 14447
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5722 13696 5778 13705
rect 5722 13631 5778 13640
rect 5736 13530 5764 13631
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5276 12345 5304 12582
rect 5262 12336 5318 12345
rect 5262 12271 5318 12280
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4986 7576 5042 7585
rect 4986 7511 5042 7520
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4066 6896 4122 6905
rect 3332 6860 3384 6866
rect 4066 6831 4122 6840
rect 3332 6802 3384 6808
rect 3344 6458 3372 6802
rect 4080 6730 4108 6831
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 5368 5953 5396 12718
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11393 5580 11494
rect 5538 11384 5594 11393
rect 5538 11319 5594 11328
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10810 5580 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9178 6040 15660
rect 6196 15570 6224 18566
rect 6380 18154 6408 19207
rect 6748 18970 6776 19994
rect 6840 19854 6868 20198
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 18970 6868 19246
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 16726 6960 18022
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6380 15910 6408 16594
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6104 15162 6132 15506
rect 6380 15502 6408 15846
rect 6368 15496 6420 15502
rect 6656 15473 6684 16594
rect 7024 15978 7052 24550
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7564 23180 7616 23186
rect 7668 23168 7696 27520
rect 8772 24818 8800 27520
rect 9784 25362 9812 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9232 24954 9260 25298
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 8850 24848 8906 24857
rect 8760 24812 8812 24818
rect 8850 24783 8906 24792
rect 8760 24754 8812 24760
rect 8864 24614 8892 24783
rect 8300 24608 8352 24614
rect 8220 24556 8300 24562
rect 8220 24550 8352 24556
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8220 24534 8340 24550
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 8024 24064 8076 24070
rect 8024 24006 8076 24012
rect 7746 23896 7802 23905
rect 7746 23831 7748 23840
rect 7800 23831 7802 23840
rect 7748 23802 7800 23808
rect 8036 23254 8064 24006
rect 8128 23662 8156 24210
rect 8116 23656 8168 23662
rect 8116 23598 8168 23604
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 7616 23140 7696 23168
rect 7564 23122 7616 23128
rect 7116 22778 7144 23122
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7760 22234 7788 23190
rect 8036 22778 8064 23190
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7484 20806 7512 22034
rect 8220 21962 8248 24534
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8864 23798 8892 24006
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8312 22234 8340 22374
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8024 21344 8076 21350
rect 8220 21321 8248 21422
rect 8404 21350 8432 23530
rect 8496 23497 8524 23598
rect 8576 23520 8628 23526
rect 8482 23488 8538 23497
rect 8576 23462 8628 23468
rect 8482 23423 8538 23432
rect 8392 21344 8444 21350
rect 8024 21286 8076 21292
rect 8206 21312 8262 21321
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 19990 7512 20742
rect 8036 20466 8064 21286
rect 8392 21286 8444 21292
rect 8206 21247 8262 21256
rect 8116 21072 8168 21078
rect 8116 21014 8168 21020
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8128 20330 8156 21014
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 7746 20224 7802 20233
rect 7746 20159 7802 20168
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7760 19310 7788 20159
rect 8128 20058 8156 20266
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 8128 19242 8156 19994
rect 8220 19242 8248 20742
rect 8496 20602 8524 23423
rect 8588 22098 8616 23462
rect 8864 23254 8892 23734
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8680 22642 8708 22918
rect 9140 22710 9168 23666
rect 9692 23322 9720 25094
rect 9784 24954 9812 25298
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9864 24744 9916 24750
rect 9864 24686 9916 24692
rect 10046 24712 10102 24721
rect 9772 24268 9824 24274
rect 9772 24210 9824 24216
rect 9784 23866 9812 24210
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9876 23610 9904 24686
rect 10046 24647 10102 24656
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9784 23582 9904 23610
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9692 22710 9720 23258
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8588 21690 8616 22034
rect 9140 21690 9168 22646
rect 9784 22642 9812 23582
rect 9864 23520 9916 23526
rect 9862 23488 9864 23497
rect 9916 23488 9918 23497
rect 9862 23423 9918 23432
rect 9968 23254 9996 24006
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 9968 22778 9996 23190
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 10060 21962 10088 24647
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10152 23594 10364 23610
rect 10152 23588 10376 23594
rect 10152 23582 10324 23588
rect 10152 23526 10180 23582
rect 10324 23530 10376 23536
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 22420 10732 25094
rect 10796 24857 10824 27520
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 10782 24848 10838 24857
rect 10782 24783 10838 24792
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10782 24168 10838 24177
rect 10782 24103 10838 24112
rect 10796 23526 10824 24103
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10796 23322 10824 23462
rect 10784 23316 10836 23322
rect 10784 23258 10836 23264
rect 10876 23044 10928 23050
rect 10876 22986 10928 22992
rect 10888 22642 10916 22986
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10704 22392 10824 22420
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10796 22114 10824 22392
rect 10704 22086 10824 22114
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 8588 21146 8616 21626
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8772 20058 8800 21422
rect 10060 21321 10088 21422
rect 10046 21312 10102 21321
rect 10046 21247 10102 21256
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 8404 19174 8432 19858
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8392 19168 8444 19174
rect 8298 19136 8354 19145
rect 8392 19110 8444 19116
rect 8298 19071 8354 19080
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 7392 18426 7420 18770
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 8036 18222 8064 18770
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 7760 17882 7788 18158
rect 8312 17882 8340 19071
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7564 17672 7616 17678
rect 7562 17640 7564 17649
rect 7616 17640 7618 17649
rect 7562 17575 7618 17584
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17202 7144 17478
rect 7576 17338 7604 17575
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7484 16130 7512 16594
rect 7300 16102 7512 16130
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7300 15910 7328 16102
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6736 15496 6788 15502
rect 6368 15438 6420 15444
rect 6642 15464 6698 15473
rect 6736 15438 6788 15444
rect 6642 15399 6698 15408
rect 6656 15162 6684 15399
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6642 14784 6698 14793
rect 6642 14719 6698 14728
rect 6656 14618 6684 14719
rect 6748 14657 6776 15438
rect 6734 14648 6790 14657
rect 6644 14612 6696 14618
rect 6734 14583 6790 14592
rect 6644 14554 6696 14560
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6104 14006 6132 14486
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6196 13530 6224 14418
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6472 13433 6500 13806
rect 6458 13424 6514 13433
rect 6458 13359 6514 13368
rect 6458 12880 6514 12889
rect 6458 12815 6514 12824
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6104 11937 6132 12242
rect 6090 11928 6146 11937
rect 6090 11863 6092 11872
rect 6144 11863 6146 11872
rect 6092 11834 6144 11840
rect 6288 11558 6316 12242
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11257 6316 11494
rect 6472 11354 6500 12815
rect 6748 12442 6776 14583
rect 6932 14498 6960 15642
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7024 14958 7052 15302
rect 7012 14952 7064 14958
rect 7064 14900 7144 14906
rect 7012 14894 7144 14900
rect 7024 14878 7144 14894
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6840 14482 6960 14498
rect 6828 14476 6960 14482
rect 6880 14470 6960 14476
rect 6828 14418 6880 14424
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6840 13818 6868 13942
rect 6840 13790 6960 13818
rect 6932 12986 6960 13790
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6932 12714 6960 12922
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11626 6776 12038
rect 6918 11792 6974 11801
rect 6918 11727 6974 11736
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6274 11248 6330 11257
rect 6274 11183 6330 11192
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6104 9722 6132 10066
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6196 9602 6224 11018
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10130 6592 10406
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9761 6592 10066
rect 6550 9752 6606 9761
rect 6550 9687 6552 9696
rect 6604 9687 6606 9696
rect 6552 9658 6604 9664
rect 6104 9574 6224 9602
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5552 8634 5580 9007
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5630 8528 5686 8537
rect 6012 8498 6040 9114
rect 5630 8463 5686 8472
rect 6000 8492 6052 8498
rect 5644 8430 5672 8463
rect 6000 8434 6052 8440
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6104 6905 6132 9574
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 9110 6500 9318
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6472 8566 6500 9046
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6564 8090 6592 8910
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6196 7206 6224 7822
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 2594 5944 2650 5953
rect 2594 5879 2596 5888
rect 2648 5879 2650 5888
rect 5354 5944 5410 5953
rect 5354 5879 5410 5888
rect 2596 5850 2648 5856
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2516 5370 2544 5714
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5262 4040 5318 4049
rect 5262 3975 5318 3984
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2686 2408 2742 2417
rect 2686 2343 2688 2352
rect 2740 2343 2742 2352
rect 2688 2314 2740 2320
rect 2884 513 2912 2450
rect 2870 504 2926 513
rect 1766 0 1822 480
rect 5276 480 5304 3975
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6196 2689 6224 7142
rect 6748 3505 6776 11562
rect 6932 11354 6960 11727
rect 7024 11626 7052 14758
rect 7116 13462 7144 14878
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7116 12986 7144 13398
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7116 12442 7144 12922
rect 7208 12850 7236 13670
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6932 10606 6960 11290
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9586 6960 9998
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7024 9058 7052 10406
rect 6840 9030 7052 9058
rect 6840 8974 6868 9030
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6840 7410 6868 7958
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 7300 4049 7328 15846
rect 7392 13326 7420 15914
rect 7576 15910 7604 17138
rect 7944 17066 7972 17750
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7746 16688 7802 16697
rect 8404 16658 8432 19110
rect 8588 18970 8616 19246
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8482 18184 8538 18193
rect 8482 18119 8538 18128
rect 8496 17338 8524 18119
rect 8680 17785 8708 19654
rect 8772 19310 8800 19994
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8772 18426 8800 19246
rect 9784 18970 9812 20334
rect 9968 20058 9996 20878
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 19514 9996 19858
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 10060 18834 10088 21247
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10612 20618 10640 21014
rect 10704 20924 10732 22086
rect 10784 22024 10836 22030
rect 10782 21992 10784 22001
rect 10836 21992 10838 22001
rect 10782 21927 10838 21936
rect 10796 21078 10824 21927
rect 10888 21146 10916 22442
rect 10980 22114 11008 24550
rect 11440 24342 11468 25094
rect 11624 24682 11652 25298
rect 11612 24676 11664 24682
rect 11612 24618 11664 24624
rect 11428 24336 11480 24342
rect 11428 24278 11480 24284
rect 11440 23866 11468 24278
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11072 23254 11100 23802
rect 11624 23662 11652 24142
rect 11808 23905 11836 27520
rect 12912 25498 12940 27520
rect 13924 25498 13952 27520
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 12624 25356 12676 25362
rect 12624 25298 12676 25304
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 12636 24750 12664 25298
rect 12624 24744 12676 24750
rect 12622 24712 12624 24721
rect 12676 24712 12678 24721
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12440 24676 12492 24682
rect 12622 24647 12678 24656
rect 12440 24618 12492 24624
rect 12636 24621 12664 24647
rect 11794 23896 11850 23905
rect 11794 23831 11850 23840
rect 12176 23730 12204 24618
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 24342 12296 24550
rect 12256 24336 12308 24342
rect 12256 24278 12308 24284
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 11612 23656 11664 23662
rect 11610 23624 11612 23633
rect 11664 23624 11666 23633
rect 11610 23559 11666 23568
rect 12176 23526 12204 23666
rect 12268 23526 12296 24278
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 11060 23248 11112 23254
rect 11060 23190 11112 23196
rect 11796 23248 11848 23254
rect 11796 23190 11848 23196
rect 11072 23066 11100 23190
rect 11336 23112 11388 23118
rect 11072 23038 11192 23066
rect 11336 23054 11388 23060
rect 11060 22160 11112 22166
rect 10980 22108 11060 22114
rect 10980 22102 11112 22108
rect 10980 22086 11100 22102
rect 10980 21690 11008 22086
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11164 21570 11192 23038
rect 11348 22234 11376 23054
rect 11808 22778 11836 23190
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11612 22500 11664 22506
rect 11612 22442 11664 22448
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11624 22166 11652 22442
rect 11886 22264 11942 22273
rect 11886 22199 11888 22208
rect 11940 22199 11942 22208
rect 11888 22170 11940 22176
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11624 21962 11652 22102
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 10980 21542 11192 21570
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10704 20896 10824 20924
rect 10612 20590 10732 20618
rect 10704 20330 10732 20590
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 19174 10180 19858
rect 10704 19242 10732 20266
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18834 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8864 18086 8892 18226
rect 9048 18154 9076 18634
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18358 9260 18566
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8666 17776 8722 17785
rect 8666 17711 8722 17720
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 7746 16623 7748 16632
rect 7800 16623 7802 16632
rect 8392 16652 8444 16658
rect 7748 16594 7800 16600
rect 8392 16594 8444 16600
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7668 14482 7696 16050
rect 7852 16046 7880 16458
rect 8680 16114 8708 17711
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 8668 15972 8720 15978
rect 8772 15960 8800 16390
rect 8864 16114 8892 18022
rect 9048 17921 9076 18090
rect 9034 17912 9090 17921
rect 9034 17847 9090 17856
rect 9140 17542 9168 18158
rect 9508 17882 9536 18770
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 10060 18086 10088 18294
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 9588 18080 9640 18086
rect 10048 18080 10100 18086
rect 9640 18028 9720 18034
rect 9588 18022 9720 18028
rect 10048 18022 10100 18028
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9600 18006 9720 18022
rect 9692 17882 9720 18006
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9862 17640 9918 17649
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17066 9168 17478
rect 9310 17232 9366 17241
rect 9310 17167 9366 17176
rect 9324 17134 9352 17167
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9324 16794 9352 17070
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9416 16522 9444 17070
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16590 9628 17002
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16250 9444 16458
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9600 16182 9628 16526
rect 9692 16250 9720 16594
rect 9784 16590 9812 17614
rect 9862 17575 9918 17584
rect 9876 17202 9904 17575
rect 10060 17542 10088 18022
rect 10152 17678 10180 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17882 10732 18090
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 17338 10088 17478
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8720 15932 8800 15960
rect 8668 15914 8720 15920
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8206 15600 8262 15609
rect 8036 15337 8064 15574
rect 8206 15535 8208 15544
rect 8260 15535 8262 15544
rect 8208 15506 8260 15512
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8022 15328 8078 15337
rect 8022 15263 8078 15272
rect 8036 15162 8064 15263
rect 8024 15156 8076 15162
rect 8220 15144 8248 15370
rect 8300 15156 8352 15162
rect 8220 15116 8300 15144
rect 8024 15098 8076 15104
rect 8300 15098 8352 15104
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 14074 7696 14418
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7562 13968 7618 13977
rect 7562 13903 7618 13912
rect 7576 13870 7604 13903
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13530 7604 13806
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7392 12850 7420 13262
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11354 7420 12174
rect 7576 11762 7604 13262
rect 7760 12238 7788 14554
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8220 14074 8248 14418
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8220 13870 8248 14010
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8680 13802 8708 15914
rect 9140 15434 9168 16118
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9232 15366 9260 15914
rect 9876 15609 9904 16730
rect 9968 16697 9996 17070
rect 9954 16688 10010 16697
rect 9954 16623 10010 16632
rect 10060 16454 10088 17274
rect 10152 16998 10180 17614
rect 10704 17338 10732 17682
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10152 16114 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10520 16046 10548 16390
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10704 15978 10732 16390
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9862 15600 9918 15609
rect 9862 15535 9918 15544
rect 9956 15564 10008 15570
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8680 13190 8708 13738
rect 8772 13297 8800 14758
rect 9126 14376 9182 14385
rect 9232 14362 9260 15302
rect 9678 15056 9734 15065
rect 9678 14991 9734 15000
rect 9692 14550 9720 14991
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9692 14362 9720 14486
rect 9182 14334 9260 14362
rect 9600 14334 9720 14362
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9126 14311 9128 14320
rect 9180 14311 9182 14320
rect 9128 14282 9180 14288
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 14006 8984 14214
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 9140 13870 9168 14282
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 8758 13288 8814 13297
rect 8758 13223 8814 13232
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8404 12986 8432 13126
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8680 12753 8708 13126
rect 8666 12744 8722 12753
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 8300 12708 8352 12714
rect 8666 12679 8722 12688
rect 8300 12650 8352 12656
rect 7944 12374 7972 12650
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7944 11898 7972 12310
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7576 10266 7604 11086
rect 7944 10470 7972 11222
rect 8208 11144 8260 11150
rect 8312 11132 8340 12650
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11626 8616 12038
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8260 11104 8340 11132
rect 8208 11086 8260 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10606 8340 10950
rect 8300 10600 8352 10606
rect 8220 10548 8300 10554
rect 8220 10542 8352 10548
rect 8220 10526 8340 10542
rect 7932 10464 7984 10470
rect 8220 10418 8248 10526
rect 7932 10406 7984 10412
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7944 10169 7972 10406
rect 8128 10390 8248 10418
rect 7930 10160 7986 10169
rect 7930 10095 7986 10104
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8362 7420 8774
rect 7484 8498 7512 9998
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9178 8064 9522
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7392 8090 7420 8298
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7342 7420 8026
rect 7484 7954 7512 8434
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 7002 7420 7278
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 6254 7604 6598
rect 8128 6322 8156 10390
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9382 8248 10134
rect 8208 9376 8260 9382
rect 8206 9344 8208 9353
rect 8260 9344 8262 9353
rect 8206 9279 8262 9288
rect 8220 9110 8248 9279
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8634 8248 8910
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8298 8256 8354 8265
rect 8298 8191 8354 8200
rect 8312 8090 8340 8191
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 7954 8432 11222
rect 8680 11014 8708 12679
rect 8772 12186 8800 13223
rect 9140 12442 9168 13806
rect 9600 13734 9628 14334
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9588 13728 9640 13734
rect 9508 13676 9588 13682
rect 9508 13670 9640 13676
rect 9508 13654 9628 13670
rect 9508 13274 9536 13654
rect 9692 13546 9720 13874
rect 9600 13530 9720 13546
rect 9588 13524 9720 13530
rect 9640 13518 9720 13524
rect 9588 13466 9640 13472
rect 9784 13410 9812 14350
rect 9600 13394 9812 13410
rect 9588 13388 9812 13394
rect 9640 13382 9812 13388
rect 9588 13330 9640 13336
rect 9680 13320 9732 13326
rect 9416 13268 9680 13274
rect 9416 13262 9732 13268
rect 9416 13246 9720 13262
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 8772 12158 8984 12186
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11762 8892 12038
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8772 11286 8800 11562
rect 8956 11506 8984 12158
rect 8864 11478 8984 11506
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8680 9722 8708 10746
rect 8760 10736 8812 10742
rect 8864 10724 8892 11478
rect 9140 11354 9168 12378
rect 9310 11656 9366 11665
rect 9310 11591 9366 11600
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9140 10810 9168 11290
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9324 10742 9352 11591
rect 8812 10696 8892 10724
rect 9312 10736 9364 10742
rect 8760 10678 8812 10684
rect 9312 10678 9364 10684
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8772 9654 8800 10678
rect 9324 10266 9352 10678
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8404 7546 8432 7890
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 7576 5778 7604 6190
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 5030 7604 5714
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5370 8064 5510
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8036 5166 8064 5306
rect 8404 5166 8432 6190
rect 8680 5234 8708 8774
rect 8772 8362 8800 8910
rect 8956 8537 8984 9998
rect 9324 9586 9352 10202
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9416 9450 9444 13246
rect 9692 12986 9720 13246
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9784 12889 9812 13382
rect 9876 13161 9904 15535
rect 9956 15506 10008 15512
rect 9968 15065 9996 15506
rect 10060 15502 10088 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15638 10732 15914
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9954 15056 10010 15065
rect 9954 14991 10010 15000
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9968 14482 9996 14826
rect 10060 14822 10088 15438
rect 10704 15337 10732 15574
rect 10690 15328 10746 15337
rect 10690 15263 10746 15272
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14521 10088 14758
rect 10046 14512 10102 14521
rect 9956 14476 10008 14482
rect 10046 14447 10102 14456
rect 9956 14418 10008 14424
rect 9968 14006 9996 14418
rect 10152 14414 10180 14826
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13190 9996 13670
rect 9956 13184 10008 13190
rect 9862 13152 9918 13161
rect 9956 13126 10008 13132
rect 9862 13087 9918 13096
rect 9770 12880 9826 12889
rect 9770 12815 9826 12824
rect 9968 12442 9996 13126
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 10060 11937 10088 14214
rect 10230 13968 10286 13977
rect 10336 13938 10364 14282
rect 10230 13903 10286 13912
rect 10324 13932 10376 13938
rect 10244 13870 10272 13903
rect 10324 13874 10376 13880
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 12238 10180 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12918 10364 13262
rect 10704 13258 10732 13806
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10612 12782 10640 13126
rect 10704 12782 10732 13194
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10046 11928 10102 11937
rect 10428 11898 10456 12174
rect 10046 11863 10102 11872
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10704 11694 10732 12582
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 9518 9536 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10796 11150 10824 20896
rect 10980 20602 11008 21542
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11440 20806 11468 21422
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11532 21185 11560 21354
rect 11518 21176 11574 21185
rect 11518 21111 11574 21120
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19378 11192 19654
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11348 18834 11376 19994
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 10888 17762 10916 18770
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11072 18358 11100 18566
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10888 17734 11008 17762
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10888 16454 10916 17274
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10980 16250 11008 17734
rect 11072 16572 11100 18294
rect 11256 18290 11284 18566
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11348 17882 11376 18770
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11244 17808 11296 17814
rect 11244 17750 11296 17756
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17338 11192 17478
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11164 17241 11192 17274
rect 11150 17232 11206 17241
rect 11150 17167 11206 17176
rect 11256 16726 11284 17750
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11072 16544 11376 16572
rect 11348 16454 11376 16544
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15366 11100 16050
rect 11256 15978 11284 16390
rect 11348 16182 11376 16390
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10968 14952 11020 14958
rect 10966 14920 10968 14929
rect 11020 14920 11022 14929
rect 10966 14855 11022 14864
rect 10874 14376 10930 14385
rect 10874 14311 10930 14320
rect 10888 13394 10916 14311
rect 10980 14074 11008 14855
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10980 13326 11008 14010
rect 11072 13802 11100 15302
rect 11164 14278 11192 15438
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11164 13326 11192 14214
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11334 13968 11390 13977
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11256 12918 11284 13942
rect 11334 13903 11390 13912
rect 11348 13530 11376 13903
rect 11440 13530 11468 20742
rect 11900 20602 11928 20946
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 12084 19990 12112 21626
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11716 18902 11744 19178
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11716 18154 11744 18838
rect 11808 18290 11836 19858
rect 12084 19514 12112 19926
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12176 19310 12204 23462
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12268 18970 12296 23462
rect 12360 21146 12388 24074
rect 12452 22778 12480 24618
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12544 23633 12572 24006
rect 12912 23730 12940 24142
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12530 23624 12586 23633
rect 12636 23594 12664 23666
rect 12530 23559 12532 23568
rect 12584 23559 12586 23568
rect 12624 23588 12676 23594
rect 12532 23530 12584 23536
rect 12624 23530 12676 23536
rect 12912 23322 12940 23666
rect 12900 23316 12952 23322
rect 12900 23258 12952 23264
rect 12530 23216 12586 23225
rect 12530 23151 12532 23160
rect 12584 23151 12586 23160
rect 12532 23122 12584 23128
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12452 22438 12480 22714
rect 12544 22642 12572 23122
rect 13188 22642 13216 24142
rect 13648 23848 13676 24550
rect 13832 24138 13860 25298
rect 14936 25242 14964 27520
rect 14844 25214 14964 25242
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 14292 24721 14320 25094
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14278 24712 14334 24721
rect 14278 24647 14280 24656
rect 14332 24647 14334 24656
rect 14280 24618 14332 24624
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13820 23860 13872 23866
rect 13648 23820 13820 23848
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12452 21690 12480 22034
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12636 21570 12664 22578
rect 13556 22545 13584 23054
rect 13542 22536 13598 22545
rect 13542 22471 13598 22480
rect 13556 22234 13584 22471
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 13004 21690 13032 22034
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12452 21542 12664 21570
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12452 21026 12480 21542
rect 12820 21486 12848 21558
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 12360 21010 12480 21026
rect 12348 21004 12480 21010
rect 12400 20998 12480 21004
rect 12348 20946 12400 20952
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12440 19712 12492 19718
rect 12636 19700 12664 21354
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 21010 12756 21286
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12728 20058 12756 20946
rect 12820 20806 12848 21422
rect 13648 21146 13676 23820
rect 13820 23802 13872 23808
rect 14384 23254 14412 24754
rect 14554 24440 14610 24449
rect 14554 24375 14556 24384
rect 14608 24375 14610 24384
rect 14556 24346 14608 24352
rect 14568 23730 14596 24346
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14660 23594 14688 24142
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 14462 23488 14518 23497
rect 14462 23423 14518 23432
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 13740 22778 13768 23190
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 14384 22642 14412 23190
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13726 21176 13782 21185
rect 13636 21140 13688 21146
rect 13726 21111 13782 21120
rect 13636 21082 13688 21088
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12492 19672 12664 19700
rect 12440 19654 12492 19660
rect 12360 18970 12388 19654
rect 12452 19292 12480 19654
rect 12532 19304 12584 19310
rect 12452 19264 12532 19292
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12452 18850 12480 19264
rect 12532 19246 12584 19252
rect 12360 18822 12480 18850
rect 12820 18834 12848 20742
rect 13280 20262 13308 21014
rect 13740 20466 13768 21111
rect 13832 20602 13860 22102
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13542 20360 13598 20369
rect 13542 20295 13598 20304
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13096 19961 13124 20198
rect 13082 19952 13138 19961
rect 13082 19887 13138 19896
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19310 13032 19790
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12808 18828 12860 18834
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 12162 18184 12218 18193
rect 11704 18148 11756 18154
rect 12162 18119 12218 18128
rect 11704 18090 11756 18096
rect 12176 17882 12204 18119
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 11886 17776 11942 17785
rect 11886 17711 11888 17720
rect 11940 17711 11942 17720
rect 11888 17682 11940 17688
rect 11900 17338 11928 17682
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 15502 11560 16526
rect 11624 15910 11652 16662
rect 11808 16590 11836 16934
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11624 13394 11652 15846
rect 11716 15570 11744 15982
rect 12176 15910 12204 16594
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11532 12986 11560 13126
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11624 12442 11652 13330
rect 11716 12986 11744 15506
rect 12084 15473 12112 15506
rect 12070 15464 12126 15473
rect 12070 15399 12126 15408
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11808 14822 11836 15302
rect 12084 15162 12112 15399
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 14618 11836 14758
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11808 13190 11836 14554
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 13870 11928 14350
rect 11992 14074 12020 14418
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12176 14006 12204 15846
rect 12360 15638 12388 18822
rect 12808 18770 12860 18776
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13096 18426 13124 18770
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13188 18290 13216 18770
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17882 12480 18022
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12452 15570 12480 17274
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 15144 12480 15506
rect 12268 15116 12480 15144
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11808 12782 11836 13126
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10980 11626 11008 12310
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 11164 11286 11192 12038
rect 11900 11898 11928 13806
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12442 12020 13262
rect 12268 13258 12296 15116
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 13462 12480 14282
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12452 12986 12480 13398
rect 12544 13002 12572 18158
rect 13188 17882 13216 18226
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17134 12940 17478
rect 13188 17134 13216 17682
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 17202 13308 17614
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12912 16046 12940 17070
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13096 16046 13124 16730
rect 13188 16658 13216 17070
rect 13266 16688 13322 16697
rect 13176 16652 13228 16658
rect 13556 16658 13584 20295
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 19990 13676 20198
rect 13924 20058 13952 22374
rect 14384 22234 14412 22578
rect 14476 22506 14504 23423
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 14752 22098 14780 24754
rect 14844 24614 14872 25214
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14844 22642 14872 23666
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15212 23338 15240 23530
rect 15396 23526 15424 24210
rect 15474 23760 15530 23769
rect 15474 23695 15530 23704
rect 15384 23520 15436 23526
rect 15382 23488 15384 23497
rect 15436 23488 15438 23497
rect 15382 23423 15438 23432
rect 15120 23322 15240 23338
rect 15108 23316 15240 23322
rect 15160 23310 15240 23316
rect 15108 23258 15160 23264
rect 15292 23248 15344 23254
rect 15292 23190 15344 23196
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14200 21690 14228 22034
rect 14844 21690 14872 22578
rect 15304 22438 15332 23190
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21690 15332 22374
rect 15488 22098 15516 23695
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15396 21622 15424 21898
rect 15580 21894 15608 22986
rect 15660 22500 15712 22506
rect 15660 22442 15712 22448
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14002 21176 14058 21185
rect 14002 21111 14004 21120
rect 14056 21111 14058 21120
rect 14004 21082 14056 21088
rect 14660 20534 14688 21422
rect 15396 21146 15424 21558
rect 15580 21457 15608 21830
rect 15672 21486 15700 22442
rect 15660 21480 15712 21486
rect 15566 21448 15622 21457
rect 15660 21422 15712 21428
rect 15566 21383 15622 21392
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20602 15332 20878
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13648 19174 13676 19926
rect 14370 19816 14426 19825
rect 14370 19751 14372 19760
rect 14424 19751 14426 19760
rect 14372 19722 14424 19728
rect 14384 19446 14412 19722
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14554 19272 14610 19281
rect 14554 19207 14556 19216
rect 14608 19207 14610 19216
rect 14556 19178 14608 19184
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13648 18086 13676 19110
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18222 13952 18566
rect 14844 18426 14872 20266
rect 15488 20262 15516 21014
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15474 19952 15530 19961
rect 15474 19887 15530 19896
rect 15488 19854 15516 19887
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15488 19446 15516 19790
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15580 19378 15608 20402
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15672 19514 15700 19926
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 15200 18352 15252 18358
rect 15198 18320 15200 18329
rect 15252 18320 15254 18329
rect 15304 18306 15332 18702
rect 15580 18358 15608 19314
rect 15764 18970 15792 25094
rect 15948 24410 15976 27520
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16316 24954 16344 25298
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16316 24857 16344 24890
rect 16302 24848 16358 24857
rect 16302 24783 16358 24792
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16868 24449 16896 24550
rect 16854 24440 16910 24449
rect 15936 24404 15988 24410
rect 16854 24375 16910 24384
rect 15936 24346 15988 24352
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16486 23760 16542 23769
rect 16486 23695 16542 23704
rect 16500 23508 16528 23695
rect 16592 23526 16620 24210
rect 16580 23520 16632 23526
rect 16210 23488 16266 23497
rect 16500 23480 16580 23508
rect 16580 23462 16632 23468
rect 16210 23423 16266 23432
rect 16224 22642 16252 23423
rect 17052 23322 17080 27520
rect 17958 24168 18014 24177
rect 17958 24103 17960 24112
rect 18012 24103 18014 24112
rect 17960 24074 18012 24080
rect 18064 23610 18092 27520
rect 18234 24304 18290 24313
rect 18234 24239 18236 24248
rect 18288 24239 18290 24248
rect 18236 24210 18288 24216
rect 18248 23866 18276 24210
rect 18970 24168 19026 24177
rect 18970 24103 19026 24112
rect 18984 23866 19012 24103
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18984 23662 19012 23802
rect 17880 23582 18092 23610
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 16316 22642 16344 23054
rect 17236 22778 17264 23054
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16118 22400 16174 22409
rect 16118 22335 16174 22344
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16040 21690 16068 21966
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 16132 20534 16160 22335
rect 16224 22234 16252 22578
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16316 21554 16344 22578
rect 16488 22160 16540 22166
rect 16394 22128 16450 22137
rect 16488 22102 16540 22108
rect 16394 22063 16450 22072
rect 16408 22030 16436 22063
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16500 21690 16528 22102
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16684 21622 16712 21966
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16592 21146 16620 21286
rect 17880 21146 17908 23582
rect 17960 23520 18012 23526
rect 17958 23488 17960 23497
rect 18012 23488 18014 23497
rect 17958 23423 18014 23432
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18524 22438 18552 23122
rect 18052 22432 18104 22438
rect 18512 22432 18564 22438
rect 18052 22374 18104 22380
rect 18510 22400 18512 22409
rect 18564 22400 18566 22409
rect 18064 22137 18092 22374
rect 18510 22335 18566 22344
rect 18050 22128 18106 22137
rect 18050 22063 18106 22072
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 18248 21690 18276 22034
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18248 21350 18276 21626
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17420 20602 17448 20946
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16132 19854 16160 20470
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19242 16620 19654
rect 17144 19242 17172 19722
rect 17328 19514 17356 19926
rect 18156 19854 18184 20334
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18800 19922 18828 20266
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 16580 19236 16632 19242
rect 17132 19236 17184 19242
rect 16580 19178 16632 19184
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15254 18278 15332 18306
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15764 18290 15792 18906
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16040 18290 16068 18838
rect 15752 18284 15804 18290
rect 15198 18255 15254 18264
rect 15752 18226 15804 18232
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16592 18222 16620 19178
rect 16960 19174 16988 19205
rect 17132 19178 17184 19184
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 16948 19168 17000 19174
rect 16946 19136 16948 19145
rect 17000 19136 17002 19145
rect 16946 19071 17002 19080
rect 16960 18970 16988 19071
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 17144 18902 17172 19178
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 13912 18216 13964 18222
rect 13910 18184 13912 18193
rect 16580 18216 16632 18222
rect 13964 18184 13966 18193
rect 16580 18158 16632 18164
rect 13910 18119 13966 18128
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13648 17814 13676 18022
rect 15120 17882 15148 18090
rect 16592 18034 16620 18158
rect 17236 18154 17264 19178
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 16500 18006 16620 18034
rect 16500 17882 16528 18006
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 13648 17338 13676 17750
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13266 16623 13322 16632
rect 13544 16652 13596 16658
rect 13176 16594 13228 16600
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12636 14482 12664 15914
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12728 14822 12756 15438
rect 12912 15366 12940 15982
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 14958 12940 15302
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12716 14816 12768 14822
rect 12714 14784 12716 14793
rect 12768 14784 12770 14793
rect 12714 14719 12770 14728
rect 12728 14618 12756 14719
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 13530 12664 14418
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 13802 12848 14350
rect 12912 13977 12940 14894
rect 13188 14618 13216 16594
rect 13280 16114 13308 16623
rect 13544 16594 13596 16600
rect 13832 16130 13860 16662
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13740 16102 13860 16130
rect 13636 15904 13688 15910
rect 13634 15872 13636 15881
rect 13740 15892 13768 16102
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13688 15872 13768 15892
rect 13690 15864 13768 15872
rect 13634 15807 13690 15816
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13464 14958 13492 15506
rect 13832 15366 13860 15982
rect 13924 15434 13952 16934
rect 14660 16794 14688 17070
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 15488 16726 15516 17614
rect 15672 16998 15700 17750
rect 17328 17746 17356 19450
rect 18052 19304 18104 19310
rect 18050 19272 18052 19281
rect 18104 19272 18106 19281
rect 18050 19207 18106 19216
rect 18156 18902 18184 19790
rect 18800 19514 18828 19858
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 17500 18896 17552 18902
rect 17500 18838 17552 18844
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 17512 18086 17540 18838
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17880 18426 17908 18702
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17882 17540 18022
rect 18156 17882 18184 18158
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 17328 17338 17356 17682
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15476 16720 15528 16726
rect 15474 16688 15476 16697
rect 15528 16688 15530 16697
rect 15474 16623 15530 16632
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14200 15706 14228 16526
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15672 15978 15700 16934
rect 15856 16794 15884 17070
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15108 15904 15160 15910
rect 15382 15872 15438 15881
rect 15160 15852 15332 15858
rect 15108 15846 15332 15852
rect 15120 15830 15332 15846
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13820 15360 13872 15366
rect 13740 15308 13820 15314
rect 13740 15302 13872 15308
rect 13740 15286 13860 15302
rect 13740 15026 13768 15286
rect 13924 15162 13952 15370
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 15304 15026 15332 15830
rect 15382 15807 15438 15816
rect 15396 15162 15424 15807
rect 15672 15638 15700 15914
rect 15764 15910 15792 16662
rect 17696 16590 17724 17206
rect 18156 17134 18184 17478
rect 18708 17270 18736 17682
rect 19076 17338 19104 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20088 24313 20116 27520
rect 20074 24304 20130 24313
rect 20074 24239 20130 24248
rect 21192 23866 21220 27520
rect 21270 24712 21326 24721
rect 21270 24647 21326 24656
rect 21284 23866 21312 24647
rect 21914 23896 21970 23905
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21272 23860 21324 23866
rect 21914 23831 21916 23840
rect 21272 23802 21324 23808
rect 21968 23831 21970 23840
rect 21916 23802 21968 23808
rect 21928 23662 21956 23802
rect 22008 23792 22060 23798
rect 22204 23746 22232 27520
rect 23216 23905 23244 27520
rect 24228 24177 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 25332 24857 25360 27520
rect 25318 24848 25374 24857
rect 25318 24783 25374 24792
rect 25502 24304 25558 24313
rect 25136 24268 25188 24274
rect 25502 24239 25558 24248
rect 25136 24210 25188 24216
rect 24214 24168 24270 24177
rect 24214 24103 24270 24112
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23202 23896 23258 23905
rect 23202 23831 23258 23840
rect 22060 23740 22232 23746
rect 22008 23734 22232 23740
rect 22020 23718 22232 23734
rect 21916 23656 21968 23662
rect 19522 23624 19578 23633
rect 21916 23598 21968 23604
rect 19522 23559 19578 23568
rect 19536 23526 19564 23559
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 19352 22273 19380 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19338 22264 19394 22273
rect 19622 22256 19918 22276
rect 19338 22199 19394 22208
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 17960 16720 18012 16726
rect 23492 16697 23520 23462
rect 23584 19281 23612 24006
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 25148 23798 25176 24210
rect 25516 23866 25544 24239
rect 26344 23882 26372 27520
rect 27356 24313 27384 27520
rect 27342 24304 27398 24313
rect 27342 24239 27398 24248
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 26160 23854 26372 23882
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25516 23662 25544 23802
rect 26160 23798 26188 23854
rect 26148 23792 26200 23798
rect 26148 23734 26200 23740
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 23570 19272 23626 19281
rect 23570 19207 23626 19216
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 17960 16662 18012 16668
rect 18602 16688 18658 16697
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15764 15570 15792 15846
rect 16592 15638 16620 15914
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15842 15328 15898 15337
rect 15842 15263 15898 15272
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 14002 14920 14058 14929
rect 14002 14855 14058 14864
rect 15658 14920 15714 14929
rect 15658 14855 15714 14864
rect 14016 14618 14044 14855
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13084 14000 13136 14006
rect 12898 13968 12954 13977
rect 13084 13942 13136 13948
rect 12898 13903 12954 13912
rect 13096 13870 13124 13942
rect 13084 13864 13136 13870
rect 13082 13832 13084 13841
rect 13136 13832 13138 13841
rect 12808 13796 12860 13802
rect 13082 13767 13138 13776
rect 12808 13738 12860 13744
rect 13832 13734 13860 14010
rect 14016 13938 14044 14554
rect 15384 14476 15436 14482
rect 15436 14436 15516 14464
rect 15384 14418 15436 14424
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15396 13977 15424 14282
rect 15382 13968 15438 13977
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14464 13932 14516 13938
rect 15488 13938 15516 14436
rect 15382 13903 15384 13912
rect 14464 13874 14516 13880
rect 15436 13903 15438 13912
rect 15476 13932 15528 13938
rect 15384 13874 15436 13880
rect 15476 13874 15528 13880
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13188 13433 13216 13466
rect 13174 13424 13230 13433
rect 13084 13388 13136 13394
rect 13174 13359 13230 13368
rect 13636 13388 13688 13394
rect 13084 13330 13136 13336
rect 13636 13330 13688 13336
rect 13096 13161 13124 13330
rect 13082 13152 13138 13161
rect 13082 13087 13138 13096
rect 12440 12980 12492 12986
rect 12544 12974 12756 13002
rect 13648 12986 13676 13330
rect 13832 13297 13860 13670
rect 14016 13530 14044 13738
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13818 13288 13874 13297
rect 13874 13246 13952 13274
rect 13818 13223 13874 13232
rect 13818 13152 13874 13161
rect 13818 13087 13874 13096
rect 12440 12922 12492 12928
rect 12452 12594 12480 12922
rect 12728 12753 12756 12974
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 12806 12880 12862 12889
rect 12806 12815 12808 12824
rect 12860 12815 12862 12824
rect 12808 12786 12860 12792
rect 12714 12744 12770 12753
rect 12714 12679 12716 12688
rect 12768 12679 12770 12688
rect 12716 12650 12768 12656
rect 12728 12619 12756 12650
rect 12452 12566 12572 12594
rect 12544 12442 12572 12566
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11992 11830 12020 12378
rect 12452 12345 12480 12378
rect 12438 12336 12494 12345
rect 12164 12300 12216 12306
rect 12438 12271 12494 12280
rect 12164 12242 12216 12248
rect 12176 11898 12204 12242
rect 12820 11898 12848 12786
rect 13096 12306 13124 12922
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13188 12374 13216 12854
rect 13832 12442 13860 13087
rect 13924 12782 13952 13246
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13096 11898 13124 12242
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 11980 11824 12032 11830
rect 12176 11801 12204 11834
rect 11980 11766 12032 11772
rect 12162 11792 12218 11801
rect 11244 11688 11296 11694
rect 11992 11665 12020 11766
rect 12162 11727 12218 11736
rect 12820 11694 12848 11834
rect 12808 11688 12860 11694
rect 11244 11630 11296 11636
rect 11978 11656 12034 11665
rect 11256 11354 11284 11630
rect 12808 11630 12860 11636
rect 11978 11591 12034 11600
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 10266 9996 10610
rect 10152 10538 10180 10950
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9678 9752 9734 9761
rect 9588 9716 9640 9722
rect 9678 9687 9734 9696
rect 9588 9658 9640 9664
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9140 8838 9168 9386
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8942 8528 8998 8537
rect 8942 8463 8944 8472
rect 8996 8463 8998 8472
rect 8944 8434 8996 8440
rect 8956 8403 8984 8434
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 9600 5545 9628 9658
rect 9692 9654 9720 9687
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9770 9344 9826 9353
rect 9770 9279 9826 9288
rect 9784 9042 9812 9279
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8634 9812 8978
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9586 5536 9642 5545
rect 9586 5471 9642 5480
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 7576 4729 7604 4966
rect 7562 4720 7618 4729
rect 7562 4655 7618 4664
rect 7286 4040 7342 4049
rect 7286 3975 7342 3984
rect 6734 3496 6790 3505
rect 6734 3431 6790 3440
rect 6182 2680 6238 2689
rect 6182 2615 6238 2624
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 8772 480 8800 4966
rect 10152 2417 10180 10474
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10796 10266 10824 11086
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10606 11100 10950
rect 11164 10606 11192 11222
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 11072 10062 11100 10542
rect 11532 10198 11560 11494
rect 11888 11280 11940 11286
rect 14476 11257 14504 13874
rect 15488 13841 15516 13874
rect 15568 13864 15620 13870
rect 15474 13832 15530 13841
rect 15568 13806 15620 13812
rect 15474 13767 15530 13776
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 11888 11222 11940 11228
rect 14462 11248 14518 11257
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10198 11744 10950
rect 11900 10470 11928 11222
rect 14462 11183 14518 11192
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11992 10674 12020 11086
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12820 10606 12848 10950
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11900 10198 11928 10406
rect 11520 10192 11572 10198
rect 11242 10160 11298 10169
rect 11520 10134 11572 10140
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11242 10095 11298 10104
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 11072 9178 11100 9998
rect 11256 9654 11284 10095
rect 11532 9722 11560 10134
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11716 9042 11744 10134
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12636 9722 12664 10066
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 11072 6225 11100 8774
rect 11348 8634 11376 8978
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 11058 6216 11114 6225
rect 11058 6151 11114 6160
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 12254 5536 12310 5545
rect 12254 5471 12310 5480
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10138 2408 10194 2417
rect 10138 2343 10194 2352
rect 12268 480 12296 5471
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15488 3369 15516 13767
rect 15580 13462 15608 13806
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15672 3482 15700 14855
rect 15856 14550 15884 15263
rect 16132 14618 16160 15438
rect 16500 14822 16528 15574
rect 16684 15502 16712 16526
rect 17052 16182 17080 16526
rect 17972 16266 18000 16662
rect 23478 16688 23534 16697
rect 18602 16623 18658 16632
rect 19340 16652 19392 16658
rect 18616 16590 18644 16623
rect 23478 16623 23534 16632
rect 19340 16594 19392 16600
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 17880 16250 18000 16266
rect 18616 16250 18644 16526
rect 19352 16250 19380 16594
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 17868 16244 18000 16250
rect 17920 16238 18000 16244
rect 18604 16244 18656 16250
rect 17868 16186 17920 16192
rect 18604 16186 18656 16192
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 17512 15162 17540 15506
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17880 15094 17908 16186
rect 19352 15337 19380 16186
rect 19536 15473 19564 16390
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19522 15464 19578 15473
rect 19522 15399 19578 15408
rect 19338 15328 19394 15337
rect 19338 15263 19394 15272
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 17868 15088 17920 15094
rect 16670 15056 16726 15065
rect 17868 15030 17920 15036
rect 16670 14991 16726 15000
rect 16684 14958 16712 14991
rect 16672 14952 16724 14958
rect 16578 14920 16634 14929
rect 16672 14894 16724 14900
rect 16578 14855 16634 14864
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15750 14376 15806 14385
rect 15750 14311 15806 14320
rect 15764 14074 15792 14311
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 16500 11626 16528 14758
rect 16592 14482 16620 14855
rect 16856 14816 16908 14822
rect 16854 14784 16856 14793
rect 16908 14784 16910 14793
rect 16854 14719 16910 14728
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16868 14521 16896 14554
rect 16854 14512 16910 14521
rect 16580 14476 16632 14482
rect 16854 14447 16910 14456
rect 16580 14418 16632 14424
rect 16592 14074 16620 14418
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 17958 13968 18014 13977
rect 17958 13903 18014 13912
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 3505 16528 11562
rect 17972 3534 18000 13903
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 17960 3528 18012 3534
rect 16486 3496 16542 3505
rect 15672 3454 15792 3482
rect 15474 3360 15530 3369
rect 14956 3292 15252 3312
rect 15474 3295 15530 3304
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15764 480 15792 3454
rect 17960 3470 18012 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 26238 3496 26294 3505
rect 16486 3431 16542 3440
rect 19260 480 19288 3470
rect 26238 3431 26294 3440
rect 22742 3360 22798 3369
rect 22742 3295 22798 3304
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 22756 480 22784 3295
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 26252 480 26280 3431
rect 2870 439 2926 448
rect 5262 0 5318 480
rect 8758 0 8814 480
rect 12254 0 12310 480
rect 15750 0 15806 480
rect 19246 0 19302 480
rect 22742 0 22798 480
rect 26238 0 26294 480
<< via2 >>
rect 1398 24248 1454 24304
rect 1490 23432 1546 23488
rect 1398 23160 1454 23216
rect 1398 22208 1454 22264
rect 478 21528 534 21584
rect 1398 21120 1454 21176
rect 1582 21120 1638 21176
rect 2042 19896 2098 19952
rect 1950 18264 2006 18320
rect 1858 17992 1914 18048
rect 1674 11736 1730 11792
rect 1582 10784 1638 10840
rect 1766 9696 1822 9752
rect 1674 9036 1730 9072
rect 1674 9016 1676 9036
rect 1676 9016 1728 9036
rect 1728 9016 1730 9036
rect 1490 7656 1546 7712
rect 1398 5616 1454 5672
rect 1766 6568 1822 6624
rect 2318 21292 2320 21312
rect 2320 21292 2372 21312
rect 2372 21292 2374 21312
rect 2318 21256 2374 21292
rect 2226 20324 2282 20360
rect 2226 20304 2228 20324
rect 2228 20304 2280 20324
rect 2280 20304 2282 20324
rect 2318 20032 2374 20088
rect 2778 27376 2834 27432
rect 2686 23588 2742 23624
rect 2686 23568 2688 23588
rect 2688 23568 2740 23588
rect 2740 23568 2742 23588
rect 2686 22500 2742 22536
rect 2686 22480 2688 22500
rect 2688 22480 2740 22500
rect 2740 22480 2742 22500
rect 2686 21412 2742 21448
rect 2686 21392 2688 21412
rect 2688 21392 2740 21412
rect 2740 21392 2742 21412
rect 2502 19760 2558 19816
rect 2870 19896 2926 19952
rect 2778 19080 2834 19136
rect 2134 16632 2190 16688
rect 2502 18536 2558 18592
rect 2410 18400 2466 18456
rect 2870 18128 2926 18184
rect 2594 14900 2596 14920
rect 2596 14900 2648 14920
rect 2648 14900 2650 14920
rect 2594 14864 2650 14900
rect 3330 23432 3386 23488
rect 4066 26308 4122 26344
rect 4066 26288 4068 26308
rect 4068 26288 4120 26308
rect 4120 26288 4122 26308
rect 4066 25356 4122 25392
rect 4066 25336 4068 25356
rect 4068 25336 4120 25356
rect 4120 25336 4122 25356
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5262 24112 5318 24168
rect 3422 21528 3478 21584
rect 3790 19080 3846 19136
rect 4066 21256 4122 21312
rect 4526 21120 4582 21176
rect 4342 18400 4398 18456
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6642 24112 6698 24168
rect 4986 19252 4988 19272
rect 4988 19252 5040 19272
rect 5040 19252 5042 19272
rect 4986 19216 5042 19252
rect 4066 17176 4122 17232
rect 4250 17040 4306 17096
rect 4066 16652 4122 16688
rect 4066 16632 4068 16652
rect 4068 16632 4120 16652
rect 4120 16632 4122 16652
rect 4250 15952 4306 16008
rect 3238 14728 3294 14784
rect 3606 13912 3662 13968
rect 3238 13640 3294 13696
rect 3514 13640 3570 13696
rect 2134 11328 2190 11384
rect 2502 11192 2558 11248
rect 2226 8200 2282 8256
rect 1766 4664 1822 4720
rect 1398 4528 1454 4584
rect 1398 3440 1454 3496
rect 1582 3440 1638 3496
rect 1398 2508 1454 2544
rect 1398 2488 1400 2508
rect 1400 2488 1452 2508
rect 1452 2488 1454 2508
rect 1582 2644 1638 2680
rect 1582 2624 1584 2644
rect 1584 2624 1636 2644
rect 1636 2624 1638 2644
rect 1490 1400 1546 1456
rect 2410 6180 2466 6216
rect 2410 6160 2412 6180
rect 2412 6160 2464 6180
rect 2464 6160 2466 6180
rect 2686 12552 2742 12608
rect 2686 9696 2742 9752
rect 3054 12552 3110 12608
rect 3054 11756 3110 11792
rect 3054 11736 3056 11756
rect 3056 11736 3108 11756
rect 3108 11736 3110 11756
rect 4894 17992 4950 18048
rect 4802 11736 4858 11792
rect 3882 8744 3938 8800
rect 3606 7540 3662 7576
rect 3606 7520 3608 7540
rect 3608 7520 3660 7540
rect 3660 7520 3662 7540
rect 4802 9696 4858 9752
rect 5630 23180 5686 23216
rect 5630 23160 5632 23180
rect 5632 23160 5684 23180
rect 5684 23160 5686 23180
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5354 17856 5410 17912
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5538 18164 5540 18184
rect 5540 18164 5592 18184
rect 5592 18164 5594 18184
rect 5538 18128 5594 18164
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5538 17176 5594 17232
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6918 21936 6974 21992
rect 6458 20204 6460 20224
rect 6460 20204 6512 20224
rect 6512 20204 6514 20224
rect 6458 20168 6514 20204
rect 6366 19216 6422 19272
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5906 14900 5908 14920
rect 5908 14900 5960 14920
rect 5960 14900 5962 14920
rect 5906 14864 5962 14900
rect 5078 11736 5134 11792
rect 5078 11192 5134 11248
rect 5262 14612 5318 14648
rect 5262 14592 5264 14612
rect 5264 14592 5316 14612
rect 5316 14592 5318 14612
rect 5538 14456 5594 14512
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5722 13640 5778 13696
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5262 12280 5318 12336
rect 4986 7520 5042 7576
rect 4066 6840 4122 6896
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5538 11328 5594 11384
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 8850 24792 8906 24848
rect 7746 23860 7802 23896
rect 7746 23840 7748 23860
rect 7748 23840 7800 23860
rect 7800 23840 7802 23860
rect 8482 23432 8538 23488
rect 8206 21256 8262 21312
rect 7746 20168 7802 20224
rect 10046 24656 10102 24712
rect 9862 23468 9864 23488
rect 9864 23468 9916 23488
rect 9916 23468 9918 23488
rect 9862 23432 9918 23468
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10782 24792 10838 24848
rect 10782 24112 10838 24168
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10046 21256 10102 21312
rect 8298 19080 8354 19136
rect 7562 17620 7564 17640
rect 7564 17620 7616 17640
rect 7616 17620 7618 17640
rect 7562 17584 7618 17620
rect 6642 15408 6698 15464
rect 6642 14728 6698 14784
rect 6734 14592 6790 14648
rect 6458 13368 6514 13424
rect 6458 12824 6514 12880
rect 6090 11892 6146 11928
rect 6090 11872 6092 11892
rect 6092 11872 6144 11892
rect 6144 11872 6146 11892
rect 6918 11736 6974 11792
rect 6274 11192 6330 11248
rect 6550 9716 6606 9752
rect 6550 9696 6552 9716
rect 6552 9696 6604 9716
rect 6604 9696 6606 9716
rect 5538 9016 5594 9072
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5630 8472 5686 8528
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6090 6840 6146 6896
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 2594 5908 2650 5944
rect 2594 5888 2596 5908
rect 2596 5888 2648 5908
rect 2648 5888 2650 5908
rect 5354 5888 5410 5944
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5262 3984 5318 4040
rect 2686 2372 2742 2408
rect 2686 2352 2688 2372
rect 2688 2352 2740 2372
rect 2740 2352 2742 2372
rect 2870 448 2926 504
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 7746 16652 7802 16688
rect 8482 18128 8538 18184
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10782 21972 10784 21992
rect 10784 21972 10836 21992
rect 10836 21972 10838 21992
rect 10782 21936 10838 21972
rect 12622 24692 12624 24712
rect 12624 24692 12676 24712
rect 12676 24692 12678 24712
rect 12622 24656 12678 24692
rect 11794 23840 11850 23896
rect 11610 23604 11612 23624
rect 11612 23604 11664 23624
rect 11664 23604 11666 23624
rect 11610 23568 11666 23604
rect 11886 22228 11942 22264
rect 11886 22208 11888 22228
rect 11888 22208 11940 22228
rect 11940 22208 11942 22228
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 8666 17720 8722 17776
rect 7746 16632 7748 16652
rect 7748 16632 7800 16652
rect 7800 16632 7802 16652
rect 9034 17856 9090 17912
rect 9310 17176 9366 17232
rect 9862 17584 9918 17640
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 8206 15564 8262 15600
rect 8206 15544 8208 15564
rect 8208 15544 8260 15564
rect 8260 15544 8262 15564
rect 8022 15272 8078 15328
rect 7562 13912 7618 13968
rect 9954 16632 10010 16688
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9862 15544 9918 15600
rect 9126 14340 9182 14376
rect 9678 15000 9734 15056
rect 9126 14320 9128 14340
rect 9128 14320 9180 14340
rect 9180 14320 9182 14340
rect 8758 13232 8814 13288
rect 8666 12688 8722 12744
rect 7930 10104 7986 10160
rect 8206 9324 8208 9344
rect 8208 9324 8260 9344
rect 8260 9324 8262 9344
rect 8206 9288 8262 9324
rect 8298 8200 8354 8256
rect 9310 11600 9366 11656
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9954 15000 10010 15056
rect 10690 15272 10746 15328
rect 10046 14456 10102 14512
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9862 13096 9918 13152
rect 9770 12824 9826 12880
rect 10230 13912 10286 13968
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10046 11872 10102 11928
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11518 21120 11574 21176
rect 11150 17176 11206 17232
rect 10966 14900 10968 14920
rect 10968 14900 11020 14920
rect 11020 14900 11022 14920
rect 10966 14864 11022 14900
rect 10874 14320 10930 14376
rect 11334 13912 11390 13968
rect 12530 23588 12586 23624
rect 12530 23568 12532 23588
rect 12532 23568 12584 23588
rect 12584 23568 12586 23588
rect 12530 23180 12586 23216
rect 12530 23160 12532 23180
rect 12532 23160 12584 23180
rect 12584 23160 12586 23180
rect 14278 24676 14334 24712
rect 14278 24656 14280 24676
rect 14280 24656 14332 24676
rect 14332 24656 14334 24676
rect 13542 22480 13598 22536
rect 14554 24404 14610 24440
rect 14554 24384 14556 24404
rect 14556 24384 14608 24404
rect 14608 24384 14610 24404
rect 14462 23432 14518 23488
rect 13726 21120 13782 21176
rect 13542 20304 13598 20360
rect 13082 19896 13138 19952
rect 12162 18128 12218 18184
rect 11886 17740 11942 17776
rect 11886 17720 11888 17740
rect 11888 17720 11940 17740
rect 11940 17720 11942 17740
rect 12070 15408 12126 15464
rect 13266 16632 13322 16688
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15474 23704 15530 23760
rect 15382 23468 15384 23488
rect 15384 23468 15436 23488
rect 15436 23468 15438 23488
rect 15382 23432 15438 23468
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14002 21140 14058 21176
rect 14002 21120 14004 21140
rect 14004 21120 14056 21140
rect 14056 21120 14058 21140
rect 15566 21392 15622 21448
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14370 19780 14426 19816
rect 14370 19760 14372 19780
rect 14372 19760 14424 19780
rect 14424 19760 14426 19780
rect 14554 19236 14610 19272
rect 14554 19216 14556 19236
rect 14556 19216 14608 19236
rect 14608 19216 14610 19236
rect 15474 19896 15530 19952
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15198 18300 15200 18320
rect 15200 18300 15252 18320
rect 15252 18300 15254 18320
rect 16302 24792 16358 24848
rect 16854 24384 16910 24440
rect 16486 23704 16542 23760
rect 16210 23432 16266 23488
rect 17958 24132 18014 24168
rect 17958 24112 17960 24132
rect 17960 24112 18012 24132
rect 18012 24112 18014 24132
rect 18234 24268 18290 24304
rect 18234 24248 18236 24268
rect 18236 24248 18288 24268
rect 18288 24248 18290 24268
rect 18970 24112 19026 24168
rect 16118 22344 16174 22400
rect 16394 22072 16450 22128
rect 17958 23468 17960 23488
rect 17960 23468 18012 23488
rect 18012 23468 18014 23488
rect 17958 23432 18014 23468
rect 18510 22380 18512 22400
rect 18512 22380 18564 22400
rect 18564 22380 18566 22400
rect 18510 22344 18566 22380
rect 18050 22072 18106 22128
rect 15198 18264 15254 18300
rect 16946 19116 16948 19136
rect 16948 19116 17000 19136
rect 17000 19116 17002 19136
rect 16946 19080 17002 19116
rect 13910 18164 13912 18184
rect 13912 18164 13964 18184
rect 13964 18164 13966 18184
rect 13910 18128 13966 18164
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 12714 14764 12716 14784
rect 12716 14764 12768 14784
rect 12768 14764 12770 14784
rect 12714 14728 12770 14764
rect 13634 15852 13636 15872
rect 13636 15852 13688 15872
rect 13688 15852 13690 15872
rect 13634 15816 13690 15852
rect 18050 19252 18052 19272
rect 18052 19252 18104 19272
rect 18104 19252 18106 19272
rect 18050 19216 18106 19252
rect 15474 16668 15476 16688
rect 15476 16668 15528 16688
rect 15528 16668 15530 16688
rect 15474 16632 15530 16668
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15382 15816 15438 15872
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20074 24248 20130 24304
rect 21270 24656 21326 24712
rect 21914 23860 21970 23896
rect 21914 23840 21916 23860
rect 21916 23840 21968 23860
rect 21968 23840 21970 23860
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 25318 24792 25374 24848
rect 25502 24248 25558 24304
rect 24214 24112 24270 24168
rect 23202 23840 23258 23896
rect 19522 23568 19578 23624
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19338 22208 19394 22264
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 27342 24248 27398 24304
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 23570 19216 23626 19272
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 15842 15272 15898 15328
rect 14002 14864 14058 14920
rect 15658 14864 15714 14920
rect 12898 13912 12954 13968
rect 13082 13812 13084 13832
rect 13084 13812 13136 13832
rect 13136 13812 13138 13832
rect 13082 13776 13138 13812
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15382 13932 15438 13968
rect 15382 13912 15384 13932
rect 15384 13912 15436 13932
rect 15436 13912 15438 13932
rect 13174 13368 13230 13424
rect 13082 13096 13138 13152
rect 13818 13232 13874 13288
rect 13818 13096 13874 13152
rect 12806 12844 12862 12880
rect 12806 12824 12808 12844
rect 12808 12824 12860 12844
rect 12860 12824 12862 12844
rect 12714 12708 12770 12744
rect 12714 12688 12716 12708
rect 12716 12688 12768 12708
rect 12768 12688 12770 12708
rect 12438 12280 12494 12336
rect 12162 11736 12218 11792
rect 11978 11600 12034 11656
rect 9678 9696 9734 9752
rect 8942 8492 8998 8528
rect 8942 8472 8944 8492
rect 8944 8472 8996 8492
rect 8996 8472 8998 8492
rect 9770 9288 9826 9344
rect 9586 5480 9642 5536
rect 7562 4664 7618 4720
rect 7286 3984 7342 4040
rect 6734 3440 6790 3496
rect 6182 2624 6238 2680
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 15474 13776 15530 13832
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14462 11192 14518 11248
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 11242 10104 11298 10160
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 11058 6160 11114 6216
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 12254 5480 12310 5536
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10138 2352 10194 2408
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 18602 16632 18658 16688
rect 23478 16632 23534 16688
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19522 15408 19578 15464
rect 19338 15272 19394 15328
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 16670 15000 16726 15056
rect 16578 14864 16634 14920
rect 15750 14320 15806 14376
rect 16854 14764 16856 14784
rect 16856 14764 16908 14784
rect 16908 14764 16910 14784
rect 16854 14728 16910 14764
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 16854 14456 16910 14512
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 17958 13912 18014 13968
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 15474 3304 15530 3360
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16486 3440 16542 3496
rect 26238 3440 26294 3496
rect 22742 3304 22798 3360
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 0 27434 480 27464
rect 2773 27434 2839 27437
rect 0 27432 2839 27434
rect 0 27376 2778 27432
rect 2834 27376 2839 27432
rect 0 27374 2839 27376
rect 0 27344 480 27374
rect 2773 27371 2839 27374
rect 0 26346 480 26376
rect 4061 26346 4127 26349
rect 0 26344 4127 26346
rect 0 26288 4066 26344
rect 4122 26288 4127 26344
rect 0 26286 4127 26288
rect 0 26256 480 26286
rect 4061 26283 4127 26286
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 4061 25394 4127 25397
rect 0 25392 4127 25394
rect 0 25336 4066 25392
rect 4122 25336 4127 25392
rect 0 25334 4127 25336
rect 0 25304 480 25334
rect 4061 25331 4127 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 8845 24850 8911 24853
rect 10777 24850 10843 24853
rect 8845 24848 10843 24850
rect 8845 24792 8850 24848
rect 8906 24792 10782 24848
rect 10838 24792 10843 24848
rect 8845 24790 10843 24792
rect 8845 24787 8911 24790
rect 10777 24787 10843 24790
rect 16297 24850 16363 24853
rect 25313 24850 25379 24853
rect 16297 24848 25379 24850
rect 16297 24792 16302 24848
rect 16358 24792 25318 24848
rect 25374 24792 25379 24848
rect 16297 24790 25379 24792
rect 16297 24787 16363 24790
rect 25313 24787 25379 24790
rect 10041 24714 10107 24717
rect 12617 24714 12683 24717
rect 10041 24712 12683 24714
rect 10041 24656 10046 24712
rect 10102 24656 12622 24712
rect 12678 24656 12683 24712
rect 10041 24654 12683 24656
rect 10041 24651 10107 24654
rect 12617 24651 12683 24654
rect 14273 24714 14339 24717
rect 21265 24714 21331 24717
rect 14273 24712 21331 24714
rect 14273 24656 14278 24712
rect 14334 24656 21270 24712
rect 21326 24656 21331 24712
rect 14273 24654 21331 24656
rect 14273 24651 14339 24654
rect 21265 24651 21331 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 14549 24442 14615 24445
rect 16849 24442 16915 24445
rect 14549 24440 16915 24442
rect 14549 24384 14554 24440
rect 14610 24384 16854 24440
rect 16910 24384 16915 24440
rect 14549 24382 16915 24384
rect 14549 24379 14615 24382
rect 16849 24379 16915 24382
rect 0 24306 480 24336
rect 1393 24306 1459 24309
rect 0 24304 1459 24306
rect 0 24248 1398 24304
rect 1454 24248 1459 24304
rect 0 24246 1459 24248
rect 0 24216 480 24246
rect 1393 24243 1459 24246
rect 18229 24306 18295 24309
rect 20069 24306 20135 24309
rect 18229 24304 20135 24306
rect 18229 24248 18234 24304
rect 18290 24248 20074 24304
rect 20130 24248 20135 24304
rect 18229 24246 20135 24248
rect 18229 24243 18295 24246
rect 20069 24243 20135 24246
rect 25497 24306 25563 24309
rect 27337 24306 27403 24309
rect 25497 24304 27403 24306
rect 25497 24248 25502 24304
rect 25558 24248 27342 24304
rect 27398 24248 27403 24304
rect 25497 24246 27403 24248
rect 25497 24243 25563 24246
rect 27337 24243 27403 24246
rect 5257 24170 5323 24173
rect 6637 24170 6703 24173
rect 5257 24168 6703 24170
rect 5257 24112 5262 24168
rect 5318 24112 6642 24168
rect 6698 24112 6703 24168
rect 5257 24110 6703 24112
rect 5257 24107 5323 24110
rect 6637 24107 6703 24110
rect 10777 24170 10843 24173
rect 17953 24170 18019 24173
rect 10777 24168 18019 24170
rect 10777 24112 10782 24168
rect 10838 24112 17958 24168
rect 18014 24112 18019 24168
rect 10777 24110 18019 24112
rect 10777 24107 10843 24110
rect 17953 24107 18019 24110
rect 18965 24170 19031 24173
rect 24209 24170 24275 24173
rect 18965 24168 24275 24170
rect 18965 24112 18970 24168
rect 19026 24112 24214 24168
rect 24270 24112 24275 24168
rect 18965 24110 24275 24112
rect 18965 24107 19031 24110
rect 24209 24107 24275 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 7741 23898 7807 23901
rect 11789 23898 11855 23901
rect 7741 23896 11855 23898
rect 7741 23840 7746 23896
rect 7802 23840 11794 23896
rect 11850 23840 11855 23896
rect 7741 23838 11855 23840
rect 7741 23835 7807 23838
rect 11789 23835 11855 23838
rect 21909 23898 21975 23901
rect 23197 23898 23263 23901
rect 21909 23896 23263 23898
rect 21909 23840 21914 23896
rect 21970 23840 23202 23896
rect 23258 23840 23263 23896
rect 21909 23838 23263 23840
rect 21909 23835 21975 23838
rect 23197 23835 23263 23838
rect 15469 23762 15535 23765
rect 16481 23762 16547 23765
rect 15469 23760 16547 23762
rect 15469 23704 15474 23760
rect 15530 23704 16486 23760
rect 16542 23704 16547 23760
rect 15469 23702 16547 23704
rect 15469 23699 15535 23702
rect 16481 23699 16547 23702
rect 2681 23626 2747 23629
rect 11605 23626 11671 23629
rect 2681 23624 11671 23626
rect 2681 23568 2686 23624
rect 2742 23568 11610 23624
rect 11666 23568 11671 23624
rect 2681 23566 11671 23568
rect 2681 23563 2747 23566
rect 11605 23563 11671 23566
rect 12525 23626 12591 23629
rect 19517 23626 19583 23629
rect 12525 23624 19583 23626
rect 12525 23568 12530 23624
rect 12586 23568 19522 23624
rect 19578 23568 19583 23624
rect 12525 23566 19583 23568
rect 12525 23563 12591 23566
rect 19517 23563 19583 23566
rect 1485 23490 1551 23493
rect 3325 23490 3391 23493
rect 1485 23488 3391 23490
rect 1485 23432 1490 23488
rect 1546 23432 3330 23488
rect 3386 23432 3391 23488
rect 1485 23430 3391 23432
rect 1485 23427 1551 23430
rect 3325 23427 3391 23430
rect 8477 23490 8543 23493
rect 9857 23490 9923 23493
rect 8477 23488 9923 23490
rect 8477 23432 8482 23488
rect 8538 23432 9862 23488
rect 9918 23432 9923 23488
rect 8477 23430 9923 23432
rect 8477 23427 8543 23430
rect 9857 23427 9923 23430
rect 14457 23490 14523 23493
rect 15377 23490 15443 23493
rect 14457 23488 15443 23490
rect 14457 23432 14462 23488
rect 14518 23432 15382 23488
rect 15438 23432 15443 23488
rect 14457 23430 15443 23432
rect 14457 23427 14523 23430
rect 15377 23427 15443 23430
rect 16205 23490 16271 23493
rect 17953 23490 18019 23493
rect 16205 23488 18019 23490
rect 16205 23432 16210 23488
rect 16266 23432 17958 23488
rect 18014 23432 18019 23488
rect 16205 23430 18019 23432
rect 16205 23427 16271 23430
rect 17953 23427 18019 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23218 480 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 480 23158
rect 1393 23155 1459 23158
rect 5625 23218 5691 23221
rect 12525 23218 12591 23221
rect 5625 23216 12591 23218
rect 5625 23160 5630 23216
rect 5686 23160 12530 23216
rect 12586 23160 12591 23216
rect 5625 23158 12591 23160
rect 5625 23155 5691 23158
rect 12525 23155 12591 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2681 22538 2747 22541
rect 13537 22538 13603 22541
rect 2681 22536 13603 22538
rect 2681 22480 2686 22536
rect 2742 22480 13542 22536
rect 13598 22480 13603 22536
rect 2681 22478 13603 22480
rect 2681 22475 2747 22478
rect 13537 22475 13603 22478
rect 16113 22402 16179 22405
rect 18505 22402 18571 22405
rect 16113 22400 18571 22402
rect 16113 22344 16118 22400
rect 16174 22344 18510 22400
rect 18566 22344 18571 22400
rect 16113 22342 18571 22344
rect 16113 22339 16179 22342
rect 18505 22339 18571 22342
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1393 22266 1459 22269
rect 0 22264 1459 22266
rect 0 22208 1398 22264
rect 1454 22208 1459 22264
rect 0 22206 1459 22208
rect 0 22176 480 22206
rect 1393 22203 1459 22206
rect 11881 22266 11947 22269
rect 19333 22266 19399 22269
rect 11881 22264 19399 22266
rect 11881 22208 11886 22264
rect 11942 22208 19338 22264
rect 19394 22208 19399 22264
rect 11881 22206 19399 22208
rect 11881 22203 11947 22206
rect 19333 22203 19399 22206
rect 16389 22130 16455 22133
rect 18045 22130 18111 22133
rect 16389 22128 18111 22130
rect 16389 22072 16394 22128
rect 16450 22072 18050 22128
rect 18106 22072 18111 22128
rect 16389 22070 18111 22072
rect 16389 22067 16455 22070
rect 18045 22067 18111 22070
rect 6913 21994 6979 21997
rect 10777 21994 10843 21997
rect 6913 21992 10843 21994
rect 6913 21936 6918 21992
rect 6974 21936 10782 21992
rect 10838 21936 10843 21992
rect 6913 21934 10843 21936
rect 6913 21931 6979 21934
rect 10777 21931 10843 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 473 21586 539 21589
rect 3417 21586 3483 21589
rect 473 21584 3483 21586
rect 473 21528 478 21584
rect 534 21528 3422 21584
rect 3478 21528 3483 21584
rect 473 21526 3483 21528
rect 473 21523 539 21526
rect 3417 21523 3483 21526
rect 2681 21450 2747 21453
rect 15561 21450 15627 21453
rect 2681 21448 15627 21450
rect 2681 21392 2686 21448
rect 2742 21392 15566 21448
rect 15622 21392 15627 21448
rect 2681 21390 15627 21392
rect 2681 21387 2747 21390
rect 15561 21387 15627 21390
rect 2313 21314 2379 21317
rect 4061 21314 4127 21317
rect 2313 21312 4127 21314
rect 2313 21256 2318 21312
rect 2374 21256 4066 21312
rect 4122 21256 4127 21312
rect 2313 21254 4127 21256
rect 2313 21251 2379 21254
rect 4061 21251 4127 21254
rect 8201 21314 8267 21317
rect 10041 21314 10107 21317
rect 8201 21312 10107 21314
rect 8201 21256 8206 21312
rect 8262 21256 10046 21312
rect 10102 21256 10107 21312
rect 8201 21254 10107 21256
rect 8201 21251 8267 21254
rect 10041 21251 10107 21254
rect 10277 21248 10597 21249
rect 0 21178 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 480 21118
rect 1393 21115 1459 21118
rect 1577 21178 1643 21181
rect 4521 21178 4587 21181
rect 1577 21176 4587 21178
rect 1577 21120 1582 21176
rect 1638 21120 4526 21176
rect 4582 21120 4587 21176
rect 1577 21118 4587 21120
rect 1577 21115 1643 21118
rect 4521 21115 4587 21118
rect 11513 21178 11579 21181
rect 13721 21178 13787 21181
rect 13997 21178 14063 21181
rect 11513 21176 14063 21178
rect 11513 21120 11518 21176
rect 11574 21120 13726 21176
rect 13782 21120 14002 21176
rect 14058 21120 14063 21176
rect 11513 21118 14063 21120
rect 11513 21115 11579 21118
rect 13721 21115 13787 21118
rect 13997 21115 14063 21118
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2221 20362 2287 20365
rect 13537 20362 13603 20365
rect 2221 20360 13603 20362
rect 2221 20304 2226 20360
rect 2282 20304 13542 20360
rect 13598 20304 13603 20360
rect 2221 20302 13603 20304
rect 2221 20299 2287 20302
rect 13537 20299 13603 20302
rect 6453 20226 6519 20229
rect 7741 20226 7807 20229
rect 6453 20224 7807 20226
rect 6453 20168 6458 20224
rect 6514 20168 7746 20224
rect 7802 20168 7807 20224
rect 6453 20166 7807 20168
rect 6453 20163 6519 20166
rect 7741 20163 7807 20166
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 2313 20090 2379 20093
rect 0 20088 2379 20090
rect 0 20032 2318 20088
rect 2374 20032 2379 20088
rect 0 20030 2379 20032
rect 0 20000 480 20030
rect 2313 20027 2379 20030
rect 2037 19954 2103 19957
rect 2865 19954 2931 19957
rect 2037 19952 2931 19954
rect 2037 19896 2042 19952
rect 2098 19896 2870 19952
rect 2926 19896 2931 19952
rect 2037 19894 2931 19896
rect 2037 19891 2103 19894
rect 2865 19891 2931 19894
rect 13077 19954 13143 19957
rect 15469 19954 15535 19957
rect 13077 19952 15535 19954
rect 13077 19896 13082 19952
rect 13138 19896 15474 19952
rect 15530 19896 15535 19952
rect 13077 19894 15535 19896
rect 13077 19891 13143 19894
rect 15469 19891 15535 19894
rect 2497 19818 2563 19821
rect 14365 19818 14431 19821
rect 2497 19816 14431 19818
rect 2497 19760 2502 19816
rect 2558 19760 14370 19816
rect 14426 19760 14431 19816
rect 2497 19758 14431 19760
rect 2497 19755 2563 19758
rect 14365 19755 14431 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 4981 19274 5047 19277
rect 6361 19274 6427 19277
rect 4981 19272 6427 19274
rect 4981 19216 4986 19272
rect 5042 19216 6366 19272
rect 6422 19216 6427 19272
rect 4981 19214 6427 19216
rect 4981 19211 5047 19214
rect 6361 19211 6427 19214
rect 14549 19274 14615 19277
rect 18045 19274 18111 19277
rect 23565 19274 23631 19277
rect 14549 19272 18111 19274
rect 14549 19216 14554 19272
rect 14610 19216 18050 19272
rect 18106 19216 18111 19272
rect 14549 19214 18111 19216
rect 14549 19211 14615 19214
rect 18045 19211 18111 19214
rect 18278 19272 23631 19274
rect 18278 19216 23570 19272
rect 23626 19216 23631 19272
rect 18278 19214 23631 19216
rect 0 19138 480 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 480 19078
rect 2773 19075 2839 19078
rect 3785 19138 3851 19141
rect 8293 19138 8359 19141
rect 3785 19136 8359 19138
rect 3785 19080 3790 19136
rect 3846 19080 8298 19136
rect 8354 19080 8359 19136
rect 3785 19078 8359 19080
rect 3785 19075 3851 19078
rect 8293 19075 8359 19078
rect 16941 19138 17007 19141
rect 18278 19138 18338 19214
rect 23565 19211 23631 19214
rect 16941 19136 18338 19138
rect 16941 19080 16946 19136
rect 17002 19080 18338 19136
rect 16941 19078 18338 19080
rect 16941 19075 17007 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2497 18594 2563 18597
rect 2497 18592 4538 18594
rect 2497 18536 2502 18592
rect 2558 18536 4538 18592
rect 2497 18534 4538 18536
rect 2497 18531 2563 18534
rect 2405 18458 2471 18461
rect 4337 18458 4403 18461
rect 2405 18456 4403 18458
rect 2405 18400 2410 18456
rect 2466 18400 4342 18456
rect 4398 18400 4403 18456
rect 2405 18398 4403 18400
rect 2405 18395 2471 18398
rect 4337 18395 4403 18398
rect 1945 18322 2011 18325
rect 4478 18322 4538 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 15193 18322 15259 18325
rect 1945 18320 3066 18322
rect 1945 18264 1950 18320
rect 2006 18264 3066 18320
rect 1945 18262 3066 18264
rect 4478 18320 15259 18322
rect 4478 18264 15198 18320
rect 15254 18264 15259 18320
rect 4478 18262 15259 18264
rect 1945 18259 2011 18262
rect 2865 18186 2931 18189
rect 1534 18184 2931 18186
rect 1534 18128 2870 18184
rect 2926 18128 2931 18184
rect 1534 18126 2931 18128
rect 3006 18186 3066 18262
rect 15193 18259 15259 18262
rect 5533 18186 5599 18189
rect 8477 18186 8543 18189
rect 3006 18184 8543 18186
rect 3006 18128 5538 18184
rect 5594 18128 8482 18184
rect 8538 18128 8543 18184
rect 3006 18126 8543 18128
rect 0 18050 480 18080
rect 1534 18050 1594 18126
rect 2865 18123 2931 18126
rect 5533 18123 5599 18126
rect 8477 18123 8543 18126
rect 12157 18186 12223 18189
rect 13905 18186 13971 18189
rect 12157 18184 13971 18186
rect 12157 18128 12162 18184
rect 12218 18128 13910 18184
rect 13966 18128 13971 18184
rect 12157 18126 13971 18128
rect 12157 18123 12223 18126
rect 13905 18123 13971 18126
rect 0 17990 1594 18050
rect 1853 18050 1919 18053
rect 4889 18050 4955 18053
rect 1853 18048 4955 18050
rect 1853 17992 1858 18048
rect 1914 17992 4894 18048
rect 4950 17992 4955 18048
rect 1853 17990 4955 17992
rect 0 17960 480 17990
rect 1853 17987 1919 17990
rect 4889 17987 4955 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5349 17914 5415 17917
rect 9029 17914 9095 17917
rect 5349 17912 9095 17914
rect 5349 17856 5354 17912
rect 5410 17856 9034 17912
rect 9090 17856 9095 17912
rect 5349 17854 9095 17856
rect 5349 17851 5415 17854
rect 9029 17851 9095 17854
rect 8661 17778 8727 17781
rect 11881 17778 11947 17781
rect 8661 17776 11947 17778
rect 8661 17720 8666 17776
rect 8722 17720 11886 17776
rect 11942 17720 11947 17776
rect 8661 17718 11947 17720
rect 8661 17715 8727 17718
rect 11881 17715 11947 17718
rect 7557 17642 7623 17645
rect 9857 17642 9923 17645
rect 7557 17640 9923 17642
rect 7557 17584 7562 17640
rect 7618 17584 9862 17640
rect 9918 17584 9923 17640
rect 7557 17582 9923 17584
rect 7557 17579 7623 17582
rect 9857 17579 9923 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 4061 17234 4127 17237
rect 5533 17234 5599 17237
rect 4061 17232 5599 17234
rect 4061 17176 4066 17232
rect 4122 17176 5538 17232
rect 5594 17176 5599 17232
rect 4061 17174 5599 17176
rect 4061 17171 4127 17174
rect 5533 17171 5599 17174
rect 9305 17234 9371 17237
rect 11145 17234 11211 17237
rect 9305 17232 11211 17234
rect 9305 17176 9310 17232
rect 9366 17176 11150 17232
rect 11206 17176 11211 17232
rect 9305 17174 11211 17176
rect 9305 17171 9371 17174
rect 11145 17171 11211 17174
rect 0 17098 480 17128
rect 4245 17098 4311 17101
rect 0 17096 4311 17098
rect 0 17040 4250 17096
rect 4306 17040 4311 17096
rect 0 17038 4311 17040
rect 0 17008 480 17038
rect 4245 17035 4311 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 2129 16690 2195 16693
rect 4061 16690 4127 16693
rect 2129 16688 4127 16690
rect 2129 16632 2134 16688
rect 2190 16632 4066 16688
rect 4122 16632 4127 16688
rect 2129 16630 4127 16632
rect 2129 16627 2195 16630
rect 4061 16627 4127 16630
rect 7741 16690 7807 16693
rect 9949 16690 10015 16693
rect 7741 16688 10015 16690
rect 7741 16632 7746 16688
rect 7802 16632 9954 16688
rect 10010 16632 10015 16688
rect 7741 16630 10015 16632
rect 7741 16627 7807 16630
rect 9949 16627 10015 16630
rect 13261 16690 13327 16693
rect 15469 16690 15535 16693
rect 13261 16688 15535 16690
rect 13261 16632 13266 16688
rect 13322 16632 15474 16688
rect 15530 16632 15535 16688
rect 13261 16630 15535 16632
rect 13261 16627 13327 16630
rect 15469 16627 15535 16630
rect 18597 16690 18663 16693
rect 23473 16690 23539 16693
rect 18597 16688 23539 16690
rect 18597 16632 18602 16688
rect 18658 16632 23478 16688
rect 23534 16632 23539 16688
rect 18597 16630 23539 16632
rect 18597 16627 18663 16630
rect 23473 16627 23539 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16010 480 16040
rect 4245 16010 4311 16013
rect 0 16008 4311 16010
rect 0 15952 4250 16008
rect 4306 15952 4311 16008
rect 0 15950 4311 15952
rect 0 15920 480 15950
rect 4245 15947 4311 15950
rect 13629 15874 13695 15877
rect 15377 15874 15443 15877
rect 13629 15872 15443 15874
rect 13629 15816 13634 15872
rect 13690 15816 15382 15872
rect 15438 15816 15443 15872
rect 13629 15814 15443 15816
rect 13629 15811 13695 15814
rect 15377 15811 15443 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 8201 15602 8267 15605
rect 9857 15602 9923 15605
rect 8158 15600 9923 15602
rect 8158 15544 8206 15600
rect 8262 15544 9862 15600
rect 9918 15544 9923 15600
rect 8158 15542 9923 15544
rect 8158 15539 8267 15542
rect 9857 15539 9923 15542
rect 6637 15466 6703 15469
rect 8158 15466 8218 15539
rect 6637 15464 8218 15466
rect 6637 15408 6642 15464
rect 6698 15408 8218 15464
rect 6637 15406 8218 15408
rect 12065 15466 12131 15469
rect 19517 15466 19583 15469
rect 12065 15464 19583 15466
rect 12065 15408 12070 15464
rect 12126 15408 19522 15464
rect 19578 15408 19583 15464
rect 12065 15406 19583 15408
rect 6637 15403 6703 15406
rect 12065 15403 12131 15406
rect 19517 15403 19583 15406
rect 8017 15330 8083 15333
rect 10685 15330 10751 15333
rect 8017 15328 10751 15330
rect 8017 15272 8022 15328
rect 8078 15272 10690 15328
rect 10746 15272 10751 15328
rect 8017 15270 10751 15272
rect 8017 15267 8083 15270
rect 10685 15267 10751 15270
rect 15837 15330 15903 15333
rect 19333 15330 19399 15333
rect 15837 15328 19399 15330
rect 15837 15272 15842 15328
rect 15898 15272 19338 15328
rect 19394 15272 19399 15328
rect 15837 15270 19399 15272
rect 15837 15267 15903 15270
rect 19333 15267 19399 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 9673 15058 9739 15061
rect 9949 15058 10015 15061
rect 16665 15058 16731 15061
rect 9673 15056 16731 15058
rect 9673 15000 9678 15056
rect 9734 15000 9954 15056
rect 10010 15000 16670 15056
rect 16726 15000 16731 15056
rect 9673 14998 16731 15000
rect 9673 14995 9739 14998
rect 9949 14995 10015 14998
rect 16665 14995 16731 14998
rect 0 14922 480 14952
rect 2589 14922 2655 14925
rect 5901 14922 5967 14925
rect 0 14862 2514 14922
rect 0 14832 480 14862
rect 2454 14514 2514 14862
rect 2589 14920 5967 14922
rect 2589 14864 2594 14920
rect 2650 14864 5906 14920
rect 5962 14864 5967 14920
rect 2589 14862 5967 14864
rect 2589 14859 2655 14862
rect 5901 14859 5967 14862
rect 10961 14922 11027 14925
rect 13997 14922 14063 14925
rect 15653 14922 15719 14925
rect 16573 14922 16639 14925
rect 10961 14920 16639 14922
rect 10961 14864 10966 14920
rect 11022 14864 14002 14920
rect 14058 14864 15658 14920
rect 15714 14864 16578 14920
rect 16634 14864 16639 14920
rect 10961 14862 16639 14864
rect 10961 14859 11027 14862
rect 13997 14859 14063 14862
rect 15653 14859 15719 14862
rect 16573 14859 16639 14862
rect 3233 14786 3299 14789
rect 6637 14786 6703 14789
rect 3233 14784 6703 14786
rect 3233 14728 3238 14784
rect 3294 14728 6642 14784
rect 6698 14728 6703 14784
rect 3233 14726 6703 14728
rect 3233 14723 3299 14726
rect 6637 14723 6703 14726
rect 12709 14786 12775 14789
rect 16849 14786 16915 14789
rect 12709 14784 16915 14786
rect 12709 14728 12714 14784
rect 12770 14728 16854 14784
rect 16910 14728 16915 14784
rect 12709 14726 16915 14728
rect 12709 14723 12775 14726
rect 16849 14723 16915 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 5257 14650 5323 14653
rect 6729 14650 6795 14653
rect 5257 14648 6795 14650
rect 5257 14592 5262 14648
rect 5318 14592 6734 14648
rect 6790 14592 6795 14648
rect 5257 14590 6795 14592
rect 5257 14587 5323 14590
rect 6729 14587 6795 14590
rect 5533 14514 5599 14517
rect 2454 14512 5599 14514
rect 2454 14456 5538 14512
rect 5594 14456 5599 14512
rect 2454 14454 5599 14456
rect 5533 14451 5599 14454
rect 10041 14514 10107 14517
rect 16849 14514 16915 14517
rect 10041 14512 16915 14514
rect 10041 14456 10046 14512
rect 10102 14456 16854 14512
rect 16910 14456 16915 14512
rect 10041 14454 16915 14456
rect 10041 14451 10107 14454
rect 16849 14451 16915 14454
rect 9121 14378 9187 14381
rect 10869 14378 10935 14381
rect 15745 14378 15811 14381
rect 9121 14376 15811 14378
rect 9121 14320 9126 14376
rect 9182 14320 10874 14376
rect 10930 14320 15750 14376
rect 15806 14320 15811 14376
rect 9121 14318 15811 14320
rect 9121 14315 9187 14318
rect 10869 14315 10935 14318
rect 15745 14315 15811 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13970 480 14000
rect 3601 13970 3667 13973
rect 0 13968 3667 13970
rect 0 13912 3606 13968
rect 3662 13912 3667 13968
rect 0 13910 3667 13912
rect 0 13880 480 13910
rect 3601 13907 3667 13910
rect 7557 13970 7623 13973
rect 10225 13970 10291 13973
rect 11329 13970 11395 13973
rect 12893 13970 12959 13973
rect 7557 13968 12959 13970
rect 7557 13912 7562 13968
rect 7618 13912 10230 13968
rect 10286 13912 11334 13968
rect 11390 13912 12898 13968
rect 12954 13912 12959 13968
rect 7557 13910 12959 13912
rect 7557 13907 7623 13910
rect 10225 13907 10291 13910
rect 11329 13907 11395 13910
rect 12893 13907 12959 13910
rect 15377 13970 15443 13973
rect 17953 13970 18019 13973
rect 15377 13968 18019 13970
rect 15377 13912 15382 13968
rect 15438 13912 17958 13968
rect 18014 13912 18019 13968
rect 15377 13910 18019 13912
rect 15377 13907 15443 13910
rect 17953 13907 18019 13910
rect 13077 13834 13143 13837
rect 15469 13834 15535 13837
rect 13077 13832 15535 13834
rect 13077 13776 13082 13832
rect 13138 13776 15474 13832
rect 15530 13776 15535 13832
rect 13077 13774 15535 13776
rect 13077 13771 13143 13774
rect 15469 13771 15535 13774
rect 3233 13698 3299 13701
rect 3509 13698 3575 13701
rect 5717 13698 5783 13701
rect 3233 13696 5783 13698
rect 3233 13640 3238 13696
rect 3294 13640 3514 13696
rect 3570 13640 5722 13696
rect 5778 13640 5783 13696
rect 3233 13638 5783 13640
rect 3233 13635 3299 13638
rect 3509 13635 3575 13638
rect 5717 13635 5783 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 6453 13426 6519 13429
rect 13169 13426 13235 13429
rect 6453 13424 13235 13426
rect 6453 13368 6458 13424
rect 6514 13368 13174 13424
rect 13230 13368 13235 13424
rect 6453 13366 13235 13368
rect 6453 13363 6519 13366
rect 13169 13363 13235 13366
rect 8753 13290 8819 13293
rect 13813 13290 13879 13293
rect 8753 13288 13879 13290
rect 8753 13232 8758 13288
rect 8814 13232 13818 13288
rect 13874 13232 13879 13288
rect 8753 13230 13879 13232
rect 8753 13227 8819 13230
rect 13813 13227 13879 13230
rect 9857 13154 9923 13157
rect 13077 13154 13143 13157
rect 13813 13154 13879 13157
rect 9857 13152 13879 13154
rect 9857 13096 9862 13152
rect 9918 13096 13082 13152
rect 13138 13096 13818 13152
rect 13874 13096 13879 13152
rect 9857 13094 13879 13096
rect 9857 13091 9923 13094
rect 13077 13091 13143 13094
rect 13813 13091 13879 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12882 480 12912
rect 6453 12882 6519 12885
rect 0 12880 6519 12882
rect 0 12824 6458 12880
rect 6514 12824 6519 12880
rect 0 12822 6519 12824
rect 0 12792 480 12822
rect 6453 12819 6519 12822
rect 9765 12882 9831 12885
rect 12801 12882 12867 12885
rect 9765 12880 12867 12882
rect 9765 12824 9770 12880
rect 9826 12824 12806 12880
rect 12862 12824 12867 12880
rect 9765 12822 12867 12824
rect 9765 12819 9831 12822
rect 12801 12819 12867 12822
rect 8661 12746 8727 12749
rect 12709 12746 12775 12749
rect 8661 12744 12775 12746
rect 8661 12688 8666 12744
rect 8722 12688 12714 12744
rect 12770 12688 12775 12744
rect 8661 12686 12775 12688
rect 8661 12683 8727 12686
rect 12709 12683 12775 12686
rect 2681 12610 2747 12613
rect 3049 12610 3115 12613
rect 2681 12608 3115 12610
rect 2681 12552 2686 12608
rect 2742 12552 3054 12608
rect 3110 12552 3115 12608
rect 2681 12550 3115 12552
rect 2681 12547 2747 12550
rect 3049 12547 3115 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5257 12338 5323 12341
rect 12433 12338 12499 12341
rect 5257 12336 12499 12338
rect 5257 12280 5262 12336
rect 5318 12280 12438 12336
rect 12494 12280 12499 12336
rect 5257 12278 12499 12280
rect 5257 12275 5323 12278
rect 12433 12275 12499 12278
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 6085 11930 6151 11933
rect 10041 11930 10107 11933
rect 6085 11928 10107 11930
rect 6085 11872 6090 11928
rect 6146 11872 10046 11928
rect 10102 11872 10107 11928
rect 6085 11870 10107 11872
rect 6085 11867 6151 11870
rect 10041 11867 10107 11870
rect 0 11794 480 11824
rect 1669 11794 1735 11797
rect 0 11792 1735 11794
rect 0 11736 1674 11792
rect 1730 11736 1735 11792
rect 0 11734 1735 11736
rect 0 11704 480 11734
rect 1669 11731 1735 11734
rect 3049 11794 3115 11797
rect 4797 11794 4863 11797
rect 3049 11792 4863 11794
rect 3049 11736 3054 11792
rect 3110 11736 4802 11792
rect 4858 11736 4863 11792
rect 3049 11734 4863 11736
rect 3049 11731 3115 11734
rect 4797 11731 4863 11734
rect 5073 11794 5139 11797
rect 6913 11794 6979 11797
rect 12157 11794 12223 11797
rect 5073 11792 12223 11794
rect 5073 11736 5078 11792
rect 5134 11736 6918 11792
rect 6974 11736 12162 11792
rect 12218 11736 12223 11792
rect 5073 11734 12223 11736
rect 5073 11731 5139 11734
rect 6913 11731 6979 11734
rect 12157 11731 12223 11734
rect 9305 11658 9371 11661
rect 11973 11658 12039 11661
rect 9305 11656 12039 11658
rect 9305 11600 9310 11656
rect 9366 11600 11978 11656
rect 12034 11600 12039 11656
rect 9305 11598 12039 11600
rect 9305 11595 9371 11598
rect 11973 11595 12039 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2129 11386 2195 11389
rect 5533 11386 5599 11389
rect 2129 11384 5599 11386
rect 2129 11328 2134 11384
rect 2190 11328 5538 11384
rect 5594 11328 5599 11384
rect 2129 11326 5599 11328
rect 2129 11323 2195 11326
rect 5533 11323 5599 11326
rect 2497 11250 2563 11253
rect 5073 11250 5139 11253
rect 2497 11248 5139 11250
rect 2497 11192 2502 11248
rect 2558 11192 5078 11248
rect 5134 11192 5139 11248
rect 2497 11190 5139 11192
rect 2497 11187 2563 11190
rect 5073 11187 5139 11190
rect 6269 11250 6335 11253
rect 14457 11250 14523 11253
rect 6269 11248 14523 11250
rect 6269 11192 6274 11248
rect 6330 11192 14462 11248
rect 14518 11192 14523 11248
rect 6269 11190 14523 11192
rect 6269 11187 6335 11190
rect 14457 11187 14523 11190
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 1577 10842 1643 10845
rect 0 10840 1643 10842
rect 0 10784 1582 10840
rect 1638 10784 1643 10840
rect 0 10782 1643 10784
rect 0 10752 480 10782
rect 1577 10779 1643 10782
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 7925 10162 7991 10165
rect 11237 10162 11303 10165
rect 7925 10160 11303 10162
rect 7925 10104 7930 10160
rect 7986 10104 11242 10160
rect 11298 10104 11303 10160
rect 7925 10102 11303 10104
rect 7925 10099 7991 10102
rect 11237 10099 11303 10102
rect 5610 9824 5930 9825
rect 0 9754 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1761 9754 1827 9757
rect 0 9752 1827 9754
rect 0 9696 1766 9752
rect 1822 9696 1827 9752
rect 0 9694 1827 9696
rect 0 9664 480 9694
rect 1761 9691 1827 9694
rect 2681 9754 2747 9757
rect 4797 9754 4863 9757
rect 2681 9752 4863 9754
rect 2681 9696 2686 9752
rect 2742 9696 4802 9752
rect 4858 9696 4863 9752
rect 2681 9694 4863 9696
rect 2681 9691 2747 9694
rect 4797 9691 4863 9694
rect 6545 9754 6611 9757
rect 9673 9754 9739 9757
rect 6545 9752 9739 9754
rect 6545 9696 6550 9752
rect 6606 9696 9678 9752
rect 9734 9696 9739 9752
rect 6545 9694 9739 9696
rect 6545 9691 6611 9694
rect 9673 9691 9739 9694
rect 8201 9346 8267 9349
rect 9765 9346 9831 9349
rect 8201 9344 9831 9346
rect 8201 9288 8206 9344
rect 8262 9288 9770 9344
rect 9826 9288 9831 9344
rect 8201 9286 9831 9288
rect 8201 9283 8267 9286
rect 9765 9283 9831 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 1669 9074 1735 9077
rect 5533 9074 5599 9077
rect 1669 9072 5599 9074
rect 1669 9016 1674 9072
rect 1730 9016 5538 9072
rect 5594 9016 5599 9072
rect 1669 9014 5599 9016
rect 1669 9011 1735 9014
rect 5533 9011 5599 9014
rect 0 8802 480 8832
rect 3877 8802 3943 8805
rect 0 8800 3943 8802
rect 0 8744 3882 8800
rect 3938 8744 3943 8800
rect 0 8742 3943 8744
rect 0 8712 480 8742
rect 3877 8739 3943 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 5625 8530 5691 8533
rect 8937 8530 9003 8533
rect 5625 8528 9003 8530
rect 5625 8472 5630 8528
rect 5686 8472 8942 8528
rect 8998 8472 9003 8528
rect 5625 8470 9003 8472
rect 5625 8467 5691 8470
rect 8937 8467 9003 8470
rect 2221 8258 2287 8261
rect 8293 8258 8359 8261
rect 2221 8256 8359 8258
rect 2221 8200 2226 8256
rect 2282 8200 8298 8256
rect 8354 8200 8359 8256
rect 2221 8198 8359 8200
rect 2221 8195 2287 8198
rect 8293 8195 8359 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 0 7714 480 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 480 7654
rect 1485 7651 1551 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 3601 7578 3667 7581
rect 4981 7578 5047 7581
rect 3601 7576 5047 7578
rect 3601 7520 3606 7576
rect 3662 7520 4986 7576
rect 5042 7520 5047 7576
rect 3601 7518 5047 7520
rect 3601 7515 3667 7518
rect 4981 7515 5047 7518
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 4061 6898 4127 6901
rect 6085 6898 6151 6901
rect 4061 6896 6151 6898
rect 4061 6840 4066 6896
rect 4122 6840 6090 6896
rect 6146 6840 6151 6896
rect 4061 6838 6151 6840
rect 4061 6835 4127 6838
rect 6085 6835 6151 6838
rect 0 6626 480 6656
rect 1761 6626 1827 6629
rect 0 6624 1827 6626
rect 0 6568 1766 6624
rect 1822 6568 1827 6624
rect 0 6566 1827 6568
rect 0 6536 480 6566
rect 1761 6563 1827 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 2405 6218 2471 6221
rect 11053 6218 11119 6221
rect 2405 6216 11119 6218
rect 2405 6160 2410 6216
rect 2466 6160 11058 6216
rect 11114 6160 11119 6216
rect 2405 6158 11119 6160
rect 2405 6155 2471 6158
rect 11053 6155 11119 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 2589 5946 2655 5949
rect 5349 5946 5415 5949
rect 2589 5944 5415 5946
rect 2589 5888 2594 5944
rect 2650 5888 5354 5944
rect 5410 5888 5415 5944
rect 2589 5886 5415 5888
rect 2589 5883 2655 5886
rect 5349 5883 5415 5886
rect 0 5674 480 5704
rect 1393 5674 1459 5677
rect 0 5672 1459 5674
rect 0 5616 1398 5672
rect 1454 5616 1459 5672
rect 0 5614 1459 5616
rect 0 5584 480 5614
rect 1393 5611 1459 5614
rect 9581 5538 9647 5541
rect 12249 5538 12315 5541
rect 9581 5536 12315 5538
rect 9581 5480 9586 5536
rect 9642 5480 12254 5536
rect 12310 5480 12315 5536
rect 9581 5478 12315 5480
rect 9581 5475 9647 5478
rect 12249 5475 12315 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 1761 4722 1827 4725
rect 7557 4722 7623 4725
rect 1761 4720 7623 4722
rect 1761 4664 1766 4720
rect 1822 4664 7562 4720
rect 7618 4664 7623 4720
rect 1761 4662 7623 4664
rect 1761 4659 1827 4662
rect 7557 4659 7623 4662
rect 0 4586 480 4616
rect 1393 4586 1459 4589
rect 0 4584 1459 4586
rect 0 4528 1398 4584
rect 1454 4528 1459 4584
rect 0 4526 1459 4528
rect 0 4496 480 4526
rect 1393 4523 1459 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 5257 4042 5323 4045
rect 7281 4042 7347 4045
rect 5257 4040 7347 4042
rect 5257 3984 5262 4040
rect 5318 3984 7286 4040
rect 7342 3984 7347 4040
rect 5257 3982 7347 3984
rect 5257 3979 5323 3982
rect 7281 3979 7347 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3498 480 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 480 3438
rect 1393 3435 1459 3438
rect 1577 3498 1643 3501
rect 6729 3498 6795 3501
rect 1577 3496 6795 3498
rect 1577 3440 1582 3496
rect 1638 3440 6734 3496
rect 6790 3440 6795 3496
rect 1577 3438 6795 3440
rect 1577 3435 1643 3438
rect 6729 3435 6795 3438
rect 16481 3498 16547 3501
rect 26233 3498 26299 3501
rect 16481 3496 26299 3498
rect 16481 3440 16486 3496
rect 16542 3440 26238 3496
rect 26294 3440 26299 3496
rect 16481 3438 26299 3440
rect 16481 3435 16547 3438
rect 26233 3435 26299 3438
rect 15469 3362 15535 3365
rect 22737 3362 22803 3365
rect 15469 3360 22803 3362
rect 15469 3304 15474 3360
rect 15530 3304 22742 3360
rect 22798 3304 22803 3360
rect 15469 3302 22803 3304
rect 15469 3299 15535 3302
rect 22737 3299 22803 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1577 2682 1643 2685
rect 6177 2682 6243 2685
rect 1577 2680 6243 2682
rect 1577 2624 1582 2680
rect 1638 2624 6182 2680
rect 6238 2624 6243 2680
rect 1577 2622 6243 2624
rect 1577 2619 1643 2622
rect 6177 2619 6243 2622
rect 0 2546 480 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 480 2486
rect 1393 2483 1459 2486
rect 2681 2410 2747 2413
rect 10133 2410 10199 2413
rect 2681 2408 10199 2410
rect 2681 2352 2686 2408
rect 2742 2352 10138 2408
rect 10194 2352 10199 2408
rect 2681 2350 10199 2352
rect 2681 2347 2747 2350
rect 10133 2347 10199 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 1458 480 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 480 1398
rect 1485 1395 1551 1398
rect 0 506 480 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 480 446
rect 2865 443 2931 446
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_17
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_21 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_14 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_54
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_buf_2  _233_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_22
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use scs8hd_inv_8  _101_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_81
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_12
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_20
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_24
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 774 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_conb_1  _209_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_21
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_25
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_47
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_69
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_109
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_113
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _158_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_78
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _153_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_99
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_103
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 590 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_60
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_4  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_88
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _122_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_18_98
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_112
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_116
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_8
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_76
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_109
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_159
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_171
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_183
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_164
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_17
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_25
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_49
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_161
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_172
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_184
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 1472 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_13
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_34
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 6900 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_72
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_165
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_172
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_176
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_25
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 406 592
use scs8hd_nor3_4  _169_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_42
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 130 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_60
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_86
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_122
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_139
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_165
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_169
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_13
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_17
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 314 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 12512 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_133
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 590 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_200
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_212
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_224
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_8
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_17
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 866 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_40
timestamp 1586364061
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_78
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_82
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_85
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_96
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_103
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_100
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_133
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_155
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_158
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_162
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_173
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 590 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_188
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_192
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_216
timestamp 1586364061
transform 1 0 20976 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_228
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_38
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_66
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_132
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_182
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_193
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_20
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_150
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_154
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_167
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_205
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_241
timestamp 1586364061
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_49
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_63
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_78
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_151
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_173
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_197
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_209
timestamp 1586364061
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_14
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_55
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 8280 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_140
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_170
timestamp 1586364061
transform 1 0 16744 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_200
timestamp 1586364061
transform 1 0 19504 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_212
timestamp 1586364061
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 774 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 314 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_17
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 4508 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_28
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_36
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_54
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_65
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_65
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_109
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_107
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_115
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_115
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_129
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_133
timestamp 1586364061
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_148
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_152
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_142
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_150
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_165
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_169
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_169
timestamp 1586364061
transform 1 0 16652 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_181
timestamp 1586364061
transform 1 0 17756 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_203
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_205
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_215
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_227
timestamp 1586364061
transform 1 0 21988 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_239
timestamp 1586364061
transform 1 0 23092 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_6
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_10
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_17
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_21
timestamp 1586364061
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_28
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_49
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_70
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 406 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_140
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_173
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_188
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_200
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_212
timestamp 1586364061
transform 1 0 20608 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_224
timestamp 1586364061
transform 1 0 21712 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 774 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_12
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_52
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_4  FILLER_36_67
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_98
timestamp 1586364061
transform 1 0 10120 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 406 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_115
timestamp 1586364061
transform 1 0 11684 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_119
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_132
timestamp 1586364061
transform 1 0 13248 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_157
timestamp 1586364061
transform 1 0 15548 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_161
timestamp 1586364061
transform 1 0 15916 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_174
timestamp 1586364061
transform 1 0 17112 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_203
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_6
timestamp 1586364061
transform 1 0 1656 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_10
timestamp 1586364061
transform 1 0 2024 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_17
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_21
timestamp 1586364061
transform 1 0 3036 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_28
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_32
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_44
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 1142 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_56
timestamp 1586364061
transform 1 0 6256 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_60
timestamp 1586364061
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_66
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_72
timestamp 1586364061
transform 1 0 7728 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_76
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_89
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_99
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  FILLER_37_138
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 590 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_187
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_215
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_239
timestamp 1586364061
transform 1 0 23092 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_17
timestamp 1586364061
transform 1 0 2668 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_29
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_48
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_52
timestamp 1586364061
transform 1 0 5888 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_63
timestamp 1586364061
transform 1 0 6900 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 17112 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_189
timestamp 1586364061
transform 1 0 18492 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_201
timestamp 1586364061
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_25
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_29
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_35
timestamp 1586364061
transform 1 0 4324 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_42
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_47
timestamp 1586364061
transform 1 0 5428 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_62
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_73
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_77
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_70
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_85
timestamp 1586364061
transform 1 0 8924 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_112
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_116
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 13800 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_136
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_144
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_147
timestamp 1586364061
transform 1 0 14628 0 -1 24480
box -38 -48 590 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_175
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_187
timestamp 1586364061
transform 1 0 18308 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_191
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_195
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_200
timestamp 1586364061
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_212
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_212
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_257
timestamp 1586364061
transform 1 0 24748 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_269
timestamp 1586364061
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_66
timestamp 1586364061
transform 1 0 7176 0 1 24480
box -38 -48 130 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_70
timestamp 1586364061
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_90
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_41_96
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 406 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 11500 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_111
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_115
timestamp 1586364061
transform 1 0 11684 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_119
timestamp 1586364061
transform 1 0 12052 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 590 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 222 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_41_167
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_41_174
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_182
timestamp 1586364061
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_84
timestamp 1586364061
transform 1 0 8832 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_92
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_97
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_116
timestamp 1586364061
transform 1 0 11776 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_153
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_162
timestamp 1586364061
transform 1 0 16008 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_174
timestamp 1586364061
transform 1 0 17112 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5262 0 5318 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8758 0 8814 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 12254 0 12310 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15750 0 15806 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 19246 0 19302 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 22742 0 22798 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[1]
port 7 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[2]
port 8 nsew default input
rlabel metal3 s 0 21088 480 21208 6 chanx_left_in[3]
port 9 nsew default input
rlabel metal3 s 0 22176 480 22296 6 chanx_left_in[4]
port 10 nsew default input
rlabel metal3 s 0 23128 480 23248 6 chanx_left_in[5]
port 11 nsew default input
rlabel metal3 s 0 24216 480 24336 6 chanx_left_in[6]
port 12 nsew default input
rlabel metal3 s 0 25304 480 25424 6 chanx_left_in[7]
port 13 nsew default input
rlabel metal3 s 0 26256 480 26376 6 chanx_left_in[8]
port 14 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[0]
port 15 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[1]
port 16 nsew default tristate
rlabel metal3 s 0 10752 480 10872 6 chanx_left_out[2]
port 17 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_left_out[3]
port 18 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[4]
port 19 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[5]
port 20 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[6]
port 21 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[7]
port 22 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[8]
port 23 nsew default tristate
rlabel metal2 s 1490 27520 1546 28000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 8758 27520 8814 28000 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 12898 27520 12954 28000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 14922 27520 14978 28000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 18050 27520 18106 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 data_in
port 42 nsew default input
rlabel metal2 s 1766 0 1822 480 6 enable
port 43 nsew default input
rlabel metal3 s 0 5584 480 5704 6 left_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 0 6536 480 6656 6 left_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal3 s 0 7624 480 7744 6 left_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 0 416 480 536 6 left_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 0 4496 480 4616 6 left_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 0 27344 480 27464 6 left_top_grid_pin_10_
port 52 nsew default input
rlabel metal2 s 478 27520 534 28000 6 top_left_grid_pin_13_
port 53 nsew default input
rlabel metal2 s 25318 27520 25374 28000 6 top_right_grid_pin_11_
port 54 nsew default input
rlabel metal2 s 26330 27520 26386 28000 6 top_right_grid_pin_13_
port 55 nsew default input
rlabel metal2 s 27342 27520 27398 28000 6 top_right_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 20074 27520 20130 28000 6 top_right_grid_pin_1_
port 57 nsew default input
rlabel metal2 s 21178 27520 21234 28000 6 top_right_grid_pin_3_
port 58 nsew default input
rlabel metal2 s 22190 27520 22246 28000 6 top_right_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 23202 27520 23258 28000 6 top_right_grid_pin_7_
port 60 nsew default input
rlabel metal2 s 24214 27520 24270 28000 6 top_right_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< properties >>
string FIXED_BBOX 0 0 27403 28000
<< end >>
