VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_left_left
  CLASS BLOCK ;
  FOREIGN grid_io_left_left ;
  ORIGIN 0.000 0.000 ;
  SIZE 39.670 BY 85.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.800 82.600 6.080 85.000 ;
    END
  END IO_ISOL_N
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.320 0.000 11.600 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.820 0.000 23.100 2.400 ;
    END
  END ccff_tail
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.270 73.480 39.670 74.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.860 0.000 34.140 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.340 82.600 28.620 85.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.280 0.000 0.560 2.400 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.270 31.320 39.670 31.920 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.270 10.240 39.670 10.840 ;
    END
  END right_width_0_height_0__pin_1_lower
  PIN right_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.270 52.400 39.670 53.000 ;
    END
  END right_width_0_height_0__pin_1_upper
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.050 10.640 6.650 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 10.710 10.640 12.310 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 10.795 33.770 73.525 ;
      LAYER met1 ;
        RECT 0.190 10.640 34.160 73.680 ;
      LAYER met2 ;
        RECT 0.290 82.320 5.520 82.600 ;
        RECT 6.360 82.320 28.060 82.600 ;
        RECT 28.900 82.320 34.130 82.600 ;
        RECT 0.290 2.680 34.130 82.320 ;
        RECT 0.840 2.400 11.040 2.680 ;
        RECT 11.880 2.400 22.540 2.680 ;
        RECT 23.380 2.400 33.580 2.680 ;
      LAYER met3 ;
        RECT 5.050 73.080 36.870 73.930 ;
        RECT 5.050 53.400 37.270 73.080 ;
        RECT 5.050 52.000 36.870 53.400 ;
        RECT 5.050 32.320 37.270 52.000 ;
        RECT 5.050 30.920 36.870 32.320 ;
        RECT 5.050 11.240 37.270 30.920 ;
        RECT 5.050 10.390 36.870 11.240 ;
      LAYER met4 ;
        RECT 16.370 10.640 29.290 73.680 ;
  END
END grid_io_left_left
END LIBRARY

