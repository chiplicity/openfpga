VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_top
  CLASS BLOCK ;
  FOREIGN grid_io_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 137.600 7.730 140.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 137.600 22.910 140.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END address[3]
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 82.320 140.000 82.920 ;
    END
  END bottom_width_0_height_0__pin_10_
  PIN bottom_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END bottom_width_0_height_0__pin_11_
  PIN bottom_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END bottom_width_0_height_0__pin_12_
  PIN bottom_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 137.600 85.010 140.000 ;
    END
  END bottom_width_0_height_0__pin_13_
  PIN bottom_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END bottom_width_0_height_0__pin_14_
  PIN bottom_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 137.600 100.650 140.000 ;
    END
  END bottom_width_0_height_0__pin_15_
  PIN bottom_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 56.480 140.000 57.080 ;
    END
  END bottom_width_0_height_0__pin_1_
  PIN bottom_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END bottom_width_0_height_0__pin_2_
  PIN bottom_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END bottom_width_0_height_0__pin_3_
  PIN bottom_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END bottom_width_0_height_0__pin_4_
  PIN bottom_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END bottom_width_0_height_0__pin_5_
  PIN bottom_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END bottom_width_0_height_0__pin_6_
  PIN bottom_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END bottom_width_0_height_0__pin_7_
  PIN bottom_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END bottom_width_0_height_0__pin_8_
  PIN bottom_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 137.600 54.190 140.000 ;
    END
  END bottom_width_0_height_0__pin_9_
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.160 140.000 6.760 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 107.480 140.000 108.080 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 116.010 137.600 116.290 140.000 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 120.400 140.000 121.000 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 133.320 140.000 133.920 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 131.650 137.600 131.930 140.000 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 138.390 128.080 ;
      LAYER met2 ;
        RECT 23.190 137.320 37.990 137.600 ;
        RECT 38.830 137.320 53.630 137.600 ;
        RECT 54.470 137.320 69.270 137.600 ;
        RECT 70.110 137.320 84.450 137.600 ;
        RECT 85.290 137.320 100.090 137.600 ;
        RECT 100.930 137.320 115.730 137.600 ;
        RECT 116.570 137.320 131.370 137.600 ;
        RECT 132.210 137.320 138.370 137.600 ;
        RECT 22.630 8.995 138.370 137.320 ;
      LAYER met3 ;
        RECT 0.310 121.400 138.610 128.005 ;
        RECT 0.310 120.000 137.200 121.400 ;
        RECT 0.310 113.920 138.610 120.000 ;
        RECT 2.800 112.520 138.610 113.920 ;
        RECT 0.310 108.480 138.610 112.520 ;
        RECT 0.310 107.080 137.200 108.480 ;
        RECT 0.310 96.240 138.610 107.080 ;
        RECT 2.800 94.840 137.200 96.240 ;
        RECT 0.310 83.320 138.610 94.840 ;
        RECT 0.310 81.920 137.200 83.320 ;
        RECT 0.310 79.240 138.610 81.920 ;
        RECT 2.800 77.840 138.610 79.240 ;
        RECT 0.310 70.400 138.610 77.840 ;
        RECT 0.310 69.000 137.200 70.400 ;
        RECT 0.310 61.560 138.610 69.000 ;
        RECT 2.800 60.160 138.610 61.560 ;
        RECT 0.310 57.480 138.610 60.160 ;
        RECT 0.310 56.080 137.200 57.480 ;
        RECT 0.310 45.240 138.610 56.080 ;
        RECT 0.310 43.880 137.200 45.240 ;
        RECT 2.800 43.840 137.200 43.880 ;
        RECT 2.800 42.480 138.610 43.840 ;
        RECT 0.310 32.320 138.610 42.480 ;
        RECT 0.310 30.920 137.200 32.320 ;
        RECT 0.310 26.200 138.610 30.920 ;
        RECT 2.800 24.800 138.610 26.200 ;
        RECT 0.310 19.400 138.610 24.800 ;
        RECT 0.310 18.000 137.200 19.400 ;
        RECT 0.310 9.200 138.610 18.000 ;
        RECT 2.800 7.800 138.610 9.200 ;
        RECT 0.310 7.160 138.610 7.800 ;
        RECT 0.310 6.760 137.200 7.160 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END grid_io_top
END LIBRARY

