magic
tech sky130A
magscale 1 2
timestamp 1606425894
<< locali >>
rect 6653 12631 6687 12869
rect 7481 9979 7515 10149
rect 7423 9945 7515 9979
rect 17785 9911 17819 10217
rect 6653 9367 6687 9469
rect 8769 9367 8803 9469
rect 15025 9027 15059 9129
rect 14013 8823 14047 8993
rect 18981 8619 19015 9537
rect 8861 8415 8895 8585
rect 8769 8279 8803 8381
rect 7849 7803 7883 8041
rect 3617 7191 3651 7429
rect 5549 7259 5583 7497
rect 5549 5151 5583 5253
rect 17601 4471 17635 4777
rect 5733 3383 5767 3689
rect 2605 2907 2639 3077
<< viali >>
rect 3433 14569 3467 14603
rect 5457 14569 5491 14603
rect 6469 14569 6503 14603
rect 2053 14501 2087 14535
rect 2789 14501 2823 14535
rect 1777 14433 1811 14467
rect 2513 14433 2547 14467
rect 3249 14433 3283 14467
rect 5273 14433 5307 14467
rect 6285 14433 6319 14467
rect 17601 14025 17635 14059
rect 18245 14025 18279 14059
rect 3249 13957 3283 13991
rect 3801 13957 3835 13991
rect 5549 13957 5583 13991
rect 17049 13957 17083 13991
rect 2605 13889 2639 13923
rect 6101 13889 6135 13923
rect 7389 13889 7423 13923
rect 8309 13889 8343 13923
rect 14473 13889 14507 13923
rect 1593 13821 1627 13855
rect 1869 13821 1903 13855
rect 2329 13821 2363 13855
rect 3065 13821 3099 13855
rect 3617 13821 3651 13855
rect 8033 13821 8067 13855
rect 14197 13821 14231 13855
rect 16865 13821 16899 13855
rect 17417 13821 17451 13855
rect 18061 13821 18095 13855
rect 5917 13753 5951 13787
rect 7205 13753 7239 13787
rect 6009 13685 6043 13719
rect 6837 13685 6871 13719
rect 7297 13685 7331 13719
rect 1869 13481 1903 13515
rect 5457 13481 5491 13515
rect 6469 13481 6503 13515
rect 10057 13413 10091 13447
rect 1685 13345 1719 13379
rect 2605 13345 2639 13379
rect 5825 13345 5859 13379
rect 6837 13345 6871 13379
rect 10149 13345 10183 13379
rect 11345 13345 11379 13379
rect 2697 13277 2731 13311
rect 2789 13277 2823 13311
rect 5917 13277 5951 13311
rect 6101 13277 6135 13311
rect 6929 13277 6963 13311
rect 7113 13277 7147 13311
rect 10241 13277 10275 13311
rect 11437 13277 11471 13311
rect 11621 13277 11655 13311
rect 2237 13141 2271 13175
rect 9689 13141 9723 13175
rect 10977 13141 11011 13175
rect 6837 12937 6871 12971
rect 4261 12869 4295 12903
rect 6653 12869 6687 12903
rect 2329 12801 2363 12835
rect 3249 12801 3283 12835
rect 4813 12801 4847 12835
rect 6101 12801 6135 12835
rect 2053 12733 2087 12767
rect 3709 12733 3743 12767
rect 5825 12733 5859 12767
rect 3065 12665 3099 12699
rect 4721 12665 4755 12699
rect 7389 12801 7423 12835
rect 8401 12801 8435 12835
rect 9689 12801 9723 12835
rect 11161 12801 11195 12835
rect 13001 12801 13035 12835
rect 14013 12801 14047 12835
rect 14105 12801 14139 12835
rect 9597 12733 9631 12767
rect 10977 12733 11011 12767
rect 8309 12665 8343 12699
rect 12817 12665 12851 12699
rect 12909 12665 12943 12699
rect 1685 12597 1719 12631
rect 2145 12597 2179 12631
rect 2697 12597 2731 12631
rect 3157 12597 3191 12631
rect 4629 12597 4663 12631
rect 5457 12597 5491 12631
rect 5917 12597 5951 12631
rect 6653 12597 6687 12631
rect 7205 12597 7239 12631
rect 7297 12597 7331 12631
rect 7849 12597 7883 12631
rect 8217 12597 8251 12631
rect 9137 12597 9171 12631
rect 9505 12597 9539 12631
rect 10609 12597 10643 12631
rect 11069 12597 11103 12631
rect 12449 12597 12483 12631
rect 13553 12597 13587 12631
rect 13921 12597 13955 12631
rect 1961 12393 1995 12427
rect 2973 12393 3007 12427
rect 6101 12393 6135 12427
rect 9045 12393 9079 12427
rect 8953 12325 8987 12359
rect 2329 12257 2363 12291
rect 3341 12257 3375 12291
rect 4445 12257 4479 12291
rect 6009 12257 6043 12291
rect 7757 12257 7791 12291
rect 7849 12257 7883 12291
rect 10793 12257 10827 12291
rect 11989 12257 12023 12291
rect 13645 12257 13679 12291
rect 2421 12189 2455 12223
rect 2513 12189 2547 12223
rect 3433 12189 3467 12223
rect 3525 12189 3559 12223
rect 4537 12189 4571 12223
rect 4629 12189 4663 12223
rect 6285 12189 6319 12223
rect 7941 12189 7975 12223
rect 9229 12189 9263 12223
rect 9689 12189 9723 12223
rect 10885 12189 10919 12223
rect 10977 12189 11011 12223
rect 12357 12189 12391 12223
rect 13737 12189 13771 12223
rect 13829 12189 13863 12223
rect 17785 12189 17819 12223
rect 5641 12121 5675 12155
rect 4077 12053 4111 12087
rect 7389 12053 7423 12087
rect 8585 12053 8619 12087
rect 10425 12053 10459 12087
rect 13277 12053 13311 12087
rect 3157 11849 3191 11883
rect 6837 11781 6871 11815
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 9045 11713 9079 11747
rect 10057 11713 10091 11747
rect 10517 11713 10551 11747
rect 13553 11713 13587 11747
rect 16221 11713 16255 11747
rect 17233 11713 17267 11747
rect 1777 11645 1811 11679
rect 2044 11645 2078 11679
rect 3433 11645 3467 11679
rect 4169 11645 4203 11679
rect 4436 11645 4470 11679
rect 8861 11645 8895 11679
rect 9873 11645 9907 11679
rect 10784 11645 10818 11679
rect 13277 11645 13311 11679
rect 13921 11645 13955 11679
rect 14177 11645 14211 11679
rect 15945 11645 15979 11679
rect 18061 11645 18095 11679
rect 8953 11577 8987 11611
rect 9965 11577 9999 11611
rect 3617 11509 3651 11543
rect 5549 11509 5583 11543
rect 7205 11509 7239 11543
rect 8493 11509 8527 11543
rect 9505 11509 9539 11543
rect 11897 11509 11931 11543
rect 12909 11509 12943 11543
rect 13369 11509 13403 11543
rect 15301 11509 15335 11543
rect 15577 11509 15611 11543
rect 16037 11509 16071 11543
rect 16589 11509 16623 11543
rect 16957 11509 16991 11543
rect 17049 11509 17083 11543
rect 18245 11509 18279 11543
rect 2789 11305 2823 11339
rect 6929 11305 6963 11339
rect 8861 11305 8895 11339
rect 11069 11305 11103 11339
rect 14289 11305 14323 11339
rect 16681 11305 16715 11339
rect 5356 11237 5390 11271
rect 7849 11237 7883 11271
rect 11713 11237 11747 11271
rect 12900 11237 12934 11271
rect 17224 11237 17258 11271
rect 1676 11169 1710 11203
rect 3065 11169 3099 11203
rect 4445 11169 4479 11203
rect 4537 11169 4571 11203
rect 5089 11169 5123 11203
rect 9945 11169 9979 11203
rect 12633 11169 12667 11203
rect 14933 11169 14967 11203
rect 15557 11169 15591 11203
rect 1409 11101 1443 11135
rect 4721 11101 4755 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 9689 11101 9723 11135
rect 11805 11101 11839 11135
rect 11989 11101 12023 11135
rect 15301 11101 15335 11135
rect 16957 11101 16991 11135
rect 6469 11033 6503 11067
rect 7481 11033 7515 11067
rect 11345 11033 11379 11067
rect 14749 11033 14783 11067
rect 3249 10965 3283 10999
rect 4077 10965 4111 10999
rect 8493 10965 8527 10999
rect 14013 10965 14047 10999
rect 18337 10965 18371 10999
rect 1409 10761 1443 10795
rect 3801 10761 3835 10795
rect 5457 10761 5491 10795
rect 5733 10761 5767 10795
rect 10333 10761 10367 10795
rect 11345 10761 11379 10795
rect 12449 10761 12483 10795
rect 8953 10693 8987 10727
rect 15393 10693 15427 10727
rect 1961 10625 1995 10659
rect 6193 10625 6227 10659
rect 6377 10625 6411 10659
rect 9689 10625 9723 10659
rect 9781 10625 9815 10659
rect 10977 10625 11011 10659
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 13093 10625 13127 10659
rect 14289 10625 14323 10659
rect 15209 10625 15243 10659
rect 15853 10625 15887 10659
rect 16037 10625 16071 10659
rect 2421 10557 2455 10591
rect 2688 10557 2722 10591
rect 4077 10557 4111 10591
rect 4344 10557 4378 10591
rect 7573 10557 7607 10591
rect 7840 10557 7874 10591
rect 9597 10557 9631 10591
rect 14105 10557 14139 10591
rect 14933 10557 14967 10591
rect 16313 10557 16347 10591
rect 18061 10557 18095 10591
rect 1777 10489 1811 10523
rect 6101 10489 6135 10523
rect 10793 10489 10827 10523
rect 12817 10489 12851 10523
rect 14197 10489 14231 10523
rect 15025 10489 15059 10523
rect 16580 10489 16614 10523
rect 1869 10421 1903 10455
rect 9229 10421 9263 10455
rect 10701 10421 10735 10455
rect 11713 10421 11747 10455
rect 12909 10421 12943 10455
rect 13737 10421 13771 10455
rect 14565 10421 14599 10455
rect 15761 10421 15795 10455
rect 17693 10421 17727 10455
rect 18245 10421 18279 10455
rect 1593 10217 1627 10251
rect 2605 10217 2639 10251
rect 5549 10217 5583 10251
rect 6929 10217 6963 10251
rect 11069 10217 11103 10251
rect 12817 10217 12851 10251
rect 13185 10217 13219 10251
rect 13645 10217 13679 10251
rect 14473 10217 14507 10251
rect 15761 10217 15795 10251
rect 16865 10217 16899 10251
rect 17785 10217 17819 10251
rect 2053 10149 2087 10183
rect 4436 10149 4470 10183
rect 7021 10149 7055 10183
rect 7481 10149 7515 10183
rect 14381 10149 14415 10183
rect 15669 10149 15703 10183
rect 1961 10081 1995 10115
rect 2973 10081 3007 10115
rect 3065 10081 3099 10115
rect 3801 10081 3835 10115
rect 2145 10013 2179 10047
rect 3157 10013 3191 10047
rect 4169 10013 4203 10047
rect 5825 10013 5859 10047
rect 7205 10013 7239 10047
rect 7840 10081 7874 10115
rect 9505 10081 9539 10115
rect 9945 10081 9979 10115
rect 11704 10081 11738 10115
rect 13553 10081 13587 10115
rect 16313 10081 16347 10115
rect 17233 10081 17267 10115
rect 7573 10013 7607 10047
rect 9689 10013 9723 10047
rect 11437 10013 11471 10047
rect 13737 10013 13771 10047
rect 14657 10013 14691 10047
rect 15945 10013 15979 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 7389 9945 7423 9979
rect 17877 10081 17911 10115
rect 18061 9945 18095 9979
rect 3617 9877 3651 9911
rect 6561 9877 6595 9911
rect 8953 9877 8987 9911
rect 9321 9877 9355 9911
rect 14013 9877 14047 9911
rect 15301 9877 15335 9911
rect 16497 9877 16531 9911
rect 17785 9877 17819 9911
rect 6469 9673 6503 9707
rect 16957 9673 16991 9707
rect 2053 9605 2087 9639
rect 3065 9605 3099 9639
rect 10241 9605 10275 9639
rect 10333 9605 10367 9639
rect 11161 9605 11195 9639
rect 13829 9605 13863 9639
rect 14105 9605 14139 9639
rect 16313 9605 16347 9639
rect 2605 9537 2639 9571
rect 3709 9537 3743 9571
rect 4537 9537 4571 9571
rect 4721 9537 4755 9571
rect 10885 9537 10919 9571
rect 11621 9537 11655 9571
rect 11805 9537 11839 9571
rect 14933 9537 14967 9571
rect 17417 9537 17451 9571
rect 17601 9537 17635 9571
rect 18981 9537 19015 9571
rect 1501 9469 1535 9503
rect 5089 9469 5123 9503
rect 6653 9469 6687 9503
rect 6837 9469 6871 9503
rect 8677 9469 8711 9503
rect 8769 9469 8803 9503
rect 8861 9469 8895 9503
rect 9128 9469 9162 9503
rect 12449 9469 12483 9503
rect 12705 9469 12739 9503
rect 14289 9469 14323 9503
rect 14381 9469 14415 9503
rect 15200 9469 15234 9503
rect 17325 9469 17359 9503
rect 18061 9469 18095 9503
rect 2421 9401 2455 9435
rect 5356 9401 5390 9435
rect 7082 9401 7116 9435
rect 10793 9401 10827 9435
rect 1685 9333 1719 9367
rect 2513 9333 2547 9367
rect 3433 9333 3467 9367
rect 3525 9333 3559 9367
rect 4077 9333 4111 9367
rect 4445 9333 4479 9367
rect 6653 9333 6687 9367
rect 8217 9333 8251 9367
rect 8493 9333 8527 9367
rect 8769 9333 8803 9367
rect 10701 9333 10735 9367
rect 11529 9333 11563 9367
rect 14565 9333 14599 9367
rect 18245 9333 18279 9367
rect 2789 9129 2823 9163
rect 4813 9129 4847 9163
rect 5181 9129 5215 9163
rect 6193 9129 6227 9163
rect 6285 9129 6319 9163
rect 6837 9129 6871 9163
rect 7573 9129 7607 9163
rect 8125 9129 8159 9163
rect 8585 9129 8619 9163
rect 10333 9129 10367 9163
rect 14565 9129 14599 9163
rect 14657 9129 14691 9163
rect 15025 9129 15059 9163
rect 17417 9129 17451 9163
rect 17785 9129 17819 9163
rect 8953 9061 8987 9095
rect 13553 9061 13587 9095
rect 17877 9061 17911 9095
rect 1676 8993 1710 9027
rect 3065 8993 3099 9027
rect 4077 8993 4111 9027
rect 7021 8993 7055 9027
rect 7481 8993 7515 9027
rect 10701 8993 10735 9027
rect 10793 8993 10827 9027
rect 11612 8993 11646 9027
rect 14013 8993 14047 9027
rect 15025 8993 15059 9027
rect 15761 8993 15795 9027
rect 16028 8993 16062 9027
rect 1409 8925 1443 8959
rect 5273 8925 5307 8959
rect 5365 8925 5399 8959
rect 6377 8925 6411 8959
rect 7757 8925 7791 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 10885 8925 10919 8959
rect 11345 8925 11379 8959
rect 13645 8925 13679 8959
rect 13829 8925 13863 8959
rect 5825 8857 5859 8891
rect 13185 8857 13219 8891
rect 14841 8925 14875 8959
rect 15301 8925 15335 8959
rect 17969 8925 18003 8959
rect 3249 8789 3283 8823
rect 4261 8789 4295 8823
rect 7113 8789 7147 8823
rect 12725 8789 12759 8823
rect 14013 8789 14047 8823
rect 14197 8789 14231 8823
rect 17141 8789 17175 8823
rect 1501 8585 1535 8619
rect 3893 8585 3927 8619
rect 6929 8585 6963 8619
rect 7941 8585 7975 8619
rect 8861 8585 8895 8619
rect 11989 8585 12023 8619
rect 13185 8585 13219 8619
rect 18245 8585 18279 8619
rect 18981 8585 19015 8619
rect 6009 8517 6043 8551
rect 2145 8449 2179 8483
rect 7389 8449 7423 8483
rect 7573 8449 7607 8483
rect 8401 8449 8435 8483
rect 8585 8449 8619 8483
rect 10333 8517 10367 8551
rect 12817 8517 12851 8551
rect 13737 8449 13771 8483
rect 16313 8449 16347 8483
rect 2513 8381 2547 8415
rect 4169 8381 4203 8415
rect 5825 8381 5859 8415
rect 7297 8381 7331 8415
rect 8309 8381 8343 8415
rect 8769 8381 8803 8415
rect 8861 8381 8895 8415
rect 8953 8381 8987 8415
rect 9220 8381 9254 8415
rect 10609 8381 10643 8415
rect 12633 8381 12667 8415
rect 13645 8381 13679 8415
rect 14197 8381 14231 8415
rect 16569 8381 16603 8415
rect 18061 8381 18095 8415
rect 1961 8313 1995 8347
rect 2780 8313 2814 8347
rect 4436 8313 4470 8347
rect 10876 8313 10910 8347
rect 13553 8313 13587 8347
rect 14464 8313 14498 8347
rect 1869 8245 1903 8279
rect 5549 8245 5583 8279
rect 8769 8245 8803 8279
rect 15577 8245 15611 8279
rect 15853 8245 15887 8279
rect 17693 8245 17727 8279
rect 2973 8041 3007 8075
rect 4905 8041 4939 8075
rect 6377 8041 6411 8075
rect 7849 8041 7883 8075
rect 8585 8041 8619 8075
rect 12173 8041 12207 8075
rect 12633 8041 12667 8075
rect 13185 8041 13219 8075
rect 13645 8041 13679 8075
rect 14657 8041 14691 8075
rect 15669 8041 15703 8075
rect 17509 8041 17543 8075
rect 1860 7973 1894 8007
rect 1593 7905 1627 7939
rect 3249 7905 3283 7939
rect 4077 7905 4111 7939
rect 5273 7905 5307 7939
rect 6285 7905 6319 7939
rect 7297 7905 7331 7939
rect 5365 7837 5399 7871
rect 5549 7837 5583 7871
rect 6469 7837 6503 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 9045 7973 9079 8007
rect 14565 7973 14599 8007
rect 15761 7973 15795 8007
rect 16865 7973 16899 8007
rect 17969 7973 18003 8007
rect 7941 7905 7975 7939
rect 8953 7905 8987 7939
rect 9873 7905 9907 7939
rect 12081 7905 12115 7939
rect 12541 7905 12575 7939
rect 13553 7905 13587 7939
rect 17877 7905 17911 7939
rect 9229 7837 9263 7871
rect 12725 7837 12759 7871
rect 13737 7837 13771 7871
rect 14841 7837 14875 7871
rect 15853 7837 15887 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 18061 7837 18095 7871
rect 4261 7769 4295 7803
rect 7849 7769 7883 7803
rect 16497 7769 16531 7803
rect 3433 7701 3467 7735
rect 5917 7701 5951 7735
rect 6929 7701 6963 7735
rect 8125 7701 8159 7735
rect 11161 7701 11195 7735
rect 11897 7701 11931 7735
rect 14197 7701 14231 7735
rect 15301 7701 15335 7735
rect 1685 7497 1719 7531
rect 2697 7497 2731 7531
rect 3709 7497 3743 7531
rect 4721 7497 4755 7531
rect 5549 7497 5583 7531
rect 5733 7497 5767 7531
rect 8217 7497 8251 7531
rect 10517 7497 10551 7531
rect 12449 7497 12483 7531
rect 16497 7497 16531 7531
rect 3617 7429 3651 7463
rect 2145 7361 2179 7395
rect 2329 7361 2363 7395
rect 3341 7361 3375 7395
rect 2053 7225 2087 7259
rect 3065 7225 3099 7259
rect 4169 7361 4203 7395
rect 4261 7361 4295 7395
rect 5181 7361 5215 7395
rect 5365 7361 5399 7395
rect 6377 7361 6411 7395
rect 10977 7361 11011 7395
rect 11161 7361 11195 7395
rect 11897 7361 11931 7395
rect 13001 7361 13035 7395
rect 15761 7361 15795 7395
rect 15853 7361 15887 7395
rect 17141 7361 17175 7395
rect 6837 7293 6871 7327
rect 7093 7293 7127 7327
rect 8493 7293 8527 7327
rect 10885 7293 10919 7327
rect 13652 7293 13686 7327
rect 15669 7293 15703 7327
rect 17509 7293 17543 7327
rect 18061 7293 18095 7327
rect 5089 7225 5123 7259
rect 5549 7225 5583 7259
rect 8738 7225 8772 7259
rect 11713 7225 11747 7259
rect 12909 7225 12943 7259
rect 13912 7225 13946 7259
rect 3157 7157 3191 7191
rect 3617 7157 3651 7191
rect 4077 7157 4111 7191
rect 6101 7157 6135 7191
rect 6193 7157 6227 7191
rect 9873 7157 9907 7191
rect 11345 7157 11379 7191
rect 11805 7157 11839 7191
rect 12817 7157 12851 7191
rect 15025 7157 15059 7191
rect 15301 7157 15335 7191
rect 16865 7157 16899 7191
rect 16957 7157 16991 7191
rect 18245 7157 18279 7191
rect 6653 6953 6687 6987
rect 7113 6953 7147 6987
rect 11713 6953 11747 6987
rect 13737 6953 13771 6987
rect 14565 6953 14599 6987
rect 17049 6953 17083 6987
rect 17693 6953 17727 6987
rect 10701 6885 10735 6919
rect 1685 6817 1719 6851
rect 2504 6817 2538 6851
rect 4629 6817 4663 6851
rect 5273 6817 5307 6851
rect 5540 6817 5574 6851
rect 6929 6817 6963 6851
rect 7665 6817 7699 6851
rect 8116 6817 8150 6851
rect 9689 6817 9723 6851
rect 12613 6817 12647 6851
rect 15669 6817 15703 6851
rect 15925 6817 15959 6851
rect 2237 6749 2271 6783
rect 4721 6749 4755 6783
rect 4905 6749 4939 6783
rect 7849 6749 7883 6783
rect 10793 6749 10827 6783
rect 10977 6749 11011 6783
rect 11805 6749 11839 6783
rect 11989 6749 12023 6783
rect 12357 6749 12391 6783
rect 14657 6749 14691 6783
rect 14841 6749 14875 6783
rect 17785 6749 17819 6783
rect 17877 6749 17911 6783
rect 3617 6681 3651 6715
rect 9873 6681 9907 6715
rect 10333 6681 10367 6715
rect 1869 6613 1903 6647
rect 4261 6613 4295 6647
rect 7481 6613 7515 6647
rect 9229 6613 9263 6647
rect 11345 6613 11379 6647
rect 14197 6613 14231 6647
rect 17325 6613 17359 6647
rect 6101 6409 6135 6443
rect 12081 6409 12115 6443
rect 12449 6409 12483 6443
rect 13645 6341 13679 6375
rect 16037 6341 16071 6375
rect 3709 6273 3743 6307
rect 7665 6273 7699 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 14657 6273 14691 6307
rect 15669 6273 15703 6307
rect 16313 6273 16347 6307
rect 1409 6205 1443 6239
rect 1676 6205 1710 6239
rect 4077 6205 4111 6239
rect 4721 6205 4755 6239
rect 4988 6205 5022 6239
rect 6561 6205 6595 6239
rect 8125 6205 8159 6239
rect 8677 6205 8711 6239
rect 10701 6205 10735 6239
rect 13461 6205 13495 6239
rect 14381 6205 14415 6239
rect 16221 6205 16255 6239
rect 16580 6205 16614 6239
rect 18061 6205 18095 6239
rect 8944 6137 8978 6171
rect 10968 6137 11002 6171
rect 15393 6137 15427 6171
rect 15485 6137 15519 6171
rect 2789 6069 2823 6103
rect 3065 6069 3099 6103
rect 3433 6069 3467 6103
rect 3525 6069 3559 6103
rect 4261 6069 4295 6103
rect 6377 6069 6411 6103
rect 7113 6069 7147 6103
rect 7481 6069 7515 6103
rect 7573 6069 7607 6103
rect 8309 6069 8343 6103
rect 10057 6069 10091 6103
rect 12817 6069 12851 6103
rect 14013 6069 14047 6103
rect 14473 6069 14507 6103
rect 15025 6069 15059 6103
rect 17693 6069 17727 6103
rect 18245 6069 18279 6103
rect 2513 5865 2547 5899
rect 2605 5865 2639 5899
rect 4445 5865 4479 5899
rect 5917 5865 5951 5899
rect 8493 5865 8527 5899
rect 8861 5865 8895 5899
rect 11713 5865 11747 5899
rect 12449 5865 12483 5899
rect 14197 5865 14231 5899
rect 14565 5865 14599 5899
rect 16681 5865 16715 5899
rect 17417 5865 17451 5899
rect 4813 5797 4847 5831
rect 9873 5797 9907 5831
rect 14657 5797 14691 5831
rect 15546 5797 15580 5831
rect 17325 5797 17359 5831
rect 1409 5729 1443 5763
rect 1685 5729 1719 5763
rect 3249 5729 3283 5763
rect 4905 5729 4939 5763
rect 5825 5729 5859 5763
rect 6745 5729 6779 5763
rect 7104 5729 7138 5763
rect 10600 5729 10634 5763
rect 12633 5729 12667 5763
rect 13185 5729 13219 5763
rect 17969 5729 18003 5763
rect 2697 5661 2731 5695
rect 3433 5661 3467 5695
rect 5089 5661 5123 5695
rect 6101 5661 6135 5695
rect 6837 5661 6871 5695
rect 8953 5661 8987 5695
rect 9045 5661 9079 5695
rect 10333 5661 10367 5695
rect 11989 5661 12023 5695
rect 13277 5661 13311 5695
rect 13369 5661 13403 5695
rect 14841 5661 14875 5695
rect 15301 5661 15335 5695
rect 17509 5661 17543 5695
rect 2145 5593 2179 5627
rect 8217 5593 8251 5627
rect 5457 5525 5491 5559
rect 6561 5525 6595 5559
rect 12817 5525 12851 5559
rect 16957 5525 16991 5559
rect 18153 5525 18187 5559
rect 4721 5321 4755 5355
rect 6837 5321 6871 5355
rect 13829 5321 13863 5355
rect 14657 5321 14691 5355
rect 16405 5321 16439 5355
rect 16681 5321 16715 5355
rect 5549 5253 5583 5287
rect 3801 5185 3835 5219
rect 4261 5185 4295 5219
rect 5365 5185 5399 5219
rect 6193 5185 6227 5219
rect 6377 5185 6411 5219
rect 7481 5185 7515 5219
rect 8309 5185 8343 5219
rect 8493 5185 8527 5219
rect 11897 5185 11931 5219
rect 17141 5185 17175 5219
rect 17233 5185 17267 5219
rect 1593 5117 1627 5151
rect 3709 5117 3743 5151
rect 5549 5117 5583 5151
rect 8861 5117 8895 5151
rect 9505 5117 9539 5151
rect 11713 5117 11747 5151
rect 12456 5117 12490 5151
rect 14473 5117 14507 5151
rect 15025 5117 15059 5151
rect 15281 5117 15315 5151
rect 18061 5117 18095 5151
rect 1838 5049 1872 5083
rect 3617 5049 3651 5083
rect 5181 5049 5215 5083
rect 6101 5049 6135 5083
rect 8217 5049 8251 5083
rect 9750 5049 9784 5083
rect 12694 5049 12728 5083
rect 2973 4981 3007 5015
rect 3249 4981 3283 5015
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 7205 4981 7239 5015
rect 7297 4981 7331 5015
rect 7849 4981 7883 5015
rect 9045 4981 9079 5015
rect 10885 4981 10919 5015
rect 11345 4981 11379 5015
rect 11805 4981 11839 5015
rect 17049 4981 17083 5015
rect 18245 4981 18279 5015
rect 4629 4777 4663 4811
rect 8769 4777 8803 4811
rect 10057 4777 10091 4811
rect 10149 4777 10183 4811
rect 11161 4777 11195 4811
rect 11805 4777 11839 4811
rect 12173 4777 12207 4811
rect 12817 4777 12851 4811
rect 13461 4777 13495 4811
rect 15301 4777 15335 4811
rect 16773 4777 16807 4811
rect 17233 4777 17267 4811
rect 17601 4777 17635 4811
rect 2136 4709 2170 4743
rect 5426 4709 5460 4743
rect 11253 4709 11287 4743
rect 13921 4709 13955 4743
rect 15761 4709 15795 4743
rect 3801 4641 3835 4675
rect 4537 4641 4571 4675
rect 6837 4641 6871 4675
rect 7656 4641 7690 4675
rect 9045 4641 9079 4675
rect 13001 4641 13035 4675
rect 13829 4641 13863 4675
rect 14473 4641 14507 4675
rect 15669 4641 15703 4675
rect 17141 4641 17175 4675
rect 1869 4573 1903 4607
rect 4813 4573 4847 4607
rect 5181 4573 5215 4607
rect 7389 4573 7423 4607
rect 10241 4573 10275 4607
rect 11437 4573 11471 4607
rect 12265 4573 12299 4607
rect 12449 4573 12483 4607
rect 14013 4573 14047 4607
rect 15853 4573 15887 4607
rect 17417 4573 17451 4607
rect 3249 4505 3283 4539
rect 10793 4505 10827 4539
rect 17785 4641 17819 4675
rect 18061 4573 18095 4607
rect 3617 4437 3651 4471
rect 4169 4437 4203 4471
rect 6561 4437 6595 4471
rect 7021 4437 7055 4471
rect 9229 4437 9263 4471
rect 9689 4437 9723 4471
rect 17601 4437 17635 4471
rect 8217 4233 8251 4267
rect 11345 4233 11379 4267
rect 14657 4233 14691 4267
rect 16865 4233 16899 4267
rect 4261 4165 4295 4199
rect 14381 4165 14415 4199
rect 2329 4097 2363 4131
rect 2421 4097 2455 4131
rect 2881 4097 2915 4131
rect 5273 4097 5307 4131
rect 6101 4097 6135 4131
rect 6193 4097 6227 4131
rect 11989 4097 12023 4131
rect 13001 4097 13035 4131
rect 15209 4097 15243 4131
rect 2237 4029 2271 4063
rect 3148 4029 3182 4063
rect 4997 4029 5031 4063
rect 5089 4029 5123 4063
rect 6837 4029 6871 4063
rect 8861 4029 8895 4063
rect 10517 4029 10551 4063
rect 11713 4029 11747 4063
rect 11805 4029 11839 4063
rect 13268 4029 13302 4063
rect 15025 4029 15059 4063
rect 16129 4029 16163 4063
rect 16681 4029 16715 4063
rect 17233 4029 17267 4063
rect 18061 4029 18095 4063
rect 6009 3961 6043 3995
rect 7082 3961 7116 3995
rect 9128 3961 9162 3995
rect 10793 3961 10827 3995
rect 15117 3961 15151 3995
rect 1869 3893 1903 3927
rect 4629 3893 4663 3927
rect 5641 3893 5675 3927
rect 10241 3893 10275 3927
rect 12449 3893 12483 3927
rect 16313 3893 16347 3927
rect 17417 3893 17451 3927
rect 18245 3893 18279 3927
rect 2789 3689 2823 3723
rect 5733 3689 5767 3723
rect 7205 3689 7239 3723
rect 7481 3689 7515 3723
rect 7941 3689 7975 3723
rect 8493 3689 8527 3723
rect 8861 3689 8895 3723
rect 9873 3689 9907 3723
rect 13645 3689 13679 3723
rect 14013 3689 14047 3723
rect 5181 3621 5215 3655
rect 1665 3553 1699 3587
rect 3249 3553 3283 3587
rect 4077 3553 4111 3587
rect 1409 3485 1443 3519
rect 3525 3485 3559 3519
rect 4353 3485 4387 3519
rect 5273 3485 5307 3519
rect 5365 3485 5399 3519
rect 10578 3621 10612 3655
rect 6081 3553 6115 3587
rect 7849 3553 7883 3587
rect 8953 3553 8987 3587
rect 9689 3553 9723 3587
rect 10333 3553 10367 3587
rect 12245 3553 12279 3587
rect 16497 3553 16531 3587
rect 17049 3553 17083 3587
rect 17785 3553 17819 3587
rect 5825 3485 5859 3519
rect 8125 3485 8159 3519
rect 9045 3485 9079 3519
rect 11989 3485 12023 3519
rect 14105 3485 14139 3519
rect 14197 3485 14231 3519
rect 17233 3485 17267 3519
rect 18061 3485 18095 3519
rect 16681 3417 16715 3451
rect 4813 3349 4847 3383
rect 5733 3349 5767 3383
rect 11713 3349 11747 3383
rect 13369 3349 13403 3383
rect 1777 3145 1811 3179
rect 3801 3145 3835 3179
rect 9689 3145 9723 3179
rect 18245 3145 18279 3179
rect 2605 3077 2639 3111
rect 2789 3077 2823 3111
rect 8677 3077 8711 3111
rect 16313 3077 16347 3111
rect 2237 3009 2271 3043
rect 2421 3009 2455 3043
rect 3433 3009 3467 3043
rect 4261 3009 4295 3043
rect 4445 3009 4479 3043
rect 5365 3009 5399 3043
rect 9229 3009 9263 3043
rect 10241 3009 10275 3043
rect 11253 3009 11287 3043
rect 13001 3009 13035 3043
rect 3249 2941 3283 2975
rect 6009 2941 6043 2975
rect 7205 2941 7239 2975
rect 7941 2941 7975 2975
rect 9045 2941 9079 2975
rect 11713 2941 11747 2975
rect 13461 2941 13495 2975
rect 14197 2941 14231 2975
rect 14933 2941 14967 2975
rect 16497 2941 16531 2975
rect 17233 2941 17267 2975
rect 18061 2941 18095 2975
rect 2145 2873 2179 2907
rect 2605 2873 2639 2907
rect 3157 2873 3191 2907
rect 5181 2873 5215 2907
rect 6285 2873 6319 2907
rect 7481 2873 7515 2907
rect 8217 2873 8251 2907
rect 9137 2873 9171 2907
rect 10057 2873 10091 2907
rect 11161 2873 11195 2907
rect 12817 2873 12851 2907
rect 13737 2873 13771 2907
rect 14473 2873 14507 2907
rect 15209 2873 15243 2907
rect 16773 2873 16807 2907
rect 17509 2873 17543 2907
rect 4169 2805 4203 2839
rect 4813 2805 4847 2839
rect 5273 2805 5307 2839
rect 10149 2805 10183 2839
rect 10701 2805 10735 2839
rect 11069 2805 11103 2839
rect 11897 2805 11931 2839
rect 12449 2805 12483 2839
rect 12909 2805 12943 2839
rect 1593 2601 1627 2635
rect 1961 2601 1995 2635
rect 2421 2601 2455 2635
rect 2973 2601 3007 2635
rect 3341 2601 3375 2635
rect 4353 2601 4387 2635
rect 4721 2601 4755 2635
rect 5365 2601 5399 2635
rect 5733 2601 5767 2635
rect 6377 2601 6411 2635
rect 8677 2601 8711 2635
rect 10149 2601 10183 2635
rect 10793 2601 10827 2635
rect 11253 2601 11287 2635
rect 16681 2601 16715 2635
rect 2329 2533 2363 2567
rect 5825 2533 5859 2567
rect 10241 2533 10275 2567
rect 1409 2465 1443 2499
rect 3433 2465 3467 2499
rect 4813 2465 4847 2499
rect 6929 2465 6963 2499
rect 7941 2465 7975 2499
rect 9045 2465 9079 2499
rect 11161 2465 11195 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 14381 2465 14415 2499
rect 16773 2465 16807 2499
rect 17509 2465 17543 2499
rect 2605 2397 2639 2431
rect 3525 2397 3559 2431
rect 4997 2397 5031 2431
rect 5917 2397 5951 2431
rect 7113 2397 7147 2431
rect 8217 2397 8251 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 11345 2397 11379 2431
rect 11989 2397 12023 2431
rect 12817 2397 12851 2431
rect 14565 2397 14599 2431
rect 17049 2397 17083 2431
rect 17785 2397 17819 2431
rect 9781 2329 9815 2363
rect 17325 2329 17359 2363
<< metal1 >>
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 6454 16572 6460 16584
rect 3384 16544 6460 16572
rect 3384 16532 3390 16544
rect 6454 16532 6460 16544
rect 6512 16532 6518 16584
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 3418 14600 3424 14612
rect 3379 14572 3424 14600
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5040 14572 5457 14600
rect 5040 14560 5046 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 6454 14600 6460 14612
rect 6415 14572 6460 14600
rect 5445 14563 5503 14569
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 2038 14532 2044 14544
rect 1999 14504 2044 14532
rect 2038 14492 2044 14504
rect 2096 14492 2102 14544
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 2832 14504 2877 14532
rect 2832 14492 2838 14504
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14464 2559 14467
rect 3237 14467 3295 14473
rect 3237 14464 3249 14467
rect 2547 14436 3249 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 3237 14433 3249 14436
rect 3283 14464 3295 14467
rect 3326 14464 3332 14476
rect 3283 14436 3332 14464
rect 3283 14433 3295 14436
rect 3237 14427 3295 14433
rect 1780 14396 1808 14427
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 5166 14424 5172 14476
rect 5224 14464 5230 14476
rect 5261 14467 5319 14473
rect 5261 14464 5273 14467
rect 5224 14436 5273 14464
rect 5224 14424 5230 14436
rect 5261 14433 5273 14436
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 8018 14464 8024 14476
rect 6319 14436 8024 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 3602 14396 3608 14408
rect 1780 14368 3608 14396
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 17586 14328 17592 14340
rect 4120 14300 17592 14328
rect 4120 14288 4126 14300
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 17586 14056 17592 14068
rect 1728 14028 16712 14056
rect 17547 14028 17592 14056
rect 1728 14016 1734 14028
rect 3234 13988 3240 14000
rect 3195 13960 3240 13988
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 3786 13988 3792 14000
rect 3747 13960 3792 13988
rect 3786 13948 3792 13960
rect 3844 13948 3850 14000
rect 5537 13991 5595 13997
rect 5537 13957 5549 13991
rect 5583 13988 5595 13991
rect 5626 13988 5632 14000
rect 5583 13960 5632 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2774 13920 2780 13932
rect 2639 13892 2780 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 6089 13923 6147 13929
rect 6089 13920 6101 13923
rect 5500 13892 6101 13920
rect 5500 13880 5506 13892
rect 6089 13889 6101 13892
rect 6135 13889 6147 13923
rect 6089 13883 6147 13889
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 6328 13892 7389 13920
rect 6328 13880 6334 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 8294 13920 8300 13932
rect 8255 13892 8300 13920
rect 7377 13883 7435 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 14918 13920 14924 13932
rect 14507 13892 14924 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 16684 13920 16712 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 18230 14056 18236 14068
rect 18191 14028 18236 14056
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 16758 13948 16764 14000
rect 16816 13988 16822 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16816 13960 17049 13988
rect 16816 13948 16822 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 16684 13892 16896 13920
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13821 1639 13855
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1581 13815 1639 13821
rect 1596 13784 1624 13815
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 3050 13852 3056 13864
rect 2363 13824 3056 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3602 13852 3608 13864
rect 3563 13824 3608 13852
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 8018 13852 8024 13864
rect 7979 13824 8024 13852
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 16868 13861 16896 13892
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 11664 13824 14197 13852
rect 11664 13812 11670 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13821 16911 13855
rect 17402 13852 17408 13864
rect 17363 13824 17408 13852
rect 16853 13815 16911 13821
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17920 13824 18061 13852
rect 17920 13812 17926 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 1762 13784 1768 13796
rect 1596 13756 1768 13784
rect 1762 13744 1768 13756
rect 1820 13744 1826 13796
rect 5905 13787 5963 13793
rect 5905 13753 5917 13787
rect 5951 13784 5963 13787
rect 7193 13787 7251 13793
rect 5951 13756 6868 13784
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 5994 13716 6000 13728
rect 5955 13688 6000 13716
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 6840 13725 6868 13756
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 7374 13784 7380 13796
rect 7239 13756 7380 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13685 6883 13719
rect 7282 13716 7288 13728
rect 7243 13688 7288 13716
rect 6825 13679 6883 13685
rect 7282 13676 7288 13688
rect 7340 13676 7346 13728
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1857 13515 1915 13521
rect 1857 13481 1869 13515
rect 1903 13512 1915 13515
rect 2866 13512 2872 13524
rect 1903 13484 2872 13512
rect 1903 13481 1915 13484
rect 1857 13475 1915 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5994 13512 6000 13524
rect 5491 13484 6000 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 7282 13512 7288 13524
rect 6503 13484 7288 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 11882 13512 11888 13524
rect 7524 13484 11888 13512
rect 7524 13472 7530 13484
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 10045 13447 10103 13453
rect 10045 13444 10057 13447
rect 9824 13416 10057 13444
rect 9824 13404 9830 13416
rect 10045 13413 10057 13416
rect 10091 13444 10103 13447
rect 15194 13444 15200 13456
rect 10091 13416 15200 13444
rect 10091 13413 10103 13416
rect 10045 13407 10103 13413
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 1762 13376 1768 13388
rect 1719 13348 1768 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 5258 13376 5264 13388
rect 3384 13348 5264 13376
rect 3384 13336 3390 13348
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5810 13376 5816 13388
rect 5771 13348 5816 13376
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6472 13348 6837 13376
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 1452 13280 2697 13308
rect 1452 13268 1458 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13277 2835 13311
rect 5902 13308 5908 13320
rect 5863 13280 5908 13308
rect 2777 13271 2835 13277
rect 2498 13200 2504 13252
rect 2556 13240 2562 13252
rect 2792 13240 2820 13271
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 6086 13308 6092 13320
rect 5999 13280 6092 13308
rect 6086 13268 6092 13280
rect 6144 13308 6150 13320
rect 6270 13308 6276 13320
rect 6144 13280 6276 13308
rect 6144 13268 6150 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 2556 13212 2820 13240
rect 2556 13200 2562 13212
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 2225 13175 2283 13181
rect 2225 13172 2237 13175
rect 2096 13144 2237 13172
rect 2096 13132 2102 13144
rect 2225 13141 2237 13144
rect 2271 13141 2283 13175
rect 2225 13135 2283 13141
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 6472 13172 6500 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 11146 13376 11152 13388
rect 10183 13348 11152 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11256 13348 11345 13376
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6604 13280 6929 13308
rect 6604 13268 6610 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 7098 13308 7104 13320
rect 7059 13280 7104 13308
rect 6917 13271 6975 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10284 13280 10329 13308
rect 10284 13268 10290 13280
rect 7742 13200 7748 13252
rect 7800 13240 7806 13252
rect 11256 13240 11284 13348
rect 11333 13345 11345 13348
rect 11379 13376 11391 13379
rect 14642 13376 14648 13388
rect 11379 13348 14648 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 11422 13308 11428 13320
rect 11383 13280 11428 13308
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 7800 13212 11284 13240
rect 7800 13200 7806 13212
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 15286 13240 15292 13252
rect 11848 13212 15292 13240
rect 11848 13200 11854 13212
rect 15286 13200 15292 13212
rect 15344 13200 15350 13252
rect 7558 13172 7564 13184
rect 3844 13144 7564 13172
rect 3844 13132 3850 13144
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 9674 13172 9680 13184
rect 9635 13144 9680 13172
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 10962 13172 10968 13184
rect 10923 13144 10968 13172
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 4706 12968 4712 12980
rect 3016 12940 4712 12968
rect 3016 12928 3022 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5810 12928 5816 12980
rect 5868 12968 5874 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 5868 12940 6837 12968
rect 5868 12928 5874 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 7466 12968 7472 12980
rect 6825 12931 6883 12937
rect 6932 12940 7472 12968
rect 4249 12903 4307 12909
rect 4249 12869 4261 12903
rect 4295 12900 4307 12903
rect 5534 12900 5540 12912
rect 4295 12872 5540 12900
rect 4295 12869 4307 12872
rect 4249 12863 4307 12869
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 5994 12860 6000 12912
rect 6052 12900 6058 12912
rect 6641 12903 6699 12909
rect 6052 12872 6132 12900
rect 6052 12860 6058 12872
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2682 12832 2688 12844
rect 2363 12804 2688 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3050 12792 3056 12844
rect 3108 12832 3114 12844
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 3108 12804 3249 12832
rect 3108 12792 3114 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 4614 12832 4620 12844
rect 3237 12795 3295 12801
rect 4264 12804 4620 12832
rect 2038 12764 2044 12776
rect 1999 12736 2044 12764
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 2406 12724 2412 12776
rect 2464 12764 2470 12776
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 2464 12736 3709 12764
rect 2464 12724 2470 12736
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 1486 12656 1492 12708
rect 1544 12696 1550 12708
rect 3053 12699 3111 12705
rect 1544 12668 2728 12696
rect 1544 12656 1550 12668
rect 1673 12631 1731 12637
rect 1673 12597 1685 12631
rect 1719 12628 1731 12631
rect 1854 12628 1860 12640
rect 1719 12600 1860 12628
rect 1719 12597 1731 12600
rect 1673 12591 1731 12597
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 2130 12588 2136 12640
rect 2188 12628 2194 12640
rect 2700 12637 2728 12668
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 4264 12696 4292 12804
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 4798 12832 4804 12844
rect 4759 12804 4804 12832
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 6104 12841 6132 12872
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 6932 12900 6960 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 16482 12968 16488 12980
rect 12860 12940 16488 12968
rect 12860 12928 12866 12940
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 6687 12872 6960 12900
rect 7024 12872 9812 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12801 6147 12835
rect 6089 12795 6147 12801
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 5813 12767 5871 12773
rect 5813 12764 5825 12767
rect 4396 12736 5825 12764
rect 4396 12724 4402 12736
rect 5813 12733 5825 12736
rect 5859 12733 5871 12767
rect 5813 12727 5871 12733
rect 3099 12668 4292 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 4522 12656 4528 12708
rect 4580 12696 4586 12708
rect 4709 12699 4767 12705
rect 4709 12696 4721 12699
rect 4580 12668 4721 12696
rect 4580 12656 4586 12668
rect 4709 12665 4721 12668
rect 4755 12665 4767 12699
rect 7024 12696 7052 12872
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7156 12804 7389 12832
rect 7156 12792 7162 12804
rect 7377 12801 7389 12804
rect 7423 12832 7435 12835
rect 7466 12832 7472 12844
rect 7423 12804 7472 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7466 12792 7472 12804
rect 7524 12832 7530 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 7524 12804 8401 12832
rect 7524 12792 7530 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 9677 12835 9735 12841
rect 9677 12832 9689 12835
rect 9364 12804 9689 12832
rect 9364 12792 9370 12804
rect 9677 12801 9689 12804
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 7926 12724 7932 12776
rect 7984 12764 7990 12776
rect 9585 12767 9643 12773
rect 9585 12764 9597 12767
rect 7984 12736 9597 12764
rect 7984 12724 7990 12736
rect 9585 12733 9597 12736
rect 9631 12733 9643 12767
rect 9585 12727 9643 12733
rect 4709 12659 4767 12665
rect 5368 12668 7052 12696
rect 2685 12631 2743 12637
rect 2188 12600 2233 12628
rect 2188 12588 2194 12600
rect 2685 12597 2697 12631
rect 2731 12597 2743 12631
rect 2685 12591 2743 12597
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 4617 12631 4675 12637
rect 3200 12600 3245 12628
rect 3200 12588 3206 12600
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 5368 12628 5396 12668
rect 7374 12656 7380 12708
rect 7432 12696 7438 12708
rect 7432 12668 7880 12696
rect 7432 12656 7438 12668
rect 4663 12600 5396 12628
rect 5445 12631 5503 12637
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 5445 12597 5457 12631
rect 5491 12628 5503 12631
rect 5718 12628 5724 12640
rect 5491 12600 5724 12628
rect 5491 12597 5503 12600
rect 5445 12591 5503 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5868 12600 5917 12628
rect 5868 12588 5874 12600
rect 5905 12597 5917 12600
rect 5951 12628 5963 12631
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 5951 12600 6653 12628
rect 5951 12597 5963 12600
rect 5905 12591 5963 12597
rect 6641 12597 6653 12600
rect 6687 12597 6699 12631
rect 6641 12591 6699 12597
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 6788 12600 7205 12628
rect 6788 12588 6794 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 7285 12631 7343 12637
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7742 12628 7748 12640
rect 7331 12600 7748 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 7852 12637 7880 12668
rect 8018 12656 8024 12708
rect 8076 12696 8082 12708
rect 8297 12699 8355 12705
rect 8297 12696 8309 12699
rect 8076 12668 8309 12696
rect 8076 12656 8082 12668
rect 8297 12665 8309 12668
rect 8343 12665 8355 12699
rect 9784 12696 9812 12872
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 11790 12900 11796 12912
rect 10744 12872 11796 12900
rect 10744 12860 10750 12872
rect 11790 12860 11796 12872
rect 11848 12860 11854 12912
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 11940 12872 14044 12900
rect 11940 12860 11946 12872
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 10928 12804 11161 12832
rect 10928 12792 10934 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 14016 12841 14044 12872
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 11664 12804 13001 12832
rect 11664 12792 11670 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 10962 12764 10968 12776
rect 10923 12736 10968 12764
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 14108 12764 14136 12795
rect 12400 12736 14136 12764
rect 12400 12724 12406 12736
rect 12802 12696 12808 12708
rect 9784 12668 12808 12696
rect 8297 12659 8355 12665
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 12897 12699 12955 12705
rect 12897 12665 12909 12699
rect 12943 12696 12955 12699
rect 17034 12696 17040 12708
rect 12943 12668 17040 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 7837 12631 7895 12637
rect 7837 12597 7849 12631
rect 7883 12597 7895 12631
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 7837 12591 7895 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 8720 12600 9137 12628
rect 8720 12588 8726 12600
rect 9125 12597 9137 12600
rect 9171 12597 9183 12631
rect 9125 12591 9183 12597
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9272 12600 9505 12628
rect 9272 12588 9278 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 10594 12628 10600 12640
rect 10555 12600 10600 12628
rect 9493 12591 9551 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 12437 12631 12495 12637
rect 12437 12628 12449 12631
rect 11103 12600 12449 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 12437 12597 12449 12600
rect 12483 12597 12495 12631
rect 13538 12628 13544 12640
rect 13499 12600 13544 12628
rect 12437 12591 12495 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12628 13967 12631
rect 15010 12628 15016 12640
rect 13955 12600 15016 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2130 12424 2136 12436
rect 1995 12396 2136 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 3142 12424 3148 12436
rect 3007 12396 3148 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 4890 12424 4896 12436
rect 4580 12396 4896 12424
rect 4580 12384 4586 12396
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6089 12427 6147 12433
rect 6089 12424 6101 12427
rect 5776 12396 6101 12424
rect 5776 12384 5782 12396
rect 6089 12393 6101 12396
rect 6135 12393 6147 12427
rect 6089 12387 6147 12393
rect 9033 12427 9091 12433
rect 9033 12393 9045 12427
rect 9079 12424 9091 12427
rect 9674 12424 9680 12436
rect 9079 12396 9680 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15194 12424 15200 12436
rect 14792 12396 15200 12424
rect 14792 12384 14798 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 3476 12328 8953 12356
rect 3476 12316 3482 12328
rect 8941 12325 8953 12328
rect 8987 12356 8999 12359
rect 11514 12356 11520 12368
rect 8987 12328 11520 12356
rect 8987 12325 8999 12328
rect 8941 12319 8999 12325
rect 11514 12316 11520 12328
rect 11572 12316 11578 12368
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2317 12291 2375 12297
rect 2317 12288 2329 12291
rect 2096 12260 2329 12288
rect 2096 12248 2102 12260
rect 2317 12257 2329 12260
rect 2363 12257 2375 12291
rect 3326 12288 3332 12300
rect 3287 12260 3332 12288
rect 2317 12251 2375 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 4430 12288 4436 12300
rect 4391 12260 4436 12288
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 6638 12288 6644 12300
rect 6043 12260 6644 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7708 12260 7757 12288
rect 7708 12248 7714 12260
rect 7745 12257 7757 12260
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 7883 12260 8984 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 8956 12232 8984 12260
rect 10502 12248 10508 12300
rect 10560 12288 10566 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10560 12260 10793 12288
rect 10560 12248 10566 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11664 12260 11989 12288
rect 11664 12248 11670 12260
rect 11977 12257 11989 12260
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 14274 12288 14280 12300
rect 13679 12260 14280 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 2556 12192 2601 12220
rect 2556 12180 2562 12192
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 2832 12192 3433 12220
rect 2832 12180 2838 12192
rect 3421 12189 3433 12192
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12189 3571 12223
rect 4522 12220 4528 12232
rect 4483 12192 4528 12220
rect 3513 12183 3571 12189
rect 2222 12112 2228 12164
rect 2280 12152 2286 12164
rect 3528 12152 3556 12183
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12220 6331 12223
rect 6362 12220 6368 12232
rect 6319 12192 6368 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 2280 12124 3556 12152
rect 2280 12112 2286 12124
rect 3786 12112 3792 12164
rect 3844 12152 3850 12164
rect 4632 12152 4660 12183
rect 6362 12180 6368 12192
rect 6420 12220 6426 12232
rect 7929 12223 7987 12229
rect 6420 12192 7420 12220
rect 6420 12180 6426 12192
rect 3844 12124 4660 12152
rect 5629 12155 5687 12161
rect 3844 12112 3850 12124
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 7282 12152 7288 12164
rect 5675 12124 7288 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 7392 12152 7420 12192
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 7944 12152 7972 12183
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12220 9275 12223
rect 9306 12220 9312 12232
rect 9263 12192 9312 12220
rect 9263 12189 9275 12192
rect 9217 12183 9275 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9456 12192 9689 12220
rect 9456 12180 9462 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 10870 12220 10876 12232
rect 10831 12192 10876 12220
rect 9677 12183 9735 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 12345 12223 12403 12229
rect 11020 12192 11065 12220
rect 11020 12180 11026 12192
rect 12345 12189 12357 12223
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 7392 12124 7972 12152
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 8812 12124 10732 12152
rect 8812 12112 8818 12124
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3660 12056 4077 12084
rect 3660 12044 3666 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 6512 12056 7389 12084
rect 6512 12044 6518 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8168 12056 8585 12084
rect 8168 12044 8174 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 8573 12047 8631 12053
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 10376 12056 10425 12084
rect 10376 12044 10382 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10704 12084 10732 12124
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 12360 12152 12388 12183
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 12768 12192 13737 12220
rect 12768 12180 12774 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13740 12152 13768 12183
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 17770 12220 17776 12232
rect 13872 12192 13917 12220
rect 17731 12192 17776 12220
rect 13872 12180 13878 12192
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 15562 12152 15568 12164
rect 10836 12124 12388 12152
rect 13096 12124 13676 12152
rect 13740 12124 15568 12152
rect 10836 12112 10842 12124
rect 11422 12084 11428 12096
rect 10704 12056 11428 12084
rect 10413 12047 10471 12053
rect 11422 12044 11428 12056
rect 11480 12084 11486 12096
rect 11882 12084 11888 12096
rect 11480 12056 11888 12084
rect 11480 12044 11486 12056
rect 11882 12044 11888 12056
rect 11940 12084 11946 12096
rect 13096 12084 13124 12124
rect 13262 12084 13268 12096
rect 11940 12056 13124 12084
rect 13223 12056 13268 12084
rect 11940 12044 11946 12056
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 13648 12084 13676 12124
rect 15562 12112 15568 12124
rect 15620 12112 15626 12164
rect 15102 12084 15108 12096
rect 13648 12056 15108 12084
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2740 11852 3157 11880
rect 2740 11840 2746 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 3694 11840 3700 11892
rect 3752 11880 3758 11892
rect 3752 11852 11560 11880
rect 3752 11840 3758 11852
rect 5902 11772 5908 11824
rect 5960 11812 5966 11824
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 5960 11784 6837 11812
rect 5960 11772 5966 11784
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 6825 11775 6883 11781
rect 9674 11772 9680 11824
rect 9732 11812 9738 11824
rect 11532 11812 11560 11852
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 16114 11880 16120 11892
rect 11664 11852 16120 11880
rect 11664 11840 11670 11852
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 13170 11812 13176 11824
rect 9732 11784 10548 11812
rect 11532 11784 13176 11812
rect 9732 11772 9738 11784
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 5592 11716 7297 11744
rect 5592 11704 5598 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7466 11744 7472 11756
rect 7427 11716 7472 11744
rect 7285 11707 7343 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8628 11716 9045 11744
rect 8628 11704 8634 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 10520 11753 10548 11784
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 9180 11716 10057 11744
rect 9180 11704 9186 11716
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 16209 11747 16267 11753
rect 13587 11716 14044 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 1765 11679 1823 11685
rect 1765 11676 1777 11679
rect 1636 11648 1777 11676
rect 1636 11636 1642 11648
rect 1765 11645 1777 11648
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 2032 11679 2090 11685
rect 2032 11645 2044 11679
rect 2078 11676 2090 11679
rect 2498 11676 2504 11688
rect 2078 11648 2504 11676
rect 2078 11645 2090 11648
rect 2032 11639 2090 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 4157 11679 4215 11685
rect 3467 11648 3740 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3605 11543 3663 11549
rect 3605 11540 3617 11543
rect 3016 11512 3617 11540
rect 3016 11500 3022 11512
rect 3605 11509 3617 11512
rect 3651 11509 3663 11543
rect 3712 11540 3740 11648
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4172 11608 4200 11639
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4424 11679 4482 11685
rect 4424 11676 4436 11679
rect 4304 11648 4436 11676
rect 4304 11636 4310 11648
rect 4424 11645 4436 11648
rect 4470 11676 4482 11679
rect 4798 11676 4804 11688
rect 4470 11648 4804 11676
rect 4470 11645 4482 11648
rect 4424 11639 4482 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 6270 11676 6276 11688
rect 4908 11648 6276 11676
rect 4338 11608 4344 11620
rect 4172 11580 4344 11608
rect 4338 11568 4344 11580
rect 4396 11568 4402 11620
rect 4908 11540 4936 11648
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 7484 11608 7512 11704
rect 14016 11688 14044 11716
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16574 11744 16580 11756
rect 16255 11716 16580 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 17218 11744 17224 11756
rect 17179 11716 17224 11744
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 8754 11676 8760 11688
rect 5552 11580 7512 11608
rect 7576 11648 8760 11676
rect 5552 11552 5580 11580
rect 5534 11540 5540 11552
rect 3712 11512 4936 11540
rect 5447 11512 5540 11540
rect 3605 11503 3663 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 5868 11512 7205 11540
rect 5868 11500 5874 11512
rect 7193 11509 7205 11512
rect 7239 11540 7251 11543
rect 7576 11540 7604 11648
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 9398 11676 9404 11688
rect 8895 11648 9404 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11676 9919 11679
rect 10318 11676 10324 11688
rect 9907 11648 10324 11676
rect 9907 11645 9919 11648
rect 9861 11639 9919 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 10772 11679 10830 11685
rect 10772 11645 10784 11679
rect 10818 11676 10830 11679
rect 11054 11676 11060 11688
rect 10818 11648 11060 11676
rect 10818 11645 10830 11648
rect 10772 11639 10830 11645
rect 11054 11636 11060 11648
rect 11112 11676 11118 11688
rect 11698 11676 11704 11688
rect 11112 11648 11704 11676
rect 11112 11636 11118 11648
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 13262 11676 13268 11688
rect 13223 11648 13268 11676
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13906 11676 13912 11688
rect 13867 11648 13912 11676
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14165 11679 14223 11685
rect 14165 11676 14177 11679
rect 14056 11648 14177 11676
rect 14056 11636 14062 11648
rect 14165 11645 14177 11648
rect 14211 11645 14223 11679
rect 14165 11639 14223 11645
rect 15102 11636 15108 11688
rect 15160 11676 15166 11688
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 15160 11648 15945 11676
rect 15160 11636 15166 11648
rect 15933 11645 15945 11648
rect 15979 11676 15991 11679
rect 17126 11676 17132 11688
rect 15979 11648 17132 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 8018 11608 8024 11620
rect 7708 11580 8024 11608
rect 7708 11568 7714 11580
rect 8018 11568 8024 11580
rect 8076 11608 8082 11620
rect 8941 11611 8999 11617
rect 8941 11608 8953 11611
rect 8076 11580 8953 11608
rect 8076 11568 8082 11580
rect 8941 11577 8953 11580
rect 8987 11608 8999 11611
rect 9953 11611 10011 11617
rect 8987 11580 9904 11608
rect 8987 11577 8999 11580
rect 8941 11571 8999 11577
rect 9876 11552 9904 11580
rect 9953 11577 9965 11611
rect 9999 11608 10011 11611
rect 10594 11608 10600 11620
rect 9999 11580 10600 11608
rect 9999 11577 10011 11580
rect 9953 11571 10011 11577
rect 10594 11568 10600 11580
rect 10652 11568 10658 11620
rect 14366 11608 14372 11620
rect 12912 11580 14372 11608
rect 7239 11512 7604 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8294 11540 8300 11552
rect 7892 11512 8300 11540
rect 7892 11500 7898 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8481 11543 8539 11549
rect 8481 11509 8493 11543
rect 8527 11540 8539 11543
rect 8846 11540 8852 11552
rect 8527 11512 8852 11540
rect 8527 11509 8539 11512
rect 8481 11503 8539 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9490 11540 9496 11552
rect 9451 11512 9496 11540
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 9858 11500 9864 11552
rect 9916 11500 9922 11552
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 12912 11549 12940 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11020 11512 11897 11540
rect 11020 11500 11026 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 11885 11503 11943 11509
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11509 12955 11543
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 12897 11503 12955 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15010 11540 15016 11552
rect 14884 11512 15016 11540
rect 14884 11500 14890 11512
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15289 11543 15347 11549
rect 15289 11540 15301 11543
rect 15160 11512 15301 11540
rect 15160 11500 15166 11512
rect 15289 11509 15301 11512
rect 15335 11509 15347 11543
rect 15562 11540 15568 11552
rect 15523 11512 15568 11540
rect 15289 11503 15347 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16577 11543 16635 11549
rect 16577 11540 16589 11543
rect 16071 11512 16589 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16577 11509 16589 11512
rect 16623 11509 16635 11543
rect 16577 11503 16635 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16724 11512 16957 11540
rect 16724 11500 16730 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17494 11540 17500 11552
rect 17092 11512 17500 11540
rect 17092 11500 17098 11512
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 18414 11540 18420 11552
rect 18279 11512 18420 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2556 11308 2789 11336
rect 2556 11296 2562 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 6917 11339 6975 11345
rect 2777 11299 2835 11305
rect 3068 11308 6868 11336
rect 1664 11203 1722 11209
rect 1664 11169 1676 11203
rect 1710 11200 1722 11203
rect 1946 11200 1952 11212
rect 1710 11172 1952 11200
rect 1710 11169 1722 11172
rect 1664 11163 1722 11169
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 3068 11209 3096 11308
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 5344 11271 5402 11277
rect 4396 11240 5120 11268
rect 4396 11228 4402 11240
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 5092 11209 5120 11240
rect 5344 11237 5356 11271
rect 5390 11268 5402 11271
rect 5534 11268 5540 11280
rect 5390 11240 5540 11268
rect 5390 11237 5402 11240
rect 5344 11231 5402 11237
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 5902 11228 5908 11280
rect 5960 11268 5966 11280
rect 6086 11268 6092 11280
rect 5960 11240 6092 11268
rect 5960 11228 5966 11240
rect 6086 11228 6092 11240
rect 6144 11268 6150 11280
rect 6840 11268 6868 11308
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 8202 11336 8208 11348
rect 6963 11308 8208 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 9180 11308 11069 11336
rect 9180 11296 9186 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 14274 11336 14280 11348
rect 11057 11299 11115 11305
rect 11164 11308 13952 11336
rect 14235 11308 14280 11336
rect 7650 11268 7656 11280
rect 6144 11240 6316 11268
rect 6840 11240 7656 11268
rect 6144 11228 6150 11240
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 5077 11203 5135 11209
rect 4571 11172 5028 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 5000 11132 5028 11172
rect 5077 11169 5089 11203
rect 5123 11169 5135 11203
rect 5718 11200 5724 11212
rect 5077 11163 5135 11169
rect 5184 11172 5724 11200
rect 5184 11132 5212 11172
rect 5718 11160 5724 11172
rect 5776 11200 5782 11212
rect 5776 11172 6132 11200
rect 5776 11160 5782 11172
rect 6104 11144 6132 11172
rect 5000 11104 5212 11132
rect 4709 11095 4767 11101
rect 1412 10996 1440 11095
rect 4154 11024 4160 11076
rect 4212 11024 4218 11076
rect 4724 11064 4752 11095
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 4982 11064 4988 11076
rect 4724 11036 4988 11064
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 6288 11064 6316 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 7800 11240 7849 11268
rect 7800 11228 7806 11240
rect 7837 11237 7849 11240
rect 7883 11268 7895 11271
rect 11164 11268 11192 11308
rect 7883 11240 11192 11268
rect 7883 11237 7895 11240
rect 7837 11231 7895 11237
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 11698 11268 11704 11280
rect 11572 11240 11704 11268
rect 11572 11228 11578 11240
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12888 11271 12946 11277
rect 12888 11268 12900 11271
rect 11992 11240 12900 11268
rect 9933 11203 9991 11209
rect 9933 11200 9945 11203
rect 8588 11172 9945 11200
rect 8588 11144 8616 11172
rect 9933 11169 9945 11172
rect 9979 11200 9991 11203
rect 10962 11200 10968 11212
rect 9979 11172 10968 11200
rect 9979 11169 9991 11172
rect 9933 11163 9991 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7892 11104 7941 11132
rect 7892 11092 7898 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8570 11132 8576 11144
rect 8159 11104 8576 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8941 11095 8999 11101
rect 9048 11104 9137 11132
rect 6457 11067 6515 11073
rect 6457 11064 6469 11067
rect 6288 11036 6469 11064
rect 6457 11033 6469 11036
rect 6503 11033 6515 11067
rect 6457 11027 6515 11033
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 8956 11064 8984 11095
rect 9048 11076 9076 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9125 11095 9183 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11790 11132 11796 11144
rect 11751 11104 11796 11132
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11992 11141 12020 11240
rect 12888 11237 12900 11240
rect 12934 11268 12946 11271
rect 13814 11268 13820 11280
rect 12934 11240 13820 11268
rect 12934 11237 12946 11240
rect 12888 11231 12946 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 13924 11268 13952 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 15010 11268 15016 11280
rect 13924 11240 15016 11268
rect 15010 11228 15016 11240
rect 15068 11228 15074 11280
rect 16684 11268 16712 11299
rect 17218 11277 17224 11280
rect 17212 11268 17224 11277
rect 16684 11240 17224 11268
rect 17212 11231 17224 11240
rect 17218 11228 17224 11231
rect 17276 11228 17282 11280
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 13906 11200 13912 11212
rect 12667 11172 13912 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 14921 11203 14979 11209
rect 14921 11200 14933 11203
rect 14148 11172 14933 11200
rect 14148 11160 14154 11172
rect 14921 11169 14933 11172
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15545 11203 15603 11209
rect 15545 11200 15557 11203
rect 15160 11172 15557 11200
rect 15160 11160 15166 11172
rect 15545 11169 15557 11172
rect 15591 11169 15603 11203
rect 15545 11163 15603 11169
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 7515 11036 8984 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 9030 11024 9036 11076
rect 9088 11024 9094 11076
rect 11333 11067 11391 11073
rect 11333 11033 11345 11067
rect 11379 11064 11391 11067
rect 12526 11064 12532 11076
rect 11379 11036 12532 11064
rect 11379 11033 11391 11036
rect 11333 11027 11391 11033
rect 12526 11024 12532 11036
rect 12584 11024 12590 11076
rect 13924 11064 13952 11160
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 16945 11135 17003 11141
rect 16945 11132 16957 11135
rect 15289 11095 15347 11101
rect 16316 11104 16957 11132
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 13924 11036 14749 11064
rect 14737 11033 14749 11036
rect 14783 11064 14795 11067
rect 15304 11064 15332 11095
rect 14783 11036 15332 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 1578 10996 1584 11008
rect 1412 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 3234 10996 3240 11008
rect 3195 10968 3240 10996
rect 3234 10956 3240 10968
rect 3292 10956 3298 11008
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 3476 10968 4077 10996
rect 3476 10956 3482 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 4172 10996 4200 11024
rect 15304 11008 15332 11036
rect 16316 11008 16344 11104
rect 16945 11101 16957 11104
rect 16991 11101 17003 11135
rect 16945 11095 17003 11101
rect 4798 10996 4804 11008
rect 4172 10968 4804 10996
rect 4065 10959 4123 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 8481 10999 8539 11005
rect 8481 10965 8493 10999
rect 8527 10996 8539 10999
rect 9582 10996 9588 11008
rect 8527 10968 9588 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 12618 10996 12624 11008
rect 10652 10968 12624 10996
rect 10652 10956 10658 10968
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13998 10996 14004 11008
rect 13959 10968 14004 10996
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 15286 10996 15292 11008
rect 15199 10968 15292 10996
rect 15286 10956 15292 10968
rect 15344 10996 15350 11008
rect 16298 10996 16304 11008
rect 15344 10968 16304 10996
rect 15344 10956 15350 10968
rect 16298 10956 16304 10968
rect 16356 10956 16362 11008
rect 17586 10956 17592 11008
rect 17644 10996 17650 11008
rect 18325 10999 18383 11005
rect 18325 10996 18337 10999
rect 17644 10968 18337 10996
rect 17644 10956 17650 10968
rect 18325 10965 18337 10968
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1394 10792 1400 10804
rect 1355 10764 1400 10792
rect 1394 10752 1400 10764
rect 1452 10752 1458 10804
rect 3789 10795 3847 10801
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 4246 10792 4252 10804
rect 3835 10764 4252 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 7742 10792 7748 10804
rect 5767 10764 7748 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 10321 10795 10379 10801
rect 8536 10764 10272 10792
rect 8536 10752 8542 10764
rect 8941 10727 8999 10733
rect 8941 10693 8953 10727
rect 8987 10724 8999 10727
rect 9122 10724 9128 10736
rect 8987 10696 9128 10724
rect 8987 10693 8999 10696
rect 8941 10687 8999 10693
rect 9122 10684 9128 10696
rect 9180 10724 9186 10736
rect 10244 10724 10272 10764
rect 10321 10761 10333 10795
rect 10367 10792 10379 10795
rect 10870 10792 10876 10804
rect 10367 10764 10876 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11790 10792 11796 10804
rect 11379 10764 11796 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 13354 10792 13360 10804
rect 12483 10764 13360 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 12802 10724 12808 10736
rect 9180 10696 9812 10724
rect 10244 10696 12808 10724
rect 9180 10684 9186 10696
rect 1946 10656 1952 10668
rect 1907 10628 1952 10656
rect 1946 10616 1952 10628
rect 2004 10656 2010 10668
rect 2130 10656 2136 10668
rect 2004 10628 2136 10656
rect 2004 10616 2010 10628
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 6178 10656 6184 10668
rect 6139 10628 6184 10656
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6362 10656 6368 10668
rect 6323 10628 6368 10656
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9784 10665 9812 10696
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 15381 10727 15439 10733
rect 15381 10693 15393 10727
rect 15427 10724 15439 10727
rect 16114 10724 16120 10736
rect 15427 10696 16120 10724
rect 15427 10693 15439 10696
rect 15381 10687 15439 10693
rect 16114 10684 16120 10696
rect 16172 10684 16178 10736
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9548 10628 9689 10656
rect 9548 10616 9554 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11054 10656 11060 10668
rect 11011 10628 11060 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11480 10628 11805 10656
rect 11480 10616 11486 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12342 10656 12348 10668
rect 12023 10628 12348 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13814 10656 13820 10668
rect 13127 10628 13820 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 14056 10628 14289 10656
rect 14056 10616 14062 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10656 15255 10659
rect 15243 10628 15516 10656
rect 15243 10625 15255 10628
rect 15197 10619 15255 10625
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 2682 10597 2688 10600
rect 2409 10591 2467 10597
rect 2409 10588 2421 10591
rect 1636 10560 2421 10588
rect 1636 10548 1642 10560
rect 2409 10557 2421 10560
rect 2455 10557 2467 10591
rect 2676 10588 2688 10597
rect 2643 10560 2688 10588
rect 2409 10551 2467 10557
rect 2676 10551 2688 10560
rect 2682 10548 2688 10551
rect 2740 10548 2746 10600
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4154 10588 4160 10600
rect 4111 10560 4160 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4332 10591 4390 10597
rect 4332 10557 4344 10591
rect 4378 10588 4390 10591
rect 5902 10588 5908 10600
rect 4378 10560 5908 10588
rect 4378 10557 4390 10560
rect 4332 10551 4390 10557
rect 5902 10548 5908 10560
rect 5960 10548 5966 10600
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7524 10560 7573 10588
rect 7524 10548 7530 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7828 10591 7886 10597
rect 7828 10557 7840 10591
rect 7874 10588 7886 10591
rect 9030 10588 9036 10600
rect 7874 10560 9036 10588
rect 7874 10557 7886 10560
rect 7828 10551 7886 10557
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 9582 10588 9588 10600
rect 9543 10560 9588 10588
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 12584 10560 14105 10588
rect 12584 10548 12590 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 14976 10560 15021 10588
rect 14976 10548 14982 10560
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 3142 10520 3148 10532
rect 1811 10492 3148 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 6089 10523 6147 10529
rect 6089 10489 6101 10523
rect 6135 10520 6147 10523
rect 7650 10520 7656 10532
rect 6135 10492 7656 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 7650 10480 7656 10492
rect 7708 10480 7714 10532
rect 10502 10520 10508 10532
rect 7944 10492 10508 10520
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 3326 10452 3332 10464
rect 1903 10424 3332 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 3326 10412 3332 10424
rect 3384 10452 3390 10464
rect 3694 10452 3700 10464
rect 3384 10424 3700 10452
rect 3384 10412 3390 10424
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 7944 10452 7972 10492
rect 10502 10480 10508 10492
rect 10560 10480 10566 10532
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 10652 10492 10793 10520
rect 10652 10480 10658 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 12802 10520 12808 10532
rect 12763 10492 12808 10520
rect 10781 10483 10839 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 14185 10523 14243 10529
rect 14185 10520 14197 10523
rect 13228 10492 14197 10520
rect 13228 10480 13234 10492
rect 14185 10489 14197 10492
rect 14231 10489 14243 10523
rect 14185 10483 14243 10489
rect 14642 10480 14648 10532
rect 14700 10520 14706 10532
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 14700 10492 15025 10520
rect 14700 10480 14706 10492
rect 15013 10489 15025 10492
rect 15059 10489 15071 10523
rect 15488 10520 15516 10628
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 15746 10656 15752 10668
rect 15620 10628 15752 10656
rect 15620 10616 15626 10628
rect 15746 10616 15752 10628
rect 15804 10656 15810 10668
rect 15838 10656 15844 10668
rect 15804 10628 15844 10656
rect 15804 10616 15810 10628
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 16298 10588 16304 10600
rect 16259 10560 16304 10588
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 16574 10529 16580 10532
rect 16568 10520 16580 10529
rect 15488 10492 16580 10520
rect 15013 10483 15071 10489
rect 16568 10483 16580 10492
rect 16632 10520 16638 10532
rect 17586 10520 17592 10532
rect 16632 10492 17592 10520
rect 16574 10480 16580 10483
rect 16632 10480 16638 10492
rect 17586 10480 17592 10492
rect 17644 10480 17650 10532
rect 4120 10424 7972 10452
rect 4120 10412 4126 10424
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8076 10424 9229 10452
rect 8076 10412 8082 10424
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 9217 10415 9275 10421
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 10686 10452 10692 10464
rect 9456 10424 10692 10452
rect 9456 10412 9462 10424
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11664 10424 11713 10452
rect 11664 10412 11670 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13446 10452 13452 10464
rect 12943 10424 13452 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 13722 10452 13728 10464
rect 13683 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 15749 10455 15807 10461
rect 15749 10452 15761 10455
rect 14599 10424 15761 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 15749 10421 15761 10424
rect 15795 10421 15807 10455
rect 17678 10452 17684 10464
rect 17639 10424 17684 10452
rect 15749 10415 15807 10421
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 18233 10455 18291 10461
rect 18233 10421 18245 10455
rect 18279 10452 18291 10455
rect 18322 10452 18328 10464
rect 18279 10424 18328 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2406 10248 2412 10260
rect 1627 10220 2412 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2590 10248 2596 10260
rect 2551 10220 2596 10248
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 5350 10248 5356 10260
rect 3712 10220 5356 10248
rect 2041 10183 2099 10189
rect 2041 10149 2053 10183
rect 2087 10180 2099 10183
rect 3418 10180 3424 10192
rect 2087 10152 3424 10180
rect 2087 10149 2099 10152
rect 2041 10143 2099 10149
rect 3418 10140 3424 10152
rect 3476 10140 3482 10192
rect 1946 10112 1952 10124
rect 1907 10084 1952 10112
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 2314 10072 2320 10124
rect 2372 10112 2378 10124
rect 2961 10115 3019 10121
rect 2961 10112 2973 10115
rect 2372 10084 2973 10112
rect 2372 10072 2378 10084
rect 2961 10081 2973 10084
rect 3007 10081 3019 10115
rect 2961 10075 3019 10081
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10112 3111 10115
rect 3712 10112 3740 10220
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5534 10248 5540 10260
rect 5447 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10248 5598 10260
rect 5994 10248 6000 10260
rect 5592 10220 6000 10248
rect 5592 10208 5598 10220
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6512 10220 6929 10248
rect 6512 10208 6518 10220
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 6917 10211 6975 10217
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 10870 10248 10876 10260
rect 8444 10220 10876 10248
rect 8444 10208 8450 10220
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11054 10248 11060 10260
rect 11015 10220 11060 10248
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12400 10220 12817 10248
rect 12400 10208 12406 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 13170 10248 13176 10260
rect 13131 10220 13176 10248
rect 12805 10211 12863 10217
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 13538 10208 13544 10260
rect 13596 10248 13602 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 13596 10220 13645 10248
rect 13596 10208 13602 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 14461 10251 14519 10257
rect 14461 10248 14473 10251
rect 13780 10220 14473 10248
rect 13780 10208 13786 10220
rect 14461 10217 14473 10220
rect 14507 10217 14519 10251
rect 14461 10211 14519 10217
rect 15749 10251 15807 10257
rect 15749 10217 15761 10251
rect 15795 10248 15807 10251
rect 16114 10248 16120 10260
rect 15795 10220 16120 10248
rect 15795 10217 15807 10220
rect 15749 10211 15807 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10217 16911 10251
rect 16853 10211 16911 10217
rect 17773 10251 17831 10257
rect 17773 10217 17785 10251
rect 17819 10248 17831 10251
rect 17862 10248 17868 10260
rect 17819 10220 17868 10248
rect 17819 10217 17831 10220
rect 17773 10211 17831 10217
rect 4424 10183 4482 10189
rect 4424 10149 4436 10183
rect 4470 10180 4482 10183
rect 5442 10180 5448 10192
rect 4470 10152 5448 10180
rect 4470 10149 4482 10152
rect 4424 10143 4482 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 7009 10183 7067 10189
rect 7009 10149 7021 10183
rect 7055 10180 7067 10183
rect 7282 10180 7288 10192
rect 7055 10152 7288 10180
rect 7055 10149 7067 10152
rect 7009 10143 7067 10149
rect 7282 10140 7288 10152
rect 7340 10140 7346 10192
rect 7469 10183 7527 10189
rect 7469 10149 7481 10183
rect 7515 10180 7527 10183
rect 9398 10180 9404 10192
rect 7515 10152 9404 10180
rect 7515 10149 7527 10152
rect 7469 10143 7527 10149
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 14090 10180 14096 10192
rect 9508 10152 14096 10180
rect 3099 10084 3740 10112
rect 3789 10115 3847 10121
rect 3099 10081 3111 10084
rect 3053 10075 3111 10081
rect 3789 10081 3801 10115
rect 3835 10112 3847 10115
rect 6730 10112 6736 10124
rect 3835 10084 6736 10112
rect 3835 10081 3847 10084
rect 3789 10075 3847 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 7828 10115 7886 10121
rect 7828 10112 7840 10115
rect 7208 10084 7840 10112
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10013 3203 10047
rect 4154 10044 4160 10056
rect 3145 10007 3203 10013
rect 3620 10016 4160 10044
rect 2148 9976 2176 10004
rect 3160 9976 3188 10007
rect 2148 9948 3188 9976
rect 1578 9868 1584 9920
rect 1636 9908 1642 9920
rect 3620 9917 3648 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5442 10044 5448 10056
rect 5224 10016 5448 10044
rect 5224 10004 5230 10016
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5810 10044 5816 10056
rect 5771 10016 5816 10044
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 7098 10044 7104 10056
rect 5920 10016 7104 10044
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5718 9976 5724 9988
rect 5408 9948 5724 9976
rect 5408 9936 5414 9948
rect 5718 9936 5724 9948
rect 5776 9936 5782 9988
rect 3605 9911 3663 9917
rect 3605 9908 3617 9911
rect 1636 9880 3617 9908
rect 1636 9868 1642 9880
rect 3605 9877 3617 9880
rect 3651 9877 3663 9911
rect 3605 9871 3663 9877
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 5920 9908 5948 10016
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7208 10053 7236 10084
rect 7828 10081 7840 10084
rect 7874 10112 7886 10115
rect 8202 10112 8208 10124
rect 7874 10084 8208 10112
rect 7874 10081 7886 10084
rect 7828 10075 7886 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9508 10121 9536 10152
rect 14090 10140 14096 10152
rect 14148 10140 14154 10192
rect 14366 10180 14372 10192
rect 14327 10152 14372 10180
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 16868 10180 16896 10211
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 15703 10152 16896 10180
rect 16960 10152 17908 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10081 9551 10115
rect 9933 10115 9991 10121
rect 9933 10112 9945 10115
rect 9493 10075 9551 10081
rect 9600 10084 9945 10112
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7524 10016 7573 10044
rect 7524 10004 7530 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 9600 10044 9628 10084
rect 9933 10081 9945 10084
rect 9979 10081 9991 10115
rect 9933 10075 9991 10081
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 11146 10112 11152 10124
rect 10560 10084 11152 10112
rect 10560 10072 10566 10084
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 11692 10115 11750 10121
rect 11692 10081 11704 10115
rect 11738 10112 11750 10115
rect 11974 10112 11980 10124
rect 11738 10084 11980 10112
rect 11738 10081 11750 10084
rect 11692 10075 11750 10081
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 12066 10072 12072 10124
rect 12124 10112 12130 10124
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 12124 10084 13553 10112
rect 12124 10072 12130 10084
rect 13541 10081 13553 10084
rect 13587 10081 13599 10115
rect 13541 10075 13599 10081
rect 14550 10072 14556 10124
rect 14608 10112 14614 10124
rect 14608 10084 16252 10112
rect 14608 10072 14614 10084
rect 7561 10007 7619 10013
rect 8956 10016 9628 10044
rect 6454 9936 6460 9988
rect 6512 9976 6518 9988
rect 7377 9979 7435 9985
rect 7377 9976 7389 9979
rect 6512 9948 7389 9976
rect 6512 9936 6518 9948
rect 7377 9945 7389 9948
rect 7423 9945 7435 9979
rect 7377 9939 7435 9945
rect 3752 9880 5948 9908
rect 6549 9911 6607 9917
rect 3752 9868 3758 9880
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 7558 9908 7564 9920
rect 6595 9880 7564 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 8956 9917 8984 10016
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 9732 10016 9825 10044
rect 10980 10016 11437 10044
rect 9732 10004 9738 10016
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8904 9880 8953 9908
rect 8904 9868 8910 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9692 9908 9720 10004
rect 10980 9920 11008 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 13814 10044 13820 10056
rect 13771 10016 13820 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 15102 10044 15108 10056
rect 14691 10016 15108 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16114 10044 16120 10056
rect 15979 10016 16120 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 16224 10044 16252 10084
rect 16298 10072 16304 10124
rect 16356 10112 16362 10124
rect 16356 10084 16401 10112
rect 16356 10072 16362 10084
rect 16960 10044 16988 10152
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17880 10121 17908 10152
rect 17865 10115 17923 10121
rect 17865 10081 17877 10115
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 17310 10044 17316 10056
rect 16224 10016 16988 10044
rect 17271 10016 17316 10044
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17678 10044 17684 10056
rect 17451 10016 17684 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 13630 9976 13636 9988
rect 13372 9948 13636 9976
rect 10962 9908 10968 9920
rect 9355 9880 10968 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 13372 9908 13400 9948
rect 13630 9936 13636 9948
rect 13688 9976 13694 9988
rect 14918 9976 14924 9988
rect 13688 9948 14924 9976
rect 13688 9936 13694 9948
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 15654 9936 15660 9988
rect 15712 9976 15718 9988
rect 17420 9976 17448 10007
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18046 9976 18052 9988
rect 15712 9948 17448 9976
rect 18007 9948 18052 9976
rect 15712 9936 15718 9948
rect 18046 9936 18052 9948
rect 18104 9936 18110 9988
rect 11112 9880 13400 9908
rect 11112 9868 11118 9880
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 13504 9880 14013 9908
rect 13504 9868 13510 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 14001 9871 14059 9877
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 14516 9880 15301 9908
rect 14516 9868 14522 9880
rect 15289 9877 15301 9880
rect 15335 9877 15347 9911
rect 16482 9908 16488 9920
rect 16443 9880 16488 9908
rect 15289 9871 15347 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 17773 9911 17831 9917
rect 17773 9908 17785 9911
rect 17736 9880 17785 9908
rect 17736 9868 17742 9880
rect 17773 9877 17785 9880
rect 17819 9877 17831 9911
rect 17773 9871 17831 9877
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 5074 9704 5080 9716
rect 3200 9676 5080 9704
rect 3200 9664 3206 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5316 9676 6316 9704
rect 5316 9664 5322 9676
rect 2038 9636 2044 9648
rect 1999 9608 2044 9636
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 4430 9636 4436 9648
rect 3099 9608 4436 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 6288 9636 6316 9676
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6457 9707 6515 9713
rect 6457 9704 6469 9707
rect 6420 9676 6469 9704
rect 6420 9664 6426 9676
rect 6457 9673 6469 9676
rect 6503 9673 6515 9707
rect 14550 9704 14556 9716
rect 6457 9667 6515 9673
rect 6564 9676 14556 9704
rect 6564 9636 6592 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 15286 9704 15292 9716
rect 14936 9676 15292 9704
rect 10226 9636 10232 9648
rect 6288 9608 6592 9636
rect 10187 9608 10232 9636
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 10321 9639 10379 9645
rect 10321 9605 10333 9639
rect 10367 9636 10379 9639
rect 11054 9636 11060 9648
rect 10367 9608 11060 9636
rect 10367 9605 10379 9608
rect 10321 9599 10379 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 12066 9636 12072 9648
rect 11195 9608 12072 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14090 9636 14096 9648
rect 14051 9608 14096 9636
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2590 9568 2596 9580
rect 2188 9540 2596 9568
rect 2188 9528 2194 9540
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 4246 9568 4252 9580
rect 3743 9540 4252 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4396 9540 4537 9568
rect 4396 9528 4402 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4755 9540 5212 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 4154 9500 4160 9512
rect 1535 9472 4160 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5184 9500 5212 9540
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 10873 9571 10931 9577
rect 6788 9540 6960 9568
rect 6788 9528 6794 9540
rect 6641 9503 6699 9509
rect 5184 9472 6408 9500
rect 5077 9463 5135 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 3970 9432 3976 9444
rect 2455 9404 3976 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 3970 9392 3976 9404
rect 4028 9392 4034 9444
rect 4706 9392 4712 9444
rect 4764 9392 4770 9444
rect 5092 9432 5120 9463
rect 6380 9444 6408 9472
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6687 9472 6837 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6932 9500 6960 9540
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 10919 9540 10999 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 9122 9509 9128 9512
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 6932 9472 8677 9500
rect 6825 9463 6883 9469
rect 8665 9469 8677 9472
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8803 9472 8861 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 9116 9500 9128 9509
rect 9083 9472 9128 9500
rect 8849 9463 8907 9469
rect 9116 9463 9128 9472
rect 9122 9460 9128 9463
rect 9180 9460 9186 9512
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 10971 9500 10999 9540
rect 11330 9528 11336 9580
rect 11388 9568 11394 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11388 9540 11621 9568
rect 11388 9528 11394 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 12342 9568 12348 9580
rect 11839 9540 12348 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 12342 9528 12348 9540
rect 12400 9568 12406 9580
rect 14936 9577 14964 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16574 9704 16580 9716
rect 16172 9676 16580 9704
rect 16172 9664 16178 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 16945 9707 17003 9713
rect 16945 9673 16957 9707
rect 16991 9704 17003 9707
rect 17218 9704 17224 9716
rect 16991 9676 17224 9704
rect 16991 9673 17003 9676
rect 16945 9667 17003 9673
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 16206 9636 16212 9648
rect 16080 9608 16212 9636
rect 16080 9596 16086 9608
rect 16206 9596 16212 9608
rect 16264 9636 16270 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 16264 9608 16313 9636
rect 16264 9596 16270 9608
rect 16301 9605 16313 9608
rect 16347 9605 16359 9639
rect 16301 9599 16359 9605
rect 14921 9571 14979 9577
rect 12400 9540 12572 9568
rect 12400 9528 12406 9540
rect 11974 9500 11980 9512
rect 9456 9472 10916 9500
rect 10971 9472 11980 9500
rect 9456 9460 9462 9472
rect 5166 9432 5172 9444
rect 5092 9404 5172 9432
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 5344 9435 5402 9441
rect 5344 9401 5356 9435
rect 5390 9432 5402 9435
rect 5534 9432 5540 9444
rect 5390 9404 5540 9432
rect 5390 9401 5402 9404
rect 5344 9395 5402 9401
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6420 9404 7082 9432
rect 6420 9392 6426 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 7070 9395 7128 9401
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 7374 9432 7380 9444
rect 7248 9404 7380 9432
rect 7248 9392 7254 9404
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 7484 9404 8524 9432
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1673 9367 1731 9373
rect 1673 9364 1685 9367
rect 1452 9336 1685 9364
rect 1452 9324 1458 9336
rect 1673 9333 1685 9336
rect 1719 9333 1731 9367
rect 1673 9327 1731 9333
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 3418 9364 3424 9376
rect 2556 9336 2601 9364
rect 3379 9336 3424 9364
rect 2556 9324 2562 9336
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 4065 9367 4123 9373
rect 3568 9336 3613 9364
rect 3568 9324 3574 9336
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 4338 9364 4344 9376
rect 4111 9336 4344 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4433 9367 4491 9373
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 4724 9364 4752 9392
rect 4982 9364 4988 9376
rect 4479 9336 4988 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5184 9364 5212 9392
rect 7484 9376 7512 9404
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 5184 9336 6653 9364
rect 6641 9333 6653 9336
rect 6687 9364 6699 9367
rect 7466 9364 7472 9376
rect 6687 9336 7472 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 8202 9364 8208 9376
rect 8163 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8496 9373 8524 9404
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 10781 9435 10839 9441
rect 10781 9432 10793 9435
rect 8628 9404 10793 9432
rect 8628 9392 8634 9404
rect 10781 9401 10793 9404
rect 10827 9401 10839 9435
rect 10781 9395 10839 9401
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9364 8539 9367
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8527 9336 8769 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 8757 9327 8815 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10888 9364 10916 9472
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12544 9500 12572 9540
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 16390 9528 16396 9580
rect 16448 9568 16454 9580
rect 17405 9571 17463 9577
rect 17405 9568 17417 9571
rect 16448 9540 17417 9568
rect 16448 9528 16454 9540
rect 17405 9537 17417 9540
rect 17451 9537 17463 9571
rect 17586 9568 17592 9580
rect 17547 9540 17592 9568
rect 17405 9531 17463 9537
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 18966 9568 18972 9580
rect 18927 9540 18972 9568
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 12693 9503 12751 9509
rect 12693 9500 12705 9503
rect 12544 9472 12705 9500
rect 12437 9463 12495 9469
rect 12693 9469 12705 9472
rect 12739 9469 12751 9503
rect 12693 9463 12751 9469
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 12452 9432 12480 9463
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 13964 9472 14289 9500
rect 13964 9460 13970 9472
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 15188 9503 15246 9509
rect 15188 9469 15200 9503
rect 15234 9500 15246 9503
rect 15654 9500 15660 9512
rect 15234 9472 15660 9500
rect 15234 9469 15246 9472
rect 15188 9463 15246 9469
rect 11020 9404 12480 9432
rect 11020 9392 11026 9404
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 14384 9432 14412 9463
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9500 17371 9503
rect 17770 9500 17776 9512
rect 17359 9472 17776 9500
rect 17359 9469 17371 9472
rect 17313 9463 17371 9469
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 14826 9432 14832 9444
rect 13320 9404 14412 9432
rect 14476 9404 14832 9432
rect 13320 9392 13326 9404
rect 11146 9364 11152 9376
rect 10888 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9364 11210 9376
rect 11422 9364 11428 9376
rect 11204 9336 11428 9364
rect 11204 9324 11210 9336
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 11606 9364 11612 9376
rect 11563 9336 11612 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11606 9324 11612 9336
rect 11664 9364 11670 9376
rect 14476 9364 14504 9404
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 18064 9432 18092 9463
rect 15068 9404 18092 9432
rect 15068 9392 15074 9404
rect 17788 9376 17816 9404
rect 11664 9336 14504 9364
rect 14553 9367 14611 9373
rect 11664 9324 11670 9336
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 15286 9364 15292 9376
rect 14599 9336 15292 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 17770 9324 17776 9376
rect 17828 9324 17834 9376
rect 18230 9364 18236 9376
rect 18191 9336 18236 9364
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2648 9132 2789 9160
rect 2648 9120 2654 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 2777 9123 2835 9129
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 4801 9163 4859 9169
rect 4801 9160 4813 9163
rect 3568 9132 4813 9160
rect 3568 9120 3574 9132
rect 4801 9129 4813 9132
rect 4847 9129 4859 9163
rect 4801 9123 4859 9129
rect 5169 9163 5227 9169
rect 5169 9129 5181 9163
rect 5215 9160 5227 9163
rect 5258 9160 5264 9172
rect 5215 9132 5264 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 5868 9132 6193 9160
rect 5868 9120 5874 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 6181 9123 6239 9129
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6328 9132 6373 9160
rect 6328 9120 6334 9132
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6788 9132 6837 9160
rect 6788 9120 6794 9132
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 7558 9160 7564 9172
rect 7519 9132 7564 9160
rect 6825 9123 6883 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7708 9132 8125 9160
rect 7708 9120 7714 9132
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 8113 9123 8171 9129
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 9214 9160 9220 9172
rect 8619 9132 9220 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 10686 9160 10692 9172
rect 10367 9132 10692 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 14366 9160 14372 9172
rect 12400 9132 14372 9160
rect 12400 9120 12406 9132
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 14550 9160 14556 9172
rect 14511 9132 14556 9160
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14645 9163 14703 9169
rect 14645 9129 14657 9163
rect 14691 9160 14703 9163
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 14691 9132 15025 9160
rect 14691 9129 14703 9132
rect 14645 9123 14703 9129
rect 15013 9129 15025 9132
rect 15059 9160 15071 9163
rect 15194 9160 15200 9172
rect 15059 9132 15200 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17405 9163 17463 9169
rect 17405 9160 17417 9163
rect 17368 9132 17417 9160
rect 17368 9120 17374 9132
rect 17405 9129 17417 9132
rect 17451 9129 17463 9163
rect 17770 9160 17776 9172
rect 17731 9132 17776 9160
rect 17405 9123 17463 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 4706 9092 4712 9104
rect 3068 9064 4712 9092
rect 1664 9027 1722 9033
rect 1664 8993 1676 9027
rect 1710 9024 1722 9027
rect 2682 9024 2688 9036
rect 1710 8996 2688 9024
rect 1710 8993 1722 8996
rect 1664 8987 1722 8993
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3068 9033 3096 9064
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 6362 9052 6368 9104
rect 6420 9092 6426 9104
rect 7834 9092 7840 9104
rect 6420 9064 7840 9092
rect 6420 9052 6426 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 8941 9095 8999 9101
rect 8941 9092 8953 9095
rect 8812 9064 8953 9092
rect 8812 9052 8818 9064
rect 8941 9061 8953 9064
rect 8987 9092 8999 9095
rect 9030 9092 9036 9104
rect 8987 9064 9036 9092
rect 8987 9061 8999 9064
rect 8941 9055 8999 9061
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9674 9092 9680 9104
rect 9131 9064 9680 9092
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 8993 3111 9027
rect 3053 8987 3111 8993
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 7466 9024 7472 9036
rect 7427 8996 7472 9024
rect 7009 8987 7067 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1412 8820 1440 8919
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 3068 8956 3096 8987
rect 2464 8928 3096 8956
rect 4080 8956 4108 8987
rect 5258 8956 5264 8968
rect 4080 8928 5264 8956
rect 2464 8916 2470 8928
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 5408 8928 6377 8956
rect 5408 8916 5414 8928
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 7024 8956 7052 8987
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 8846 9024 8852 9036
rect 7760 8996 8852 9024
rect 7374 8956 7380 8968
rect 7024 8928 7380 8956
rect 6365 8919 6423 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7760 8965 7788 8996
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 9131 9024 9159 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 13538 9092 13544 9104
rect 13451 9064 13544 9092
rect 13538 9052 13544 9064
rect 13596 9092 13602 9104
rect 17678 9092 17684 9104
rect 13596 9064 17684 9092
rect 13596 9052 13602 9064
rect 17678 9052 17684 9064
rect 17736 9092 17742 9104
rect 17865 9095 17923 9101
rect 17865 9092 17877 9095
rect 17736 9064 17877 9092
rect 17736 9052 17742 9064
rect 17865 9061 17877 9064
rect 17911 9061 17923 9095
rect 17865 9055 17923 9061
rect 10226 9024 10232 9036
rect 8947 8996 9159 9024
rect 9232 8996 10232 9024
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 3418 8848 3424 8900
rect 3476 8888 3482 8900
rect 5813 8891 5871 8897
rect 5813 8888 5825 8891
rect 3476 8860 5825 8888
rect 3476 8848 3482 8860
rect 5813 8857 5825 8860
rect 5859 8857 5871 8891
rect 8947 8888 8975 8996
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8956 9091 8959
rect 9122 8956 9128 8968
rect 9079 8928 9128 8956
rect 9079 8925 9091 8928
rect 9033 8919 9091 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9232 8965 9260 8996
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10686 9024 10692 9036
rect 10647 8996 10692 9024
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 9024 10839 9027
rect 11422 9024 11428 9036
rect 10827 8996 11428 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11606 9033 11612 9036
rect 11600 8987 11612 9033
rect 11664 9024 11670 9036
rect 14001 9027 14059 9033
rect 11664 8996 11700 9024
rect 11606 8984 11612 8987
rect 11664 8984 11670 8996
rect 14001 8993 14013 9027
rect 14047 9024 14059 9027
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 14047 8996 15025 9024
rect 14047 8993 14059 8996
rect 14001 8987 14059 8993
rect 15013 8993 15025 8996
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 15378 8984 15384 9036
rect 15436 9024 15442 9036
rect 16022 9033 16028 9036
rect 15749 9027 15807 9033
rect 15749 9024 15761 9027
rect 15436 8996 15761 9024
rect 15436 8984 15442 8996
rect 15749 8993 15761 8996
rect 15795 8993 15807 9027
rect 16016 9024 16028 9033
rect 15983 8996 16028 9024
rect 15749 8987 15807 8993
rect 16016 8987 16028 8996
rect 16022 8984 16028 8987
rect 16080 8984 16086 9036
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 10410 8956 10416 8968
rect 9217 8919 9275 8925
rect 9324 8928 10416 8956
rect 5813 8851 5871 8857
rect 5920 8860 8975 8888
rect 9140 8888 9168 8916
rect 9324 8888 9352 8928
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10870 8956 10876 8968
rect 10831 8928 10876 8956
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11020 8928 11345 8956
rect 11020 8916 11026 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 13630 8956 13636 8968
rect 13591 8928 13636 8956
rect 11333 8919 11391 8925
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13814 8956 13820 8968
rect 13775 8928 13820 8956
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 14826 8956 14832 8968
rect 14787 8928 14832 8956
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14976 8928 15301 8956
rect 14976 8916 14982 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17644 8928 17969 8956
rect 17644 8916 17650 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 9140 8860 9352 8888
rect 13173 8891 13231 8897
rect 1578 8820 1584 8832
rect 1412 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3200 8792 3249 8820
rect 3200 8780 3206 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4798 8820 4804 8832
rect 4295 8792 4804 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5920 8820 5948 8860
rect 13173 8857 13185 8891
rect 13219 8888 13231 8891
rect 13219 8860 15792 8888
rect 13219 8857 13231 8860
rect 13173 8851 13231 8857
rect 5040 8792 5948 8820
rect 5040 8780 5046 8792
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6546 8820 6552 8832
rect 6420 8792 6552 8820
rect 6420 8780 6426 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 7101 8823 7159 8829
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 7282 8820 7288 8832
rect 7147 8792 7288 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 9306 8820 9312 8832
rect 8444 8792 9312 8820
rect 8444 8780 8450 8792
rect 9306 8780 9312 8792
rect 9364 8820 9370 8832
rect 10318 8820 10324 8832
rect 9364 8792 10324 8820
rect 9364 8780 9370 8792
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 12713 8823 12771 8829
rect 12713 8820 12725 8823
rect 10928 8792 12725 8820
rect 10928 8780 10934 8792
rect 12713 8789 12725 8792
rect 12759 8789 12771 8823
rect 12713 8783 12771 8789
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 14001 8823 14059 8829
rect 14001 8820 14013 8823
rect 13596 8792 14013 8820
rect 13596 8780 13602 8792
rect 14001 8789 14013 8792
rect 14047 8789 14059 8823
rect 14182 8820 14188 8832
rect 14143 8792 14188 8820
rect 14001 8783 14059 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 15378 8820 15384 8832
rect 14332 8792 15384 8820
rect 14332 8780 14338 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15764 8820 15792 8860
rect 16942 8820 16948 8832
rect 15764 8792 16948 8820
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17126 8820 17132 8832
rect 17087 8792 17132 8820
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 2498 8616 2504 8628
rect 1535 8588 2504 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3844 8588 3893 8616
rect 3844 8576 3850 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 6917 8619 6975 8625
rect 4396 8588 5764 8616
rect 4396 8576 4402 8588
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2179 8452 2636 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2608 8424 2636 8452
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 5736 8480 5764 8588
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 7466 8616 7472 8628
rect 6963 8588 7472 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 7926 8616 7932 8628
rect 7887 8588 7932 8616
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 10962 8616 10968 8628
rect 8895 8588 10968 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 5902 8508 5908 8560
rect 5960 8548 5966 8560
rect 5997 8551 6055 8557
rect 5997 8548 6009 8551
rect 5960 8520 6009 8548
rect 5960 8508 5966 8520
rect 5997 8517 6009 8520
rect 6043 8517 6055 8551
rect 5997 8511 6055 8517
rect 6362 8508 6368 8560
rect 6420 8548 6426 8560
rect 8938 8548 8944 8560
rect 6420 8520 8944 8548
rect 6420 8508 6426 8520
rect 8938 8508 8944 8520
rect 8996 8508 9002 8560
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 3752 8452 4292 8480
rect 5736 8452 7389 8480
rect 3752 8440 3758 8452
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 1636 8384 2513 8412
rect 1636 8372 1642 8384
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 1949 8347 2007 8353
rect 1949 8344 1961 8347
rect 1728 8316 1961 8344
rect 1728 8304 1734 8316
rect 1949 8313 1961 8316
rect 1995 8313 2007 8347
rect 2516 8344 2544 8375
rect 2590 8372 2596 8424
rect 2648 8372 2654 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 2700 8384 4169 8412
rect 2700 8344 2728 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4264 8412 4292 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 8202 8480 8208 8492
rect 7607 8452 8208 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8478 8480 8484 8492
rect 8435 8452 8484 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8619 8452 9076 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 5718 8412 5724 8424
rect 4264 8384 5724 8412
rect 4157 8375 4215 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8381 5871 8415
rect 5813 8375 5871 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7742 8412 7748 8424
rect 7331 8384 7748 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 2516 8316 2728 8344
rect 2768 8347 2826 8353
rect 1949 8307 2007 8313
rect 2768 8313 2780 8347
rect 2814 8344 2826 8347
rect 4246 8344 4252 8356
rect 2814 8316 4252 8344
rect 2814 8313 2826 8316
rect 2768 8307 2826 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 4430 8353 4436 8356
rect 4424 8344 4436 8353
rect 4391 8316 4436 8344
rect 4424 8307 4436 8316
rect 4488 8344 4494 8356
rect 5350 8344 5356 8356
rect 4488 8316 5356 8344
rect 4430 8304 4436 8307
rect 4488 8304 4494 8316
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5828 8344 5856 8375
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 7984 8384 8309 8412
rect 7984 8372 7990 8384
rect 8297 8381 8309 8384
rect 8343 8412 8355 8415
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8343 8384 8769 8412
rect 8343 8381 8355 8384
rect 8297 8375 8355 8381
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8895 8384 8953 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 9048 8412 9076 8452
rect 9208 8415 9266 8421
rect 9208 8412 9220 8415
rect 9048 8384 9220 8412
rect 8941 8375 8999 8381
rect 9208 8381 9220 8384
rect 9254 8412 9266 8415
rect 10042 8412 10048 8424
rect 9254 8384 10048 8412
rect 9254 8381 9266 8384
rect 9208 8375 9266 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10152 8412 10180 8588
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11974 8616 11980 8628
rect 11935 8588 11980 8616
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 15562 8616 15568 8628
rect 13219 8588 15568 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18279 8588 18981 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18969 8585 18981 8588
rect 19015 8585 19027 8619
rect 18969 8579 19027 8585
rect 10318 8548 10324 8560
rect 10279 8520 10324 8548
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8548 12863 8551
rect 13814 8548 13820 8560
rect 12851 8520 13820 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 13538 8480 13544 8492
rect 10284 8452 10732 8480
rect 10284 8440 10290 8452
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 10152 8384 10609 8412
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10704 8412 10732 8452
rect 11624 8452 13544 8480
rect 11624 8412 11652 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13722 8480 13728 8492
rect 13683 8452 13728 8480
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 15378 8440 15384 8492
rect 15436 8480 15442 8492
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 15436 8452 16313 8480
rect 15436 8440 15442 8452
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 10704 8384 11652 8412
rect 10597 8375 10655 8381
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 11756 8384 12633 8412
rect 11756 8372 11762 8384
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 12621 8375 12679 8381
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8412 13691 8415
rect 13998 8412 14004 8424
rect 13679 8384 14004 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14185 8415 14243 8421
rect 14185 8381 14197 8415
rect 14231 8412 14243 8415
rect 14274 8412 14280 8424
rect 14231 8384 14280 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 16206 8412 16212 8424
rect 14384 8384 16212 8412
rect 5828 8316 9536 8344
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 4062 8276 4068 8288
rect 1903 8248 4068 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4264 8276 4292 8304
rect 5534 8276 5540 8288
rect 4264 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 8478 8276 8484 8288
rect 6144 8248 8484 8276
rect 6144 8236 6150 8248
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8757 8279 8815 8285
rect 8757 8245 8769 8279
rect 8803 8276 8815 8279
rect 9398 8276 9404 8288
rect 8803 8248 9404 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9508 8276 9536 8316
rect 9582 8304 9588 8356
rect 9640 8344 9646 8356
rect 10870 8353 10876 8356
rect 10864 8344 10876 8353
rect 9640 8316 10876 8344
rect 9640 8304 9646 8316
rect 10864 8307 10876 8316
rect 10870 8304 10876 8307
rect 10928 8304 10934 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 12158 8344 12164 8356
rect 11112 8316 12164 8344
rect 11112 8304 11118 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 13541 8347 13599 8353
rect 13541 8313 13553 8347
rect 13587 8344 13599 8347
rect 14384 8344 14412 8384
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16557 8415 16615 8421
rect 16557 8412 16569 8415
rect 16448 8384 16569 8412
rect 16448 8372 16454 8384
rect 16557 8381 16569 8384
rect 16603 8412 16615 8415
rect 16603 8384 17264 8412
rect 16603 8381 16615 8384
rect 16557 8375 16615 8381
rect 17236 8356 17264 8384
rect 17494 8372 17500 8424
rect 17552 8412 17558 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17552 8384 18061 8412
rect 17552 8372 17558 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 13587 8316 14412 8344
rect 14452 8347 14510 8353
rect 13587 8313 13599 8316
rect 13541 8307 13599 8313
rect 14452 8313 14464 8347
rect 14498 8344 14510 8347
rect 14826 8344 14832 8356
rect 14498 8316 14832 8344
rect 14498 8313 14510 8316
rect 14452 8307 14510 8313
rect 10226 8276 10232 8288
rect 9508 8248 10232 8276
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 13722 8236 13728 8288
rect 13780 8276 13786 8288
rect 14476 8276 14504 8307
rect 14826 8304 14832 8316
rect 14884 8344 14890 8356
rect 14884 8316 16528 8344
rect 14884 8304 14890 8316
rect 13780 8248 14504 8276
rect 13780 8236 13786 8248
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 15565 8279 15623 8285
rect 15565 8276 15577 8279
rect 15252 8248 15577 8276
rect 15252 8236 15258 8248
rect 15565 8245 15577 8248
rect 15611 8245 15623 8279
rect 15565 8239 15623 8245
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15712 8248 15853 8276
rect 15712 8236 15718 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 16500 8276 16528 8316
rect 17218 8304 17224 8356
rect 17276 8304 17282 8356
rect 17678 8276 17684 8288
rect 16500 8248 17684 8276
rect 15841 8239 15899 8245
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2740 8044 2973 8072
rect 2740 8032 2746 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4893 8075 4951 8081
rect 4893 8072 4905 8075
rect 4580 8044 4905 8072
rect 4580 8032 4586 8044
rect 4893 8041 4905 8044
rect 4939 8041 4951 8075
rect 4893 8035 4951 8041
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 5776 8044 6377 8072
rect 5776 8032 5782 8044
rect 6365 8041 6377 8044
rect 6411 8072 6423 8075
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 6411 8044 7849 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 8570 8072 8576 8084
rect 8531 8044 8576 8072
rect 7837 8035 7895 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 10410 8072 10416 8084
rect 8996 8044 10416 8072
rect 8996 8032 9002 8044
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 11480 8044 12173 8072
rect 11480 8032 11486 8044
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12492 8044 12633 8072
rect 12492 8032 12498 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8041 13231 8075
rect 13173 8035 13231 8041
rect 1848 8007 1906 8013
rect 1848 7973 1860 8007
rect 1894 8004 1906 8007
rect 3786 8004 3792 8016
rect 1894 7976 3792 8004
rect 1894 7973 1906 7976
rect 1848 7967 1906 7973
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 5994 7964 6000 8016
rect 6052 8004 6058 8016
rect 6638 8004 6644 8016
rect 6052 7976 6644 8004
rect 6052 7964 6058 7976
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 9033 8007 9091 8013
rect 9033 7973 9045 8007
rect 9079 8004 9091 8007
rect 11238 8004 11244 8016
rect 9079 7976 11244 8004
rect 9079 7973 9091 7976
rect 9033 7967 9091 7973
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 13188 8004 13216 8035
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13412 8044 13645 8072
rect 13412 8032 13418 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14240 8044 14657 8072
rect 14240 8032 14246 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 15703 8044 17509 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 14553 8007 14611 8013
rect 14553 8004 14565 8007
rect 13188 7976 14565 8004
rect 14553 7973 14565 7976
rect 14599 7973 14611 8007
rect 14553 7967 14611 7973
rect 15562 7964 15568 8016
rect 15620 8004 15626 8016
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 15620 7976 15761 8004
rect 15620 7964 15626 7976
rect 15749 7973 15761 7976
rect 15795 7973 15807 8007
rect 16853 8007 16911 8013
rect 16853 8004 16865 8007
rect 15749 7967 15807 7973
rect 16776 7976 16865 8004
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7905 3295 7939
rect 4062 7936 4068 7948
rect 4023 7908 4068 7936
rect 3237 7899 3295 7905
rect 3252 7868 3280 7899
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 4304 7908 5273 7936
rect 4304 7896 4310 7908
rect 5261 7905 5273 7908
rect 5307 7905 5319 7939
rect 5261 7899 5319 7905
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 6546 7936 6552 7948
rect 6319 7908 6552 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7742 7936 7748 7948
rect 7331 7908 7748 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7926 7936 7932 7948
rect 7887 7908 7932 7936
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9861 7939 9919 7945
rect 8987 7908 9812 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 4522 7868 4528 7880
rect 3252 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 4764 7840 5365 7868
rect 4764 7828 4770 7840
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5534 7868 5540 7880
rect 5495 7840 5540 7868
rect 5353 7831 5411 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6503 7840 6592 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 4982 7800 4988 7812
rect 4295 7772 4988 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4982 7760 4988 7772
rect 5040 7760 5046 7812
rect 6564 7800 6592 7840
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7248 7840 7389 7868
rect 7248 7828 7254 7840
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9582 7868 9588 7880
rect 9263 7840 9588 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 6822 7800 6828 7812
rect 6564 7772 6828 7800
rect 6822 7760 6828 7772
rect 6880 7800 6886 7812
rect 7576 7800 7604 7831
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9784 7868 9812 7908
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 10778 7936 10784 7948
rect 9907 7908 10784 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11164 7908 12081 7936
rect 10962 7868 10968 7880
rect 9784 7840 10968 7868
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 6880 7772 7604 7800
rect 7837 7803 7895 7809
rect 6880 7760 6886 7772
rect 7837 7769 7849 7803
rect 7883 7800 7895 7803
rect 10594 7800 10600 7812
rect 7883 7772 10600 7800
rect 7883 7769 7895 7772
rect 7837 7763 7895 7769
rect 10594 7760 10600 7772
rect 10652 7800 10658 7812
rect 11054 7800 11060 7812
rect 10652 7772 11060 7800
rect 10652 7760 10658 7772
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 3418 7732 3424 7744
rect 3379 7704 3424 7732
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 5905 7735 5963 7741
rect 5905 7732 5917 7735
rect 4396 7704 5917 7732
rect 4396 7692 4402 7704
rect 5905 7701 5917 7704
rect 5951 7701 5963 7735
rect 5905 7695 5963 7701
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6052 7704 6929 7732
rect 6052 7692 6058 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 6917 7695 6975 7701
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 8113 7735 8171 7741
rect 8113 7732 8125 7735
rect 7524 7704 8125 7732
rect 7524 7692 7530 7704
rect 8113 7701 8125 7704
rect 8159 7701 8171 7735
rect 8113 7695 8171 7701
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 9030 7732 9036 7744
rect 8536 7704 9036 7732
rect 8536 7692 8542 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 11164 7741 11192 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 13170 7936 13176 7948
rect 12575 7908 13176 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 16666 7936 16672 7948
rect 13587 7908 16672 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12308 7840 12725 7868
rect 12308 7828 12314 7840
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14829 7871 14887 7877
rect 13780 7840 13825 7868
rect 13780 7828 13786 7840
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 15194 7868 15200 7880
rect 14875 7840 15200 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 15194 7828 15200 7840
rect 15252 7868 15258 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15252 7840 15853 7868
rect 15252 7828 15258 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16356 7840 16620 7868
rect 16356 7828 16362 7840
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 15010 7800 15016 7812
rect 13872 7772 15016 7800
rect 13872 7760 13878 7772
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 15562 7800 15568 7812
rect 15396 7772 15568 7800
rect 11149 7735 11207 7741
rect 11149 7732 11161 7735
rect 9640 7704 11161 7732
rect 9640 7692 9646 7704
rect 11149 7701 11161 7704
rect 11195 7701 11207 7735
rect 11149 7695 11207 7701
rect 11885 7735 11943 7741
rect 11885 7701 11897 7735
rect 11931 7732 11943 7735
rect 13906 7732 13912 7744
rect 11931 7704 13912 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 15102 7732 15108 7744
rect 14231 7704 15108 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15396 7732 15424 7772
rect 15562 7760 15568 7772
rect 15620 7760 15626 7812
rect 16206 7760 16212 7812
rect 16264 7800 16270 7812
rect 16485 7803 16543 7809
rect 16485 7800 16497 7803
rect 16264 7772 16497 7800
rect 16264 7760 16270 7772
rect 16485 7769 16497 7772
rect 16531 7769 16543 7803
rect 16485 7763 16543 7769
rect 15335 7704 15424 7732
rect 16592 7732 16620 7840
rect 16776 7800 16804 7976
rect 16853 7973 16865 7976
rect 16899 7973 16911 8007
rect 16853 7967 16911 7973
rect 16942 7964 16948 8016
rect 17000 8004 17006 8016
rect 17957 8007 18015 8013
rect 17957 8004 17969 8007
rect 17000 7976 17969 8004
rect 17000 7964 17006 7976
rect 17957 7973 17969 7976
rect 18003 7973 18015 8007
rect 17957 7967 18015 7973
rect 17310 7936 17316 7948
rect 16960 7908 17316 7936
rect 16960 7880 16988 7908
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 17865 7939 17923 7945
rect 17865 7936 17877 7939
rect 17512 7908 17877 7936
rect 16942 7868 16948 7880
rect 16903 7840 16948 7868
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 17218 7868 17224 7880
rect 17175 7840 17224 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 16850 7800 16856 7812
rect 16776 7772 16856 7800
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 17512 7732 17540 7908
rect 17865 7905 17877 7908
rect 17911 7905 17923 7939
rect 17865 7899 17923 7905
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17736 7840 18061 7868
rect 17736 7828 17742 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 16592 7704 17540 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 1946 7528 1952 7540
rect 1719 7500 1952 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 2682 7528 2688 7540
rect 2643 7500 2688 7528
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 4246 7528 4252 7540
rect 3743 7500 4252 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4706 7528 4712 7540
rect 4667 7500 4712 7528
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5583 7500 5733 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 5721 7491 5779 7497
rect 6104 7500 8217 7528
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 3605 7463 3663 7469
rect 3605 7460 3617 7463
rect 2924 7432 3617 7460
rect 2924 7420 2930 7432
rect 3605 7429 3617 7432
rect 3651 7429 3663 7463
rect 4338 7460 4344 7472
rect 3605 7423 3663 7429
rect 4172 7432 4344 7460
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2590 7392 2596 7404
rect 2363 7364 2596 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 4172 7401 4200 7432
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 5994 7460 6000 7472
rect 5184 7432 6000 7460
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4430 7392 4436 7404
rect 4295 7364 4436 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 2222 7324 2228 7336
rect 1912 7296 2228 7324
rect 1912 7284 1918 7296
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 3344 7324 3372 7355
rect 4430 7352 4436 7364
rect 4488 7392 4494 7404
rect 5184 7401 5212 7432
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 5169 7395 5227 7401
rect 4488 7364 5120 7392
rect 4488 7352 4494 7364
rect 4890 7324 4896 7336
rect 3344 7296 4896 7324
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5092 7324 5120 7364
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 6104 7392 6132 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 10505 7531 10563 7537
rect 10505 7497 10517 7531
rect 10551 7528 10563 7531
rect 10686 7528 10692 7540
rect 10551 7500 10692 7528
rect 10551 7497 10563 7500
rect 10505 7491 10563 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10778 7488 10784 7540
rect 10836 7528 10842 7540
rect 11974 7528 11980 7540
rect 10836 7500 11980 7528
rect 10836 7488 10842 7500
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12492 7500 12537 7528
rect 12492 7488 12498 7500
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 16485 7531 16543 7537
rect 16485 7528 16497 7531
rect 14056 7500 16497 7528
rect 14056 7488 14062 7500
rect 16485 7497 16497 7500
rect 16531 7497 16543 7531
rect 16485 7491 16543 7497
rect 6822 7420 6828 7472
rect 6880 7420 6886 7472
rect 12250 7460 12256 7472
rect 11624 7432 12256 7460
rect 5399 7364 6132 7392
rect 6365 7395 6423 7401
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6546 7392 6552 7404
rect 6411 7364 6552 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 5368 7324 5396 7355
rect 6546 7352 6552 7364
rect 6604 7392 6610 7404
rect 6840 7392 6868 7420
rect 11624 7404 11652 7432
rect 12250 7420 12256 7432
rect 12308 7460 12314 7472
rect 12308 7432 13032 7460
rect 12308 7420 12314 7432
rect 6604 7364 6960 7392
rect 6604 7352 6610 7364
rect 5092 7296 5396 7324
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6932 7324 6960 7364
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 10284 7364 10977 7392
rect 10284 7352 10290 7364
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11606 7392 11612 7404
rect 11195 7364 11612 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 13004 7401 13032 7432
rect 15010 7420 15016 7472
rect 15068 7460 15074 7472
rect 15068 7432 15884 7460
rect 15068 7420 15074 7432
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11756 7364 11897 7392
rect 11756 7352 11762 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 15102 7352 15108 7404
rect 15160 7392 15166 7404
rect 15160 7364 15424 7392
rect 15160 7352 15166 7364
rect 7081 7327 7139 7333
rect 7081 7324 7093 7327
rect 6932 7296 7093 7324
rect 6825 7287 6883 7293
rect 7081 7293 7093 7296
rect 7127 7293 7139 7327
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 7081 7287 7139 7293
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 10778 7324 10784 7336
rect 8628 7296 10784 7324
rect 8628 7284 8634 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10919 7296 13492 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 2314 7256 2320 7268
rect 2087 7228 2320 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 2314 7216 2320 7228
rect 2372 7216 2378 7268
rect 3053 7259 3111 7265
rect 3053 7225 3065 7259
rect 3099 7256 3111 7259
rect 5077 7259 5135 7265
rect 3099 7228 5028 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2406 7188 2412 7200
rect 2280 7160 2412 7188
rect 2280 7148 2286 7160
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 3145 7191 3203 7197
rect 3145 7157 3157 7191
rect 3191 7188 3203 7191
rect 3326 7188 3332 7200
rect 3191 7160 3332 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3651 7160 4077 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 4065 7157 4077 7160
rect 4111 7188 4123 7191
rect 4430 7188 4436 7200
rect 4111 7160 4436 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 5000 7188 5028 7228
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5123 7228 5549 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5537 7225 5549 7228
rect 5583 7225 5595 7259
rect 8110 7256 8116 7268
rect 5537 7219 5595 7225
rect 5828 7228 8116 7256
rect 5828 7188 5856 7228
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 8386 7216 8392 7268
rect 8444 7256 8450 7268
rect 8726 7259 8784 7265
rect 8726 7256 8738 7259
rect 8444 7228 8738 7256
rect 8444 7216 8450 7228
rect 8726 7225 8738 7228
rect 8772 7225 8784 7259
rect 8726 7219 8784 7225
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 11664 7228 11713 7256
rect 11664 7216 11670 7228
rect 11701 7225 11713 7228
rect 11747 7256 11759 7259
rect 12066 7256 12072 7268
rect 11747 7228 12072 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 12710 7216 12716 7268
rect 12768 7256 12774 7268
rect 12897 7259 12955 7265
rect 12897 7256 12909 7259
rect 12768 7228 12909 7256
rect 12768 7216 12774 7228
rect 12897 7225 12909 7228
rect 12943 7225 12955 7259
rect 12897 7219 12955 7225
rect 5000 7160 5856 7188
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6089 7191 6147 7197
rect 6089 7188 6101 7191
rect 6052 7160 6101 7188
rect 6052 7148 6058 7160
rect 6089 7157 6101 7160
rect 6135 7157 6147 7191
rect 6089 7151 6147 7157
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6638 7188 6644 7200
rect 6227 7160 6644 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 9490 7188 9496 7200
rect 8352 7160 9496 7188
rect 8352 7148 8358 7160
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 9861 7191 9919 7197
rect 9861 7188 9873 7191
rect 9824 7160 9873 7188
rect 9824 7148 9830 7160
rect 9861 7157 9873 7160
rect 9907 7157 9919 7191
rect 9861 7151 9919 7157
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11112 7160 11345 7188
rect 11112 7148 11118 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11790 7188 11796 7200
rect 11751 7160 11796 7188
rect 11333 7151 11391 7157
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 12526 7188 12532 7200
rect 11940 7160 12532 7188
rect 11940 7148 11946 7160
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12676 7160 12817 7188
rect 12676 7148 12682 7160
rect 12805 7157 12817 7160
rect 12851 7188 12863 7191
rect 13354 7188 13360 7200
rect 12851 7160 13360 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13464 7188 13492 7296
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 13640 7327 13698 7333
rect 13640 7324 13652 7327
rect 13596 7296 13652 7324
rect 13596 7284 13602 7296
rect 13640 7293 13652 7296
rect 13686 7293 13698 7327
rect 15396 7324 15424 7364
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15856 7401 15884 7432
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 15620 7364 15761 7392
rect 15620 7352 15626 7364
rect 15749 7361 15761 7364
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17218 7392 17224 7404
rect 17175 7364 17224 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 15657 7327 15715 7333
rect 15657 7324 15669 7327
rect 15396 7296 15669 7324
rect 13640 7287 13698 7293
rect 15657 7293 15669 7296
rect 15703 7293 15715 7327
rect 15657 7287 15715 7293
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 17497 7327 17555 7333
rect 17497 7324 17509 7327
rect 16724 7296 17509 7324
rect 16724 7284 16730 7296
rect 17497 7293 17509 7296
rect 17543 7293 17555 7327
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 17497 7287 17555 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 13900 7259 13958 7265
rect 13900 7225 13912 7259
rect 13946 7256 13958 7259
rect 15194 7256 15200 7268
rect 13946 7228 15200 7256
rect 13946 7225 13958 7228
rect 13900 7219 13958 7225
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 16632 7228 16988 7256
rect 16632 7216 16638 7228
rect 14918 7188 14924 7200
rect 13464 7160 14924 7188
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15286 7188 15292 7200
rect 15068 7160 15113 7188
rect 15247 7160 15292 7188
rect 15068 7148 15074 7160
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 16482 7188 16488 7200
rect 15620 7160 16488 7188
rect 15620 7148 15626 7160
rect 16482 7148 16488 7160
rect 16540 7188 16546 7200
rect 16960 7197 16988 7228
rect 16853 7191 16911 7197
rect 16853 7188 16865 7191
rect 16540 7160 16865 7188
rect 16540 7148 16546 7160
rect 16853 7157 16865 7160
rect 16899 7157 16911 7191
rect 16853 7151 16911 7157
rect 16945 7191 17003 7197
rect 16945 7157 16957 7191
rect 16991 7188 17003 7191
rect 17586 7188 17592 7200
rect 16991 7160 17592 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18233 7191 18291 7197
rect 18233 7188 18245 7191
rect 17920 7160 18245 7188
rect 17920 7148 17926 7160
rect 18233 7157 18245 7160
rect 18279 7157 18291 7191
rect 18233 7151 18291 7157
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 4614 6944 4620 6996
rect 4672 6984 4678 6996
rect 5074 6984 5080 6996
rect 4672 6956 5080 6984
rect 4672 6944 4678 6956
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 6604 6956 6653 6984
rect 6604 6944 6610 6956
rect 6641 6953 6653 6956
rect 6687 6953 6699 6987
rect 6641 6947 6699 6953
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 1302 6876 1308 6928
rect 1360 6916 1366 6928
rect 7116 6916 7144 6947
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8846 6984 8852 6996
rect 7800 6956 8852 6984
rect 7800 6944 7806 6956
rect 8846 6944 8852 6956
rect 8904 6984 8910 6996
rect 8904 6956 10732 6984
rect 8904 6944 8910 6956
rect 9582 6916 9588 6928
rect 1360 6888 7144 6916
rect 8036 6888 9588 6916
rect 1360 6876 1366 6888
rect 1670 6848 1676 6860
rect 1631 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2498 6857 2504 6860
rect 2492 6848 2504 6857
rect 1912 6820 2504 6848
rect 1912 6808 1918 6820
rect 2492 6811 2504 6820
rect 2498 6808 2504 6811
rect 2556 6808 2562 6860
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 4614 6848 4620 6860
rect 3108 6820 3280 6848
rect 4575 6820 4620 6848
rect 3108 6808 3114 6820
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1636 6752 2237 6780
rect 1636 6740 1642 6752
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 3252 6712 3280 6820
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 5224 6820 5273 6848
rect 5224 6808 5230 6820
rect 5261 6817 5273 6820
rect 5307 6817 5319 6851
rect 5261 6811 5319 6817
rect 5528 6851 5586 6857
rect 5528 6817 5540 6851
rect 5574 6848 5586 6851
rect 6086 6848 6092 6860
rect 5574 6820 6092 6848
rect 5574 6817 5586 6820
rect 5528 6811 5586 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6914 6848 6920 6860
rect 6875 6820 6920 6848
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 8036 6848 8064 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 10704 6925 10732 6956
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11701 6987 11759 6993
rect 11701 6984 11713 6987
rect 11112 6956 11713 6984
rect 11112 6944 11118 6956
rect 11701 6953 11713 6956
rect 11747 6953 11759 6987
rect 11701 6947 11759 6953
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 12308 6956 13737 6984
rect 12308 6944 12314 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 14553 6987 14611 6993
rect 14553 6953 14565 6987
rect 14599 6984 14611 6987
rect 15654 6984 15660 6996
rect 14599 6956 15660 6984
rect 14599 6953 14611 6956
rect 14553 6947 14611 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 17037 6987 17095 6993
rect 17037 6953 17049 6987
rect 17083 6984 17095 6987
rect 17218 6984 17224 6996
rect 17083 6956 17224 6984
rect 17083 6953 17095 6956
rect 17037 6947 17095 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17681 6987 17739 6993
rect 17681 6953 17693 6987
rect 17727 6984 17739 6987
rect 17770 6984 17776 6996
rect 17727 6956 17776 6984
rect 17727 6953 17739 6956
rect 17681 6947 17739 6953
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 10689 6919 10747 6925
rect 10689 6885 10701 6919
rect 10735 6916 10747 6919
rect 11882 6916 11888 6928
rect 10735 6888 11888 6916
rect 10735 6885 10747 6888
rect 10689 6879 10747 6885
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 11974 6876 11980 6928
rect 12032 6916 12038 6928
rect 13170 6916 13176 6928
rect 12032 6888 13176 6916
rect 12032 6876 12038 6888
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 17494 6916 17500 6928
rect 14332 6888 17500 6916
rect 14332 6876 14338 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 7699 6820 8064 6848
rect 8104 6851 8162 6857
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8104 6817 8116 6851
rect 8150 6848 8162 6851
rect 8570 6848 8576 6860
rect 8150 6820 8576 6848
rect 8150 6817 8162 6820
rect 8104 6811 8162 6817
rect 8570 6808 8576 6820
rect 8628 6848 8634 6860
rect 8628 6820 8892 6848
rect 8628 6808 8634 6820
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 7466 6780 7472 6792
rect 6328 6752 7472 6780
rect 6328 6740 6334 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8864 6780 8892 6820
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 8996 6820 9689 6848
rect 8996 6808 9002 6820
rect 9677 6817 9689 6820
rect 9723 6848 9735 6851
rect 9858 6848 9864 6860
rect 9723 6820 9864 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 12601 6851 12659 6857
rect 12601 6848 12613 6851
rect 11716 6820 12613 6848
rect 11716 6792 11744 6820
rect 12601 6817 12613 6820
rect 12647 6817 12659 6851
rect 12601 6811 12659 6817
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 12952 6820 13400 6848
rect 12952 6808 12958 6820
rect 9766 6780 9772 6792
rect 8864 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11698 6780 11704 6792
rect 11011 6752 11704 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12250 6780 12256 6792
rect 12023 6752 12256 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 3605 6715 3663 6721
rect 3605 6712 3617 6715
rect 3252 6684 3617 6712
rect 3605 6681 3617 6684
rect 3651 6712 3663 6715
rect 3694 6712 3700 6724
rect 3651 6684 3700 6712
rect 3651 6681 3663 6684
rect 3605 6675 3663 6681
rect 3694 6672 3700 6684
rect 3752 6672 3758 6724
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 9861 6715 9919 6721
rect 9861 6712 9873 6715
rect 3844 6684 4384 6712
rect 3844 6672 3850 6684
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2866 6644 2872 6656
rect 1903 6616 2872 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 4246 6644 4252 6656
rect 4207 6616 4252 6644
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4356 6644 4384 6684
rect 6288 6684 7604 6712
rect 6288 6644 6316 6684
rect 4356 6616 6316 6644
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 7432 6616 7481 6644
rect 7432 6604 7438 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7576 6644 7604 6684
rect 8772 6684 9873 6712
rect 8772 6644 8800 6684
rect 9861 6681 9873 6684
rect 9907 6681 9919 6715
rect 9861 6675 9919 6681
rect 10321 6715 10379 6721
rect 10321 6681 10333 6715
rect 10367 6712 10379 6715
rect 11808 6712 11836 6743
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6749 12403 6783
rect 13372 6780 13400 6820
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 15562 6848 15568 6860
rect 13596 6820 15568 6848
rect 13596 6808 13602 6820
rect 15562 6808 15568 6820
rect 15620 6848 15626 6860
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 15620 6820 15669 6848
rect 15620 6808 15626 6820
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 15913 6851 15971 6857
rect 15913 6848 15925 6851
rect 15804 6820 15925 6848
rect 15804 6808 15810 6820
rect 15913 6817 15925 6820
rect 15959 6817 15971 6851
rect 15913 6811 15971 6817
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 17954 6848 17960 6860
rect 16264 6820 17960 6848
rect 16264 6808 16270 6820
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 13372 6752 14657 6780
rect 12345 6743 12403 6749
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14826 6780 14832 6792
rect 14787 6752 14832 6780
rect 14645 6743 14703 6749
rect 10367 6684 11836 6712
rect 10367 6681 10379 6684
rect 10321 6675 10379 6681
rect 7576 6616 8800 6644
rect 7469 6607 7527 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 9088 6616 9229 6644
rect 9088 6604 9094 6616
rect 9217 6613 9229 6616
rect 9263 6644 9275 6647
rect 10226 6644 10232 6656
rect 9263 6616 10232 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11296 6616 11345 6644
rect 11296 6604 11302 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 12360 6644 12388 6743
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 14660 6712 14688 6743
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17552 6752 17785 6780
rect 17552 6740 17558 6752
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 15470 6712 15476 6724
rect 14056 6684 14504 6712
rect 14660 6684 15476 6712
rect 14056 6672 14062 6684
rect 13538 6644 13544 6656
rect 12360 6616 13544 6644
rect 11333 6607 11391 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14366 6644 14372 6656
rect 14231 6616 14372 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14476 6644 14504 6684
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 17126 6672 17132 6724
rect 17184 6712 17190 6724
rect 17880 6712 17908 6743
rect 17184 6684 17908 6712
rect 17184 6672 17190 6684
rect 15378 6644 15384 6656
rect 14476 6616 15384 6644
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 17313 6647 17371 6653
rect 17313 6613 17325 6647
rect 17359 6644 17371 6647
rect 17402 6644 17408 6656
rect 17359 6616 17408 6644
rect 17359 6613 17371 6616
rect 17313 6607 17371 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2958 6440 2964 6452
rect 1728 6412 2964 6440
rect 1728 6400 1734 6412
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4890 6400 4896 6452
rect 4948 6440 4954 6452
rect 6086 6440 6092 6452
rect 4948 6412 5672 6440
rect 6047 6412 6092 6440
rect 4948 6400 4954 6412
rect 3050 6372 3056 6384
rect 2608 6344 3056 6372
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 1664 6239 1722 6245
rect 1664 6205 1676 6239
rect 1710 6236 1722 6239
rect 2608 6236 2636 6344
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 5644 6372 5672 6412
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 6972 6412 11652 6440
rect 6972 6400 6978 6412
rect 8570 6372 8576 6384
rect 5644 6344 8576 6372
rect 8570 6332 8576 6344
rect 8628 6332 8634 6384
rect 11624 6372 11652 6412
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 11756 6412 12081 6440
rect 11756 6400 11762 6412
rect 12069 6409 12081 6412
rect 12115 6409 12127 6443
rect 12069 6403 12127 6409
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 12710 6440 12716 6452
rect 12483 6412 12716 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 11974 6372 11980 6384
rect 11624 6344 11980 6372
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 3694 6304 3700 6316
rect 3655 6276 3700 6304
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6362 6304 6368 6316
rect 5776 6276 6368 6304
rect 5776 6264 5782 6276
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 6472 6276 7665 6304
rect 1710 6208 2636 6236
rect 1710 6205 1722 6208
rect 1664 6199 1722 6205
rect 1412 6168 1440 6199
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3568 6208 4077 6236
rect 3568 6196 3574 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 4976 6239 5034 6245
rect 4976 6205 4988 6239
rect 5022 6236 5034 6239
rect 6472 6236 6500 6276
rect 7653 6273 7665 6276
rect 7699 6304 7711 6307
rect 8202 6304 8208 6316
rect 7699 6276 8208 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 12084 6304 12112 6403
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 12912 6412 18092 6440
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 12912 6372 12940 6412
rect 12308 6344 12940 6372
rect 12308 6332 12314 6344
rect 12912 6313 12940 6344
rect 13633 6375 13691 6381
rect 13633 6341 13645 6375
rect 13679 6372 13691 6375
rect 15102 6372 15108 6384
rect 13679 6344 15108 6372
rect 13679 6341 13691 6344
rect 13633 6335 13691 6341
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 15562 6332 15568 6384
rect 15620 6372 15626 6384
rect 16025 6375 16083 6381
rect 16025 6372 16037 6375
rect 15620 6344 16037 6372
rect 15620 6332 15626 6344
rect 16025 6341 16037 6344
rect 16071 6341 16083 6375
rect 16025 6335 16083 6341
rect 12897 6307 12955 6313
rect 8588 6276 8800 6304
rect 12084 6276 12848 6304
rect 5022 6208 6500 6236
rect 6549 6239 6607 6245
rect 5022 6205 5034 6208
rect 4976 6199 5034 6205
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 7374 6236 7380 6248
rect 6595 6208 7380 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 1578 6168 1584 6180
rect 1412 6140 1584 6168
rect 1578 6128 1584 6140
rect 1636 6128 1642 6180
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 2222 6168 2228 6180
rect 1912 6140 2228 6168
rect 1912 6128 1918 6140
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 4724 6168 4752 6199
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7524 6208 8125 6236
rect 7524 6196 7530 6208
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8588 6236 8616 6276
rect 8159 6208 8616 6236
rect 8665 6239 8723 6245
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8772 6236 8800 6276
rect 8772 6208 9168 6236
rect 8665 6199 8723 6205
rect 5166 6168 5172 6180
rect 4028 6140 4384 6168
rect 4724 6140 5172 6168
rect 4028 6128 4034 6140
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 2777 6103 2835 6109
rect 2777 6100 2789 6103
rect 2740 6072 2789 6100
rect 2740 6060 2746 6072
rect 2777 6069 2789 6072
rect 2823 6069 2835 6103
rect 3050 6100 3056 6112
rect 3011 6072 3056 6100
rect 2777 6063 2835 6069
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3421 6103 3479 6109
rect 3421 6100 3433 6103
rect 3384 6072 3433 6100
rect 3384 6060 3390 6072
rect 3421 6069 3433 6072
rect 3467 6069 3479 6103
rect 3421 6063 3479 6069
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 4246 6100 4252 6112
rect 3568 6072 3613 6100
rect 4207 6072 4252 6100
rect 3568 6060 3574 6072
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4356 6100 4384 6140
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 6270 6168 6276 6180
rect 5276 6140 6276 6168
rect 5276 6100 5304 6140
rect 6270 6128 6276 6140
rect 6328 6128 6334 6180
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 7834 6168 7840 6180
rect 6788 6140 7840 6168
rect 6788 6128 6794 6140
rect 7834 6128 7840 6140
rect 7892 6168 7898 6180
rect 8478 6168 8484 6180
rect 7892 6140 8484 6168
rect 7892 6128 7898 6140
rect 8478 6128 8484 6140
rect 8536 6168 8542 6180
rect 8680 6168 8708 6199
rect 8536 6140 8708 6168
rect 8932 6171 8990 6177
rect 8536 6128 8542 6140
rect 8932 6137 8944 6171
rect 8978 6168 8990 6171
rect 9030 6168 9036 6180
rect 8978 6140 9036 6168
rect 8978 6137 8990 6140
rect 8932 6131 8990 6137
rect 9030 6128 9036 6140
rect 9088 6128 9094 6180
rect 9140 6168 9168 6208
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 10376 6208 10701 6236
rect 10376 6196 10382 6208
rect 10689 6205 10701 6208
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12434 6236 12440 6248
rect 12032 6208 12440 6236
rect 12032 6196 12038 6208
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12820 6236 12848 6276
rect 12897 6273 12909 6307
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13004 6236 13032 6267
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 14645 6307 14703 6313
rect 13228 6276 14504 6304
rect 13228 6264 13234 6276
rect 12820 6208 13032 6236
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 13412 6208 13461 6236
rect 13412 6196 13418 6208
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 13998 6236 14004 6248
rect 13449 6199 13507 6205
rect 13924 6208 14004 6236
rect 9140 6140 9260 6168
rect 9232 6112 9260 6140
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 10956 6171 11014 6177
rect 9364 6140 10180 6168
rect 9364 6128 9370 6140
rect 6362 6100 6368 6112
rect 4356 6072 5304 6100
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 7101 6103 7159 6109
rect 7101 6100 7113 6103
rect 6512 6072 7113 6100
rect 6512 6060 6518 6072
rect 7101 6069 7113 6072
rect 7147 6069 7159 6103
rect 7466 6100 7472 6112
rect 7427 6072 7472 6100
rect 7101 6063 7159 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8294 6100 8300 6112
rect 7616 6072 7661 6100
rect 8255 6072 8300 6100
rect 7616 6060 7622 6072
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 9122 6100 9128 6112
rect 8444 6072 9128 6100
rect 8444 6060 8450 6072
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9214 6060 9220 6112
rect 9272 6060 9278 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9824 6072 10057 6100
rect 9824 6060 9830 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10152 6100 10180 6140
rect 10956 6137 10968 6171
rect 11002 6168 11014 6171
rect 11790 6168 11796 6180
rect 11002 6140 11796 6168
rect 11002 6137 11014 6140
rect 10956 6131 11014 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 10152 6072 12817 6100
rect 10045 6063 10103 6069
rect 12805 6069 12817 6072
rect 12851 6100 12863 6103
rect 13630 6100 13636 6112
rect 12851 6072 13636 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13630 6060 13636 6072
rect 13688 6100 13694 6112
rect 13924 6100 13952 6208
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14366 6236 14372 6248
rect 14327 6208 14372 6236
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 14476 6236 14504 6276
rect 14645 6273 14657 6307
rect 14691 6304 14703 6307
rect 15470 6304 15476 6316
rect 14691 6276 15476 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 15654 6304 15660 6316
rect 15615 6276 15660 6304
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16040 6304 16068 6335
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 16040 6276 16313 6304
rect 16301 6273 16313 6276
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 16209 6239 16267 6245
rect 16209 6236 16221 6239
rect 14476 6208 16221 6236
rect 16209 6205 16221 6208
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 16568 6239 16626 6245
rect 16568 6205 16580 6239
rect 16614 6236 16626 6239
rect 17126 6236 17132 6248
rect 16614 6208 17132 6236
rect 16614 6205 16626 6208
rect 16568 6199 16626 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 18064 6245 18092 6412
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 15381 6171 15439 6177
rect 15381 6168 15393 6171
rect 14016 6140 15393 6168
rect 14016 6109 14044 6140
rect 15381 6137 15393 6140
rect 15427 6137 15439 6171
rect 15381 6131 15439 6137
rect 15473 6171 15531 6177
rect 15473 6137 15485 6171
rect 15519 6168 15531 6171
rect 15519 6140 16528 6168
rect 15519 6137 15531 6140
rect 15473 6131 15531 6137
rect 13688 6072 13952 6100
rect 14001 6103 14059 6109
rect 13688 6060 13694 6072
rect 14001 6069 14013 6103
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 14182 6060 14188 6112
rect 14240 6100 14246 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 14240 6072 14473 6100
rect 14240 6060 14246 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 14700 6072 15025 6100
rect 14700 6060 14706 6072
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 16500 6100 16528 6140
rect 16666 6100 16672 6112
rect 16500 6072 16672 6100
rect 15013 6063 15071 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 17678 6100 17684 6112
rect 17639 6072 17684 6100
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 17828 6072 18245 6100
rect 17828 6060 17834 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 18233 6063 18291 6069
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 2501 5899 2559 5905
rect 2501 5896 2513 5899
rect 1544 5868 2513 5896
rect 1544 5856 1550 5868
rect 2501 5865 2513 5868
rect 2547 5865 2559 5899
rect 2501 5859 2559 5865
rect 2593 5899 2651 5905
rect 2593 5865 2605 5899
rect 2639 5896 2651 5899
rect 3050 5896 3056 5908
rect 2639 5868 3056 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4614 5896 4620 5908
rect 4479 5868 4620 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5626 5896 5632 5908
rect 4724 5868 5632 5896
rect 2958 5788 2964 5840
rect 3016 5828 3022 5840
rect 4724 5828 4752 5868
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 5905 5899 5963 5905
rect 5905 5865 5917 5899
rect 5951 5896 5963 5899
rect 6454 5896 6460 5908
rect 5951 5868 6460 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 7524 5868 8493 5896
rect 7524 5856 7530 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8812 5868 8861 5896
rect 8812 5856 8818 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 11606 5896 11612 5908
rect 9272 5868 11612 5896
rect 9272 5856 9278 5868
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 11790 5896 11796 5908
rect 11747 5868 11796 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 12437 5899 12495 5905
rect 12437 5865 12449 5899
rect 12483 5896 12495 5899
rect 12618 5896 12624 5908
rect 12483 5868 12624 5896
rect 12483 5865 12495 5868
rect 12437 5859 12495 5865
rect 12618 5856 12624 5868
rect 12676 5896 12682 5908
rect 13170 5896 13176 5908
rect 12676 5868 13176 5896
rect 12676 5856 12682 5868
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14274 5856 14280 5908
rect 14332 5896 14338 5908
rect 14553 5899 14611 5905
rect 14553 5896 14565 5899
rect 14332 5868 14565 5896
rect 14332 5856 14338 5868
rect 14553 5865 14565 5868
rect 14599 5896 14611 5899
rect 14734 5896 14740 5908
rect 14599 5868 14740 5896
rect 14599 5865 14611 5868
rect 14553 5859 14611 5865
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 15712 5868 16681 5896
rect 15712 5856 15718 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 16669 5859 16727 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 3016 5800 4752 5828
rect 4801 5831 4859 5837
rect 3016 5788 3022 5800
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 4847 5800 9873 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 9861 5797 9873 5800
rect 9907 5797 9919 5831
rect 13906 5828 13912 5840
rect 9861 5791 9919 5797
rect 10520 5800 11744 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 2130 5760 2136 5772
rect 1719 5732 2136 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 1412 5624 1440 5723
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 3694 5760 3700 5772
rect 3283 5732 3700 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 5810 5760 5816 5772
rect 4939 5732 5672 5760
rect 5771 5732 5816 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 2682 5692 2688 5704
rect 2643 5664 2688 5692
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 3016 5664 3433 5692
rect 3016 5652 3022 5664
rect 3421 5661 3433 5664
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 5442 5692 5448 5704
rect 5123 5664 5448 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5644 5692 5672 5732
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 6178 5760 6184 5772
rect 5920 5732 6184 5760
rect 5920 5692 5948 5732
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 6362 5720 6368 5772
rect 6420 5760 6426 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6420 5732 6745 5760
rect 6420 5720 6426 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7092 5763 7150 5769
rect 7092 5760 7104 5763
rect 6972 5732 7104 5760
rect 6972 5720 6978 5732
rect 7092 5729 7104 5732
rect 7138 5760 7150 5763
rect 7138 5732 8340 5760
rect 7138 5729 7150 5732
rect 7092 5723 7150 5729
rect 6086 5692 6092 5704
rect 5644 5664 5948 5692
rect 6047 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 2133 5627 2191 5633
rect 2133 5624 2145 5627
rect 1412 5596 2145 5624
rect 2133 5593 2145 5596
rect 2179 5593 2191 5627
rect 2133 5587 2191 5593
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 8202 5624 8208 5636
rect 4396 5596 6868 5624
rect 8163 5596 8208 5624
rect 4396 5584 4402 5596
rect 2498 5516 2504 5568
rect 2556 5556 2562 5568
rect 2774 5556 2780 5568
rect 2556 5528 2780 5556
rect 2556 5516 2562 5528
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 4764 5528 5457 5556
rect 4764 5516 4770 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5445 5519 5503 5525
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 6270 5556 6276 5568
rect 5776 5528 6276 5556
rect 5776 5516 5782 5528
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6549 5559 6607 5565
rect 6549 5525 6561 5559
rect 6595 5556 6607 5559
rect 6730 5556 6736 5568
rect 6595 5528 6736 5556
rect 6595 5525 6607 5528
rect 6549 5519 6607 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 6840 5556 6868 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8312 5624 8340 5732
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 10520 5760 10548 5800
rect 8444 5732 10548 5760
rect 10588 5763 10646 5769
rect 8444 5720 8450 5732
rect 10588 5729 10600 5763
rect 10634 5760 10646 5763
rect 10634 5732 11652 5760
rect 10634 5729 10646 5732
rect 10588 5723 10646 5729
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8812 5664 8953 5692
rect 8812 5652 8818 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 10318 5692 10324 5704
rect 10279 5664 10324 5692
rect 9033 5655 9091 5661
rect 8478 5624 8484 5636
rect 8312 5596 8484 5624
rect 8478 5584 8484 5596
rect 8536 5624 8542 5636
rect 9048 5624 9076 5655
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 8536 5596 9076 5624
rect 8536 5584 8542 5596
rect 9214 5584 9220 5636
rect 9272 5624 9278 5636
rect 11624 5624 11652 5732
rect 11716 5692 11744 5800
rect 12636 5800 13912 5828
rect 12636 5769 12664 5800
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 14090 5788 14096 5840
rect 14148 5828 14154 5840
rect 14645 5831 14703 5837
rect 14645 5828 14657 5831
rect 14148 5800 14657 5828
rect 14148 5788 14154 5800
rect 14645 5797 14657 5800
rect 14691 5797 14703 5831
rect 14645 5791 14703 5797
rect 15470 5788 15476 5840
rect 15528 5837 15534 5840
rect 15528 5831 15592 5837
rect 15528 5797 15546 5831
rect 15580 5828 15592 5831
rect 16390 5828 16396 5840
rect 15580 5800 16396 5828
rect 15580 5797 15592 5800
rect 15528 5791 15592 5797
rect 15528 5788 15534 5791
rect 16390 5788 16396 5800
rect 16448 5788 16454 5840
rect 17310 5828 17316 5840
rect 17271 5800 17316 5828
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 12621 5763 12679 5769
rect 12621 5729 12633 5763
rect 12667 5729 12679 5763
rect 13170 5760 13176 5772
rect 13131 5732 13176 5760
rect 12621 5723 12679 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 17954 5760 17960 5772
rect 14844 5732 16344 5760
rect 17915 5732 17960 5760
rect 14844 5704 14872 5732
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11716 5664 11989 5692
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 11977 5655 12035 5661
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5661 13415 5695
rect 14826 5692 14832 5704
rect 14787 5664 14832 5692
rect 13357 5655 13415 5661
rect 12526 5624 12532 5636
rect 9272 5596 10364 5624
rect 11624 5596 12532 5624
rect 9272 5584 9278 5596
rect 9582 5556 9588 5568
rect 6840 5528 9588 5556
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10336 5556 10364 5596
rect 12526 5584 12532 5596
rect 12584 5624 12590 5636
rect 13372 5624 13400 5655
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 16316 5692 16344 5732
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 16316 5664 17509 5692
rect 15289 5655 15347 5661
rect 17497 5661 17509 5664
rect 17543 5692 17555 5695
rect 17678 5692 17684 5704
rect 17543 5664 17684 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 13814 5624 13820 5636
rect 12584 5596 13820 5624
rect 12584 5584 12590 5596
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 12250 5556 12256 5568
rect 10336 5528 12256 5556
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12400 5528 12817 5556
rect 12400 5516 12406 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 15010 5516 15016 5568
rect 15068 5556 15074 5568
rect 15304 5556 15332 5655
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 15562 5556 15568 5568
rect 15068 5528 15568 5556
rect 15068 5516 15074 5528
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 16942 5556 16948 5568
rect 16903 5528 16948 5556
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18141 5559 18199 5565
rect 18141 5556 18153 5559
rect 17920 5528 18153 5556
rect 17920 5516 17926 5528
rect 18141 5525 18153 5528
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 5718 5352 5724 5364
rect 4755 5324 5724 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 5868 5324 6837 5352
rect 5868 5312 5874 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 11514 5352 11520 5364
rect 6825 5315 6883 5321
rect 8312 5324 11520 5352
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 3620 5256 4016 5284
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 3620 5148 3648 5256
rect 3786 5216 3792 5228
rect 3747 5188 3792 5216
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 3697 5151 3755 5157
rect 3697 5148 3709 5151
rect 2648 5120 3709 5148
rect 2648 5108 2654 5120
rect 3697 5117 3709 5120
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 3878 5108 3884 5160
rect 3936 5108 3942 5160
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 1826 5083 1884 5089
rect 1826 5080 1838 5083
rect 1728 5052 1838 5080
rect 1728 5040 1734 5052
rect 1826 5049 1838 5052
rect 1872 5049 1884 5083
rect 1826 5043 1884 5049
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5080 3663 5083
rect 3896 5080 3924 5108
rect 3651 5052 3924 5080
rect 3988 5080 4016 5256
rect 4264 5256 5549 5284
rect 4264 5225 4292 5256
rect 5537 5253 5549 5256
rect 5583 5253 5595 5287
rect 5537 5247 5595 5253
rect 5644 5256 7420 5284
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 5644 5216 5672 5256
rect 5399 5188 5672 5216
rect 6181 5219 6239 5225
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6270 5216 6276 5228
rect 6227 5188 6276 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 6914 5216 6920 5228
rect 6411 5188 6920 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 5537 5151 5595 5157
rect 4120 5120 5304 5148
rect 4120 5108 4126 5120
rect 5169 5083 5227 5089
rect 5169 5080 5181 5083
rect 3988 5052 5181 5080
rect 3651 5049 3663 5052
rect 3605 5043 3663 5049
rect 5169 5049 5181 5052
rect 5215 5049 5227 5083
rect 5276 5080 5304 5120
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5810 5148 5816 5160
rect 5583 5120 5816 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 7392 5148 7420 5256
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 8202 5216 8208 5228
rect 7515 5188 8208 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8312 5225 8340 5324
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14645 5355 14703 5361
rect 14645 5321 14657 5355
rect 14691 5352 14703 5355
rect 15194 5352 15200 5364
rect 14691 5324 15200 5352
rect 14691 5321 14703 5324
rect 14645 5315 14703 5321
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 16390 5352 16396 5364
rect 16351 5324 16396 5352
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 12434 5284 12440 5296
rect 11440 5256 12440 5284
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8536 5188 8581 5216
rect 8536 5176 8542 5188
rect 8846 5148 8852 5160
rect 7392 5120 8340 5148
rect 8807 5120 8852 5148
rect 5626 5080 5632 5092
rect 5276 5052 5632 5080
rect 5169 5043 5227 5049
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 6086 5080 6092 5092
rect 6047 5052 6092 5080
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 7650 5040 7656 5092
rect 7708 5080 7714 5092
rect 8202 5080 8208 5092
rect 7708 5052 8208 5080
rect 7708 5040 7714 5052
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 8312 5080 8340 5120
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 10318 5148 10324 5160
rect 9539 5120 10324 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 10318 5108 10324 5120
rect 10376 5148 10382 5160
rect 11440 5148 11468 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 16408 5284 16436 5312
rect 16408 5256 17264 5284
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11848 5188 11897 5216
rect 11848 5176 11854 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 13780 5188 14504 5216
rect 13780 5176 13786 5188
rect 10376 5120 11468 5148
rect 11701 5151 11759 5157
rect 10376 5108 10382 5120
rect 11701 5117 11713 5151
rect 11747 5148 11759 5151
rect 12342 5148 12348 5160
rect 11747 5120 12348 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12434 5108 12440 5160
rect 12492 5157 12498 5160
rect 14476 5157 14504 5188
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 14884 5188 15148 5216
rect 14884 5176 14890 5188
rect 12492 5148 12502 5157
rect 14461 5151 14519 5157
rect 12492 5120 12537 5148
rect 12492 5111 12502 5120
rect 14461 5117 14473 5151
rect 14507 5117 14519 5151
rect 15010 5148 15016 5160
rect 14971 5120 15016 5148
rect 14461 5111 14519 5117
rect 12492 5108 12498 5111
rect 15010 5108 15016 5120
rect 15068 5108 15074 5160
rect 15120 5148 15148 5188
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 16850 5216 16856 5228
rect 16724 5188 16856 5216
rect 16724 5176 16730 5188
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17236 5225 17264 5256
rect 17129 5219 17187 5225
rect 17129 5216 17141 5219
rect 17000 5188 17141 5216
rect 17000 5176 17006 5188
rect 17129 5185 17141 5188
rect 17175 5185 17187 5219
rect 17129 5179 17187 5185
rect 17221 5219 17279 5225
rect 17221 5185 17233 5219
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 15269 5151 15327 5157
rect 15269 5148 15281 5151
rect 15120 5120 15281 5148
rect 15269 5117 15281 5120
rect 15315 5117 15327 5151
rect 15269 5111 15327 5117
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17368 5120 18061 5148
rect 17368 5108 17374 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 9766 5089 9772 5092
rect 9738 5083 9772 5089
rect 9738 5080 9750 5083
rect 8312 5052 9750 5080
rect 9738 5049 9750 5052
rect 9824 5080 9830 5092
rect 9824 5052 9886 5080
rect 9738 5043 9772 5049
rect 9766 5040 9772 5043
rect 9824 5040 9830 5052
rect 12066 5040 12072 5092
rect 12124 5080 12130 5092
rect 12682 5083 12740 5089
rect 12682 5080 12694 5083
rect 12124 5052 12694 5080
rect 12124 5040 12130 5052
rect 12682 5049 12694 5052
rect 12728 5080 12740 5083
rect 13998 5080 14004 5092
rect 12728 5052 14004 5080
rect 12728 5049 12740 5052
rect 12682 5043 12740 5049
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2961 5015 3019 5021
rect 2961 5012 2973 5015
rect 2464 4984 2973 5012
rect 2464 4972 2470 4984
rect 2961 4981 2973 4984
rect 3007 4981 3019 5015
rect 3234 5012 3240 5024
rect 3195 4984 3240 5012
rect 2961 4975 3019 4981
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4798 5012 4804 5024
rect 3936 4984 4804 5012
rect 3936 4972 3942 4984
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 4948 4984 5089 5012
rect 4948 4972 4954 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5077 4975 5135 4981
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 5767 4984 7205 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7331 4984 7849 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 7837 4975 7895 4981
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 8720 4984 9045 5012
rect 8720 4972 8726 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 10686 5012 10692 5024
rect 9180 4984 10692 5012
rect 9180 4972 9186 4984
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 10870 5012 10876 5024
rect 10831 4984 10876 5012
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11333 5015 11391 5021
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 11606 5012 11612 5024
rect 11379 4984 11612 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 11848 4984 11893 5012
rect 11848 4972 11854 4984
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 15746 5012 15752 5024
rect 12032 4984 15752 5012
rect 12032 4972 12038 4984
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16816 4984 17049 5012
rect 16816 4972 16822 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 17037 4975 17095 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 3292 4780 4629 4808
rect 3292 4768 3298 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 6362 4808 6368 4820
rect 4617 4771 4675 4777
rect 5276 4780 6368 4808
rect 2124 4743 2182 4749
rect 2124 4709 2136 4743
rect 2170 4740 2182 4743
rect 2682 4740 2688 4752
rect 2170 4712 2688 4740
rect 2170 4709 2182 4712
rect 2124 4703 2182 4709
rect 2682 4700 2688 4712
rect 2740 4700 2746 4752
rect 5276 4740 5304 4780
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 8757 4811 8815 4817
rect 8757 4808 8769 4811
rect 8536 4780 8769 4808
rect 8536 4768 8542 4780
rect 8757 4777 8769 4780
rect 8803 4777 8815 4811
rect 8757 4771 8815 4777
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 10045 4811 10103 4817
rect 10045 4808 10057 4811
rect 9640 4780 10057 4808
rect 9640 4768 9646 4780
rect 10045 4777 10057 4780
rect 10091 4777 10103 4811
rect 10045 4771 10103 4777
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10410 4808 10416 4820
rect 10183 4780 10416 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 11149 4811 11207 4817
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 11422 4808 11428 4820
rect 11195 4780 11428 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12158 4808 12164 4820
rect 12119 4780 12164 4808
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12710 4808 12716 4820
rect 12492 4780 12716 4808
rect 12492 4768 12498 4780
rect 12710 4768 12716 4780
rect 12768 4808 12774 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12768 4780 12817 4808
rect 12768 4768 12774 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 13228 4780 13461 4808
rect 13228 4768 13234 4780
rect 13449 4777 13461 4780
rect 13495 4777 13507 4811
rect 13449 4771 13507 4777
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 15378 4808 15384 4820
rect 15335 4780 15384 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 16114 4808 16120 4820
rect 15488 4780 16120 4808
rect 3804 4712 5304 4740
rect 3804 4681 3832 4712
rect 5350 4700 5356 4752
rect 5408 4749 5414 4752
rect 5408 4743 5472 4749
rect 5408 4709 5426 4743
rect 5460 4709 5472 4743
rect 5408 4703 5472 4709
rect 5408 4700 5414 4703
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 8294 4740 8300 4752
rect 7484 4712 8300 4740
rect 3789 4675 3847 4681
rect 3789 4641 3801 4675
rect 3835 4641 3847 4675
rect 3789 4635 3847 4641
rect 4525 4675 4583 4681
rect 4525 4641 4537 4675
rect 4571 4672 4583 4675
rect 4614 4672 4620 4684
rect 4571 4644 4620 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 5368 4672 5396 4700
rect 4816 4644 5396 4672
rect 5644 4672 5672 4700
rect 5644 4644 6224 4672
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 4816 4613 4844 4644
rect 1857 4607 1915 4613
rect 1857 4604 1869 4607
rect 1636 4576 1869 4604
rect 1636 4564 1642 4576
rect 1857 4573 1869 4576
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4573 4859 4607
rect 5166 4604 5172 4616
rect 5127 4576 5172 4604
rect 4801 4567 4859 4573
rect 1872 4468 1900 4567
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 6196 4604 6224 4644
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 6604 4644 6837 4672
rect 6604 4632 6610 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 7484 4672 7512 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 11241 4743 11299 4749
rect 11241 4709 11253 4743
rect 11287 4740 11299 4743
rect 12894 4740 12900 4752
rect 11287 4712 12900 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 12894 4700 12900 4712
rect 12952 4700 12958 4752
rect 13906 4740 13912 4752
rect 13819 4712 13912 4740
rect 13906 4700 13912 4712
rect 13964 4740 13970 4752
rect 15488 4740 15516 4780
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 16758 4808 16764 4820
rect 16719 4780 16764 4808
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 17221 4811 17279 4817
rect 17221 4777 17233 4811
rect 17267 4808 17279 4811
rect 17589 4811 17647 4817
rect 17589 4808 17601 4811
rect 17267 4780 17601 4808
rect 17267 4777 17279 4780
rect 17221 4771 17279 4777
rect 17589 4777 17601 4780
rect 17635 4808 17647 4811
rect 18138 4808 18144 4820
rect 17635 4780 18144 4808
rect 17635 4777 17647 4780
rect 17589 4771 17647 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 15746 4740 15752 4752
rect 13964 4712 15516 4740
rect 15707 4712 15752 4740
rect 13964 4700 13970 4712
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 6825 4635 6883 4641
rect 6932 4644 7512 4672
rect 7644 4675 7702 4681
rect 6932 4604 6960 4644
rect 7644 4641 7656 4675
rect 7690 4672 7702 4675
rect 8202 4672 8208 4684
rect 7690 4644 8208 4672
rect 7690 4641 7702 4644
rect 7644 4635 7702 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8812 4644 9045 4672
rect 8812 4632 8818 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 9548 4644 12572 4672
rect 9548 4632 9554 4644
rect 6196 4576 6960 4604
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 7377 4567 7435 4573
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 3237 4539 3295 4545
rect 3237 4536 3249 4539
rect 3200 4508 3249 4536
rect 3200 4496 3206 4508
rect 3237 4505 3249 4508
rect 3283 4536 3295 4539
rect 3786 4536 3792 4548
rect 3283 4508 3792 4536
rect 3283 4505 3295 4508
rect 3237 4499 3295 4505
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 5184 4536 5212 4564
rect 4080 4508 5212 4536
rect 2590 4468 2596 4480
rect 1872 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4468 2654 4480
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 2648 4440 3617 4468
rect 2648 4428 2654 4440
rect 3605 4437 3617 4440
rect 3651 4468 3663 4471
rect 4080 4468 4108 4508
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7392 4536 7420 4567
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 11974 4604 11980 4616
rect 11471 4576 11980 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4573 12311 4607
rect 12434 4604 12440 4616
rect 12395 4576 12440 4604
rect 12253 4567 12311 4573
rect 6972 4508 7420 4536
rect 6972 4496 6978 4508
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 10686 4536 10692 4548
rect 8628 4508 10692 4536
rect 8628 4496 8634 4508
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4536 10839 4539
rect 12268 4536 12296 4567
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 12544 4604 12572 4644
rect 12618 4632 12624 4684
rect 12676 4672 12682 4684
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12676 4644 13001 4672
rect 12676 4632 12682 4644
rect 12989 4641 13001 4644
rect 13035 4641 13047 4675
rect 12989 4635 13047 4641
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4672 13875 4675
rect 14461 4675 14519 4681
rect 14461 4672 14473 4675
rect 13863 4644 14473 4672
rect 13863 4641 13875 4644
rect 13817 4635 13875 4641
rect 14461 4641 14473 4644
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14792 4644 15669 4672
rect 14792 4632 14798 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16172 4644 17141 4672
rect 16172 4632 16178 4644
rect 17129 4641 17141 4644
rect 17175 4641 17187 4675
rect 17770 4672 17776 4684
rect 17731 4644 17776 4672
rect 17129 4635 17187 4641
rect 17770 4632 17776 4644
rect 17828 4632 17834 4684
rect 13998 4604 14004 4616
rect 12544 4576 12664 4604
rect 13959 4576 14004 4604
rect 10827 4508 12296 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 3651 4440 4108 4468
rect 4157 4471 4215 4477
rect 3651 4437 3663 4440
rect 3605 4431 3663 4437
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 6086 4468 6092 4480
rect 4203 4440 6092 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6546 4468 6552 4480
rect 6507 4440 6552 4468
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 7006 4468 7012 4480
rect 6967 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 9214 4468 9220 4480
rect 9175 4440 9220 4468
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 9766 4468 9772 4480
rect 9723 4440 9772 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 12636 4468 12664 4576
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 17678 4604 17684 4616
rect 17451 4576 17684 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18506 4604 18512 4616
rect 18095 4576 18512 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 15194 4468 15200 4480
rect 12636 4440 15200 4468
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15378 4428 15384 4480
rect 15436 4468 15442 4480
rect 17589 4471 17647 4477
rect 17589 4468 17601 4471
rect 15436 4440 17601 4468
rect 15436 4428 15442 4440
rect 17589 4437 17601 4440
rect 17635 4437 17647 4471
rect 17589 4431 17647 4437
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 1210 4224 1216 4276
rect 1268 4264 1274 4276
rect 1268 4236 4200 4264
rect 1268 4224 1274 4236
rect 1670 4156 1676 4208
rect 1728 4196 1734 4208
rect 2774 4196 2780 4208
rect 1728 4168 2780 4196
rect 1728 4156 1734 4168
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2424 4137 2452 4168
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 2096 4100 2329 4128
rect 2096 4088 2102 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 2590 4088 2596 4140
rect 2648 4128 2654 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2648 4100 2881 4128
rect 2648 4088 2654 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 3142 4069 3148 4072
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 1912 4032 2237 4060
rect 1912 4020 1918 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 3136 4060 3148 4069
rect 3103 4032 3148 4060
rect 2225 4023 2283 4029
rect 3136 4023 3148 4032
rect 3142 4020 3148 4023
rect 3200 4020 3206 4072
rect 4172 4060 4200 4236
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 7006 4264 7012 4276
rect 4488 4236 7012 4264
rect 4488 4224 4494 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 8202 4264 8208 4276
rect 8163 4236 8208 4264
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 11333 4267 11391 4273
rect 11333 4233 11345 4267
rect 11379 4264 11391 4267
rect 12158 4264 12164 4276
rect 11379 4236 12164 4264
rect 11379 4233 11391 4236
rect 11333 4227 11391 4233
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 14645 4267 14703 4273
rect 14645 4264 14657 4267
rect 12952 4236 14657 4264
rect 12952 4224 12958 4236
rect 14645 4233 14657 4236
rect 14691 4233 14703 4267
rect 14645 4227 14703 4233
rect 15194 4224 15200 4276
rect 15252 4224 15258 4276
rect 16850 4264 16856 4276
rect 16811 4236 16856 4264
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 4249 4199 4307 4205
rect 4249 4165 4261 4199
rect 4295 4165 4307 4199
rect 5994 4196 6000 4208
rect 4249 4159 4307 4165
rect 5920 4168 6000 4196
rect 4264 4128 4292 4159
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 4264 4100 5273 4128
rect 5261 4097 5273 4100
rect 5307 4128 5319 4131
rect 5350 4128 5356 4140
rect 5307 4100 5356 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5920 4128 5948 4168
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 13998 4156 14004 4208
rect 14056 4196 14062 4208
rect 14369 4199 14427 4205
rect 14369 4196 14381 4199
rect 14056 4168 14381 4196
rect 14056 4156 14062 4168
rect 14369 4165 14381 4168
rect 14415 4165 14427 4199
rect 15212 4196 15240 4224
rect 17770 4196 17776 4208
rect 15212 4168 17776 4196
rect 14369 4159 14427 4165
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 6086 4128 6092 4140
rect 5644 4100 5948 4128
rect 6047 4100 6092 4128
rect 4890 4060 4896 4072
rect 4172 4032 4896 4060
rect 4890 4020 4896 4032
rect 4948 4060 4954 4072
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4948 4032 4997 4060
rect 4948 4020 4954 4032
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5644 4060 5672 4100
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6546 4128 6552 4140
rect 6227 4100 6552 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 5123 4032 5672 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6196 4060 6224 4091
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 11974 4128 11980 4140
rect 11935 4100 11980 4128
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12526 4128 12532 4140
rect 12084 4100 12532 4128
rect 5776 4032 6224 4060
rect 5776 4020 5782 4032
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4060 6883 4063
rect 6914 4060 6920 4072
rect 6871 4032 6920 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 6914 4020 6920 4032
rect 6972 4060 6978 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 6972 4032 8861 4060
rect 6972 4020 6978 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 9398 4060 9404 4072
rect 8849 4023 8907 4029
rect 8956 4032 9404 4060
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2682 3992 2688 4004
rect 2372 3964 2688 3992
rect 2372 3952 2378 3964
rect 2682 3952 2688 3964
rect 2740 3952 2746 4004
rect 5997 3995 6055 4001
rect 5997 3992 6009 3995
rect 4632 3964 6009 3992
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 4632 3933 4660 3964
rect 5997 3961 6009 3964
rect 6043 3961 6055 3995
rect 5997 3955 6055 3961
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6788 3964 7082 3992
rect 6788 3952 6794 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 8956 3992 8984 4032
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 9732 4032 10517 4060
rect 9732 4020 9738 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11204 4032 11713 4060
rect 11204 4020 11210 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 12084 4060 12112 4100
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12768 4100 13001 4128
rect 12768 4088 12774 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 12989 4091 13047 4097
rect 14016 4100 15209 4128
rect 11839 4032 12112 4060
rect 13256 4063 13314 4069
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 13256 4029 13268 4063
rect 13302 4060 13314 4063
rect 13814 4060 13820 4072
rect 13302 4032 13820 4060
rect 13302 4029 13314 4032
rect 13256 4023 13314 4029
rect 9122 4001 9128 4004
rect 7248 3964 8984 3992
rect 7248 3952 7254 3964
rect 9116 3955 9128 4001
rect 9180 3992 9186 4004
rect 9180 3964 9216 3992
rect 9122 3952 9128 3955
rect 9180 3952 9186 3964
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 9640 3964 10364 3992
rect 9640 3952 9646 3964
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 10226 3924 10232 3936
rect 5684 3896 5729 3924
rect 10187 3896 10232 3924
rect 5684 3884 5690 3896
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10336 3924 10364 3964
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 10781 3995 10839 4001
rect 10781 3992 10793 3995
rect 10468 3964 10793 3992
rect 10468 3952 10474 3964
rect 10781 3961 10793 3964
rect 10827 3961 10839 3995
rect 11716 3992 11744 4023
rect 13814 4020 13820 4032
rect 13872 4060 13878 4072
rect 14016 4060 14044 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 15197 4091 15255 4097
rect 16942 4088 16948 4140
rect 17000 4128 17006 4140
rect 17586 4128 17592 4140
rect 17000 4100 17592 4128
rect 17000 4088 17006 4100
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 13872 4032 14044 4060
rect 13872 4020 13878 4032
rect 14550 4020 14556 4072
rect 14608 4060 14614 4072
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14608 4032 15025 4060
rect 14608 4020 14614 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 16114 4060 16120 4072
rect 15620 4032 16120 4060
rect 15620 4020 15626 4032
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 16666 4060 16672 4072
rect 16627 4032 16672 4060
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 17221 4063 17279 4069
rect 17221 4029 17233 4063
rect 17267 4060 17279 4063
rect 17678 4060 17684 4072
rect 17267 4032 17684 4060
rect 17267 4029 17279 4032
rect 17221 4023 17279 4029
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 11974 3992 11980 4004
rect 11716 3964 11980 3992
rect 10781 3955 10839 3961
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 15105 3995 15163 4001
rect 15105 3992 15117 3995
rect 12084 3964 15117 3992
rect 11146 3924 11152 3936
rect 10336 3896 11152 3924
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 12084 3924 12112 3964
rect 15105 3961 15117 3964
rect 15151 3992 15163 3995
rect 17494 3992 17500 4004
rect 15151 3964 17500 3992
rect 15151 3961 15163 3964
rect 15105 3955 15163 3961
rect 17494 3952 17500 3964
rect 17552 3992 17558 4004
rect 18064 3992 18092 4023
rect 17552 3964 18092 3992
rect 17552 3952 17558 3964
rect 11388 3896 12112 3924
rect 11388 3884 11394 3896
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 16298 3924 16304 3936
rect 12492 3896 12537 3924
rect 16259 3896 16304 3924
rect 12492 3884 12498 3896
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 17402 3924 17408 3936
rect 17363 3896 17408 3924
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 2774 3720 2780 3732
rect 2735 3692 2780 3720
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 5721 3723 5779 3729
rect 4396 3692 5028 3720
rect 4396 3680 4402 3692
rect 4706 3652 4712 3664
rect 3252 3624 4712 3652
rect 382 3544 388 3596
rect 440 3584 446 3596
rect 3252 3593 3280 3624
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 5000 3652 5028 3692
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 6730 3720 6736 3732
rect 5767 3692 6736 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 6730 3680 6736 3692
rect 6788 3720 6794 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 6788 3692 7205 3720
rect 6788 3680 6794 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 7469 3723 7527 3729
rect 7469 3689 7481 3723
rect 7515 3720 7527 3723
rect 7558 3720 7564 3732
rect 7515 3692 7564 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 7975 3692 8493 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 8849 3723 8907 3729
rect 8849 3689 8861 3723
rect 8895 3720 8907 3723
rect 9306 3720 9312 3732
rect 8895 3692 9312 3720
rect 8895 3689 8907 3692
rect 8849 3683 8907 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3689 9919 3723
rect 9861 3683 9919 3689
rect 9968 3692 10732 3720
rect 5169 3655 5227 3661
rect 5169 3652 5181 3655
rect 5000 3624 5181 3652
rect 5169 3621 5181 3624
rect 5215 3621 5227 3655
rect 6638 3652 6644 3664
rect 5169 3615 5227 3621
rect 5644 3624 6644 3652
rect 1653 3587 1711 3593
rect 1653 3584 1665 3587
rect 440 3556 1665 3584
rect 440 3544 446 3556
rect 1653 3553 1665 3556
rect 1699 3553 1711 3587
rect 1653 3547 1711 3553
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 3602 3544 3608 3596
rect 3660 3584 3666 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3660 3556 4077 3584
rect 3660 3544 3666 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 4522 3544 4528 3596
rect 4580 3584 4586 3596
rect 4580 3556 5028 3584
rect 4580 3544 4586 3556
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3786 3516 3792 3528
rect 3559 3488 3792 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4890 3516 4896 3528
rect 4387 3488 4896 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5000 3516 5028 3556
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5000 3488 5273 3516
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5644 3516 5672 3624
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 9876 3652 9904 3683
rect 8444 3624 9904 3652
rect 8444 3612 8450 3624
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 6069 3587 6127 3593
rect 6069 3584 6081 3587
rect 5776 3556 6081 3584
rect 5776 3544 5782 3556
rect 6069 3553 6081 3556
rect 6115 3553 6127 3587
rect 7834 3584 7840 3596
rect 7795 3556 7840 3584
rect 6069 3547 6127 3553
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9677 3587 9735 3593
rect 8996 3556 9168 3584
rect 8996 3544 9002 3556
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5408 3488 5453 3516
rect 5644 3488 5825 3516
rect 5408 3476 5414 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8478 3516 8484 3528
rect 8159 3488 8484 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9140 3516 9168 3556
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9968 3584 9996 3692
rect 10226 3612 10232 3664
rect 10284 3652 10290 3664
rect 10502 3652 10508 3664
rect 10284 3624 10508 3652
rect 10284 3612 10290 3624
rect 10502 3612 10508 3624
rect 10560 3661 10566 3664
rect 10560 3655 10624 3661
rect 10560 3621 10578 3655
rect 10612 3621 10624 3655
rect 10704 3652 10732 3692
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13320 3692 13645 3720
rect 13320 3680 13326 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 14001 3723 14059 3729
rect 14001 3720 14013 3723
rect 13780 3692 14013 3720
rect 13780 3680 13786 3692
rect 14001 3689 14013 3692
rect 14047 3720 14059 3723
rect 16114 3720 16120 3732
rect 14047 3692 16120 3720
rect 14047 3689 14059 3692
rect 14001 3683 14059 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16264 3692 17080 3720
rect 16264 3680 16270 3692
rect 11514 3652 11520 3664
rect 10704 3624 11520 3652
rect 10560 3615 10624 3621
rect 10560 3612 10566 3615
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 16666 3652 16672 3664
rect 11624 3624 16672 3652
rect 10318 3584 10324 3596
rect 9723 3556 9996 3584
rect 10279 3556 10324 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11330 3584 11336 3596
rect 10428 3556 11336 3584
rect 10428 3516 10456 3556
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 9140 3488 10456 3516
rect 9033 3479 9091 3485
rect 2332 3420 5856 3448
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 2332 3380 2360 3420
rect 1820 3352 2360 3380
rect 1820 3340 1826 3352
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3602 3380 3608 3392
rect 2832 3352 3608 3380
rect 2832 3340 2838 3352
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 4764 3352 4813 3380
rect 4764 3340 4770 3352
rect 4801 3349 4813 3352
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 5721 3383 5779 3389
rect 5721 3380 5733 3383
rect 5224 3352 5733 3380
rect 5224 3340 5230 3352
rect 5721 3349 5733 3352
rect 5767 3349 5779 3383
rect 5828 3380 5856 3420
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 9048 3448 9076 3479
rect 8260 3420 9076 3448
rect 8260 3408 8266 3420
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 11624 3448 11652 3624
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 12233 3587 12291 3593
rect 12233 3584 12245 3587
rect 9456 3420 10364 3448
rect 9456 3408 9462 3420
rect 10226 3380 10232 3392
rect 5828 3352 10232 3380
rect 5721 3343 5779 3349
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10336 3380 10364 3420
rect 11256 3420 11652 3448
rect 11716 3556 12245 3584
rect 11256 3380 11284 3420
rect 10336 3352 11284 3380
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 11716 3389 11744 3556
rect 12233 3553 12245 3556
rect 12279 3553 12291 3587
rect 12233 3547 12291 3553
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 13630 3584 13636 3596
rect 12768 3556 13636 3584
rect 12768 3544 12774 3556
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14056 3556 14228 3584
rect 14056 3544 14062 3556
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11848 3488 11989 3516
rect 11848 3476 11854 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 11977 3479 12035 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 14200 3525 14228 3556
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 17052 3593 17080 3692
rect 17218 3612 17224 3664
rect 17276 3612 17282 3664
rect 16485 3587 16543 3593
rect 16485 3584 16497 3587
rect 14332 3556 16497 3584
rect 14332 3544 14338 3556
rect 16485 3553 16497 3556
rect 16531 3553 16543 3587
rect 16485 3547 16543 3553
rect 17037 3587 17095 3593
rect 17037 3553 17049 3587
rect 17083 3553 17095 3587
rect 17236 3584 17264 3612
rect 17773 3587 17831 3593
rect 17773 3584 17785 3587
rect 17236 3556 17785 3584
rect 17037 3547 17095 3553
rect 17773 3553 17785 3556
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3485 17279 3519
rect 18046 3516 18052 3528
rect 18007 3488 18052 3516
rect 17221 3479 17279 3485
rect 16574 3408 16580 3460
rect 16632 3448 16638 3460
rect 16669 3451 16727 3457
rect 16669 3448 16681 3451
rect 16632 3420 16681 3448
rect 16632 3408 16638 3420
rect 16669 3417 16681 3420
rect 16715 3417 16727 3451
rect 16669 3411 16727 3417
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 11388 3352 11713 3380
rect 11388 3340 11394 3352
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 13814 3380 13820 3392
rect 13403 3352 13820 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 17236 3380 17264 3479
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 16540 3352 17264 3380
rect 16540 3340 16546 3352
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 3510 3176 3516 3188
rect 1811 3148 3516 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3752 3148 3801 3176
rect 3752 3136 3758 3148
rect 3789 3145 3801 3148
rect 3835 3145 3847 3179
rect 3789 3139 3847 3145
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 8570 3176 8576 3188
rect 5500 3148 8576 3176
rect 5500 3136 5506 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 16206 3176 16212 3188
rect 10284 3148 16212 3176
rect 10284 3136 10290 3148
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18414 3176 18420 3188
rect 18279 3148 18420 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 2314 3068 2320 3120
rect 2372 3108 2378 3120
rect 2593 3111 2651 3117
rect 2372 3080 2544 3108
rect 2372 3068 2378 3080
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1912 3012 2237 3040
rect 1912 3000 1918 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 2225 3003 2283 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2516 3040 2544 3080
rect 2593 3077 2605 3111
rect 2639 3108 2651 3111
rect 2777 3111 2835 3117
rect 2777 3108 2789 3111
rect 2639 3080 2789 3108
rect 2639 3077 2651 3080
rect 2593 3071 2651 3077
rect 2777 3077 2789 3080
rect 2823 3077 2835 3111
rect 5626 3108 5632 3120
rect 2777 3071 2835 3077
rect 4264 3080 5632 3108
rect 3421 3043 3479 3049
rect 2516 3012 3096 3040
rect 3068 2972 3096 3012
rect 3421 3009 3433 3043
rect 3467 3040 3479 3043
rect 3602 3040 3608 3052
rect 3467 3012 3608 3040
rect 3467 3009 3479 3012
rect 3421 3003 3479 3009
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4264 3049 4292 3080
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 8665 3111 8723 3117
rect 8665 3077 8677 3111
rect 8711 3108 8723 3111
rect 10042 3108 10048 3120
rect 8711 3080 10048 3108
rect 8711 3077 8723 3080
rect 8665 3071 8723 3077
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 11330 3108 11336 3120
rect 10244 3080 11336 3108
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 5166 3040 5172 3052
rect 4479 3012 5172 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5350 3040 5356 3052
rect 5311 3012 5356 3040
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 7834 3040 7840 3052
rect 5460 3012 7840 3040
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 3068 2944 3249 2972
rect 3237 2941 3249 2944
rect 3283 2972 3295 2975
rect 5460 2972 5488 3012
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 9180 3012 9229 3040
rect 9180 3000 9186 3012
rect 9217 3009 9229 3012
rect 9263 3040 9275 3043
rect 9306 3040 9312 3052
rect 9263 3012 9312 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 10244 3049 10272 3080
rect 11330 3068 11336 3080
rect 11388 3068 11394 3120
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 14090 3108 14096 3120
rect 11572 3080 14096 3108
rect 11572 3068 11578 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 16298 3108 16304 3120
rect 16259 3080 16304 3108
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 10560 3012 11253 3040
rect 10560 3000 10566 3012
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 11480 3012 13001 3040
rect 11480 3000 11486 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13372 3012 18092 3040
rect 3283 2944 5488 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 5592 2944 6009 2972
rect 5592 2932 5598 2944
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7282 2972 7288 2984
rect 7239 2944 7288 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2972 7987 2975
rect 8018 2972 8024 2984
rect 7975 2944 8024 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 9030 2972 9036 2984
rect 8991 2944 9036 2972
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 11698 2972 11704 2984
rect 9140 2944 11704 2972
rect 2133 2907 2191 2913
rect 2133 2873 2145 2907
rect 2179 2904 2191 2907
rect 2593 2907 2651 2913
rect 2593 2904 2605 2907
rect 2179 2876 2605 2904
rect 2179 2873 2191 2876
rect 2133 2867 2191 2873
rect 2593 2873 2605 2876
rect 2639 2873 2651 2907
rect 2593 2867 2651 2873
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 3145 2907 3203 2913
rect 3145 2904 3157 2907
rect 2924 2876 3157 2904
rect 2924 2864 2930 2876
rect 3145 2873 3157 2876
rect 3191 2873 3203 2907
rect 3145 2867 3203 2873
rect 5169 2907 5227 2913
rect 5169 2873 5181 2907
rect 5215 2904 5227 2907
rect 6178 2904 6184 2916
rect 5215 2876 6184 2904
rect 5215 2873 5227 2876
rect 5169 2867 5227 2873
rect 6178 2864 6184 2876
rect 6236 2864 6242 2916
rect 6273 2907 6331 2913
rect 6273 2873 6285 2907
rect 6319 2904 6331 2907
rect 6730 2904 6736 2916
rect 6319 2876 6736 2904
rect 6319 2873 6331 2876
rect 6273 2867 6331 2873
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 7469 2907 7527 2913
rect 7469 2873 7481 2907
rect 7515 2904 7527 2907
rect 7558 2904 7564 2916
rect 7515 2876 7564 2904
rect 7515 2873 7527 2876
rect 7469 2867 7527 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8205 2907 8263 2913
rect 8205 2873 8217 2907
rect 8251 2904 8263 2907
rect 8478 2904 8484 2916
rect 8251 2876 8484 2904
rect 8251 2873 8263 2876
rect 8205 2867 8263 2873
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 9140 2913 9168 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 13372 2972 13400 3012
rect 12032 2944 13400 2972
rect 12032 2932 12038 2944
rect 13446 2932 13452 2984
rect 13504 2972 13510 2984
rect 14185 2975 14243 2981
rect 13504 2944 13549 2972
rect 13504 2932 13510 2944
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 14642 2972 14648 2984
rect 14231 2944 14648 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2972 14979 2975
rect 15286 2972 15292 2984
rect 14967 2944 15292 2972
rect 14967 2941 14979 2944
rect 14921 2935 14979 2941
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 16298 2932 16304 2984
rect 16356 2972 16362 2984
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 16356 2944 16497 2972
rect 16356 2932 16362 2944
rect 16485 2941 16497 2944
rect 16531 2941 16543 2975
rect 17218 2972 17224 2984
rect 17179 2944 17224 2972
rect 16485 2935 16543 2941
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 18064 2981 18092 3012
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 9125 2907 9183 2913
rect 9125 2904 9137 2907
rect 8588 2876 9137 2904
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 3326 2836 3332 2848
rect 2096 2808 3332 2836
rect 2096 2796 2102 2808
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 4154 2836 4160 2848
rect 4115 2808 4160 2836
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4798 2836 4804 2848
rect 4759 2808 4804 2836
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5258 2836 5264 2848
rect 5219 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 5810 2836 5816 2848
rect 5684 2808 5816 2836
rect 5684 2796 5690 2808
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 8588 2836 8616 2876
rect 9125 2873 9137 2876
rect 9171 2873 9183 2907
rect 9125 2867 9183 2873
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2904 10103 2907
rect 11149 2907 11207 2913
rect 10091 2876 10732 2904
rect 10091 2873 10103 2876
rect 10045 2867 10103 2873
rect 6052 2808 8616 2836
rect 6052 2796 6058 2808
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10192 2808 10237 2836
rect 10192 2796 10198 2808
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10502 2836 10508 2848
rect 10376 2808 10508 2836
rect 10376 2796 10382 2808
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 10704 2845 10732 2876
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 12805 2907 12863 2913
rect 11195 2876 12480 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 10689 2839 10747 2845
rect 10689 2805 10701 2839
rect 10735 2805 10747 2839
rect 11054 2836 11060 2848
rect 11015 2808 11060 2836
rect 10689 2799 10747 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11882 2836 11888 2848
rect 11843 2808 11888 2836
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12452 2845 12480 2876
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 12851 2876 13124 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2805 12495 2839
rect 12437 2799 12495 2805
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12768 2808 12909 2836
rect 12768 2796 12774 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 13096 2836 13124 2876
rect 13170 2864 13176 2916
rect 13228 2904 13234 2916
rect 13725 2907 13783 2913
rect 13725 2904 13737 2907
rect 13228 2876 13737 2904
rect 13228 2864 13234 2876
rect 13725 2873 13737 2876
rect 13771 2873 13783 2907
rect 13725 2867 13783 2873
rect 14461 2907 14519 2913
rect 14461 2873 14473 2907
rect 14507 2904 14519 2907
rect 14826 2904 14832 2916
rect 14507 2876 14832 2904
rect 14507 2873 14519 2876
rect 14461 2867 14519 2873
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 15197 2907 15255 2913
rect 15197 2873 15209 2907
rect 15243 2904 15255 2907
rect 15654 2904 15660 2916
rect 15243 2876 15660 2904
rect 15243 2873 15255 2876
rect 15197 2867 15255 2873
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 16758 2904 16764 2916
rect 16719 2876 16764 2904
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 17497 2907 17555 2913
rect 17497 2873 17509 2907
rect 17543 2904 17555 2907
rect 19426 2904 19432 2916
rect 17543 2876 19432 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 13538 2836 13544 2848
rect 13096 2808 13544 2836
rect 12897 2799 12955 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2038 2632 2044 2644
rect 1995 2604 2044 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2961 2635 3019 2641
rect 2961 2632 2973 2635
rect 2455 2604 2973 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2961 2601 2973 2604
rect 3007 2601 3019 2635
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 2961 2595 3019 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4341 2635 4399 2641
rect 4341 2632 4353 2635
rect 4212 2604 4353 2632
rect 4212 2592 4218 2604
rect 4341 2601 4353 2604
rect 4387 2601 4399 2635
rect 4341 2595 4399 2601
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 4798 2632 4804 2644
rect 4755 2604 4804 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5132 2604 5365 2632
rect 5132 2592 5138 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5684 2604 5733 2632
rect 5684 2592 5690 2604
rect 5721 2601 5733 2604
rect 5767 2601 5779 2635
rect 5721 2595 5779 2601
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 6236 2604 6377 2632
rect 6236 2592 6242 2604
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 8711 2604 8984 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 5442 2564 5448 2576
rect 2363 2536 5448 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 7834 2564 7840 2576
rect 5859 2536 7840 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8956 2564 8984 2604
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9766 2632 9772 2644
rect 9088 2604 9772 2632
rect 9088 2592 9094 2604
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 10100 2604 10149 2632
rect 10100 2592 10106 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 11054 2632 11060 2644
rect 10827 2604 11060 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11241 2635 11299 2641
rect 11241 2632 11253 2635
rect 11204 2604 11253 2632
rect 11204 2592 11210 2604
rect 11241 2601 11253 2604
rect 11287 2601 11299 2635
rect 12434 2632 12440 2644
rect 11241 2595 11299 2601
rect 11532 2604 12440 2632
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 8956 2536 10241 2564
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 2832 2468 3433 2496
rect 2832 2456 2838 2468
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 3602 2456 3608 2508
rect 3660 2496 3666 2508
rect 4430 2496 4436 2508
rect 3660 2468 4436 2496
rect 3660 2456 3666 2468
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4764 2468 4813 2496
rect 4764 2456 4770 2468
rect 4801 2465 4813 2468
rect 4847 2465 4859 2499
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 4801 2459 4859 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2496 7987 2499
rect 8846 2496 8852 2508
rect 7975 2468 8852 2496
rect 7975 2465 7987 2468
rect 7929 2459 7987 2465
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 9030 2496 9036 2508
rect 8991 2468 9036 2496
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 10870 2496 10876 2508
rect 9324 2468 10876 2496
rect 9324 2440 9352 2468
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 11532 2496 11560 2604
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 16669 2635 16727 2641
rect 16669 2601 16681 2635
rect 16715 2632 16727 2635
rect 16850 2632 16856 2644
rect 16715 2604 16856 2632
rect 16715 2601 16727 2604
rect 16669 2595 16727 2601
rect 11195 2468 11560 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11664 2468 11805 2496
rect 11664 2456 11670 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12400 2468 12633 2496
rect 12400 2456 12406 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 14458 2496 14464 2508
rect 14415 2468 14464 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 16776 2505 16804 2604
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2465 16819 2499
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 16761 2459 16819 2465
rect 17328 2468 17509 2496
rect 2406 2388 2412 2440
rect 2464 2428 2470 2440
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2464 2400 2605 2428
rect 2464 2388 2470 2400
rect 2593 2397 2605 2400
rect 2639 2428 2651 2431
rect 3510 2428 3516 2440
rect 2639 2400 3188 2428
rect 3471 2400 3516 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 3160 2360 3188 2400
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5718 2428 5724 2440
rect 5031 2400 5724 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 5920 2360 5948 2391
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6144 2400 7113 2428
rect 6144 2388 6150 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 3160 2332 5948 2360
rect 8220 2360 8248 2391
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8812 2400 9137 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 9125 2391 9183 2397
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10888 2428 10916 2456
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 10888 2400 11345 2428
rect 11333 2397 11345 2400
rect 11379 2428 11391 2431
rect 11422 2428 11428 2440
rect 11379 2400 11428 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 9398 2360 9404 2372
rect 8220 2332 9404 2360
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 10134 2360 10140 2372
rect 9815 2332 10140 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 10134 2320 10140 2332
rect 10192 2320 10198 2372
rect 11238 2320 11244 2372
rect 11296 2360 11302 2372
rect 11992 2360 12020 2391
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12216 2400 12817 2428
rect 12216 2388 12222 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 13964 2400 14565 2428
rect 13964 2388 13970 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 17034 2428 17040 2440
rect 16995 2400 17040 2428
rect 14553 2391 14611 2397
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 11296 2332 12020 2360
rect 11296 2320 11302 2332
rect 16482 2320 16488 2372
rect 16540 2360 16546 2372
rect 17328 2369 17356 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 17770 2428 17776 2440
rect 17731 2400 17776 2428
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 17313 2363 17371 2369
rect 17313 2360 17325 2363
rect 16540 2332 17325 2360
rect 16540 2320 16546 2332
rect 17313 2329 17325 2332
rect 17359 2329 17371 2363
rect 17313 2323 17371 2329
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 3694 2048 3700 2100
rect 3752 2088 3758 2100
rect 8386 2088 8392 2100
rect 3752 2060 8392 2088
rect 3752 2048 3758 2060
rect 8386 2048 8392 2060
rect 8444 2048 8450 2100
rect 1946 1980 1952 2032
rect 2004 2020 2010 2032
rect 6914 2020 6920 2032
rect 2004 1992 6920 2020
rect 2004 1980 2010 1992
rect 6914 1980 6920 1992
rect 6972 1980 6978 2032
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 8662 1340 8668 1352
rect 3384 1312 8668 1340
rect 3384 1300 3390 1312
rect 8662 1300 8668 1312
rect 8720 1300 8726 1352
rect 4062 1164 4068 1216
rect 4120 1204 4126 1216
rect 11882 1204 11888 1216
rect 4120 1176 11888 1204
rect 4120 1164 4126 1176
rect 11882 1164 11888 1176
rect 11940 1164 11946 1216
rect 3694 1028 3700 1080
rect 3752 1068 3758 1080
rect 9214 1068 9220 1080
rect 3752 1040 9220 1068
rect 3752 1028 3758 1040
rect 9214 1028 9220 1040
rect 9272 1028 9278 1080
<< via1 >>
rect 3332 16532 3384 16584
rect 6460 16532 6512 16584
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 3424 14603 3476 14612
rect 3424 14569 3433 14603
rect 3433 14569 3467 14603
rect 3467 14569 3476 14603
rect 3424 14560 3476 14569
rect 4988 14560 5040 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 2044 14535 2096 14544
rect 2044 14501 2053 14535
rect 2053 14501 2087 14535
rect 2087 14501 2096 14535
rect 2044 14492 2096 14501
rect 2780 14535 2832 14544
rect 2780 14501 2789 14535
rect 2789 14501 2823 14535
rect 2823 14501 2832 14535
rect 2780 14492 2832 14501
rect 3332 14424 3384 14476
rect 5172 14424 5224 14476
rect 8024 14424 8076 14476
rect 3608 14356 3660 14408
rect 4068 14288 4120 14340
rect 17592 14288 17644 14340
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 1676 14016 1728 14068
rect 17592 14059 17644 14068
rect 3240 13991 3292 14000
rect 3240 13957 3249 13991
rect 3249 13957 3283 13991
rect 3283 13957 3292 13991
rect 3240 13948 3292 13957
rect 3792 13991 3844 14000
rect 3792 13957 3801 13991
rect 3801 13957 3835 13991
rect 3835 13957 3844 13991
rect 3792 13948 3844 13957
rect 5632 13948 5684 14000
rect 2780 13880 2832 13932
rect 5448 13880 5500 13932
rect 6276 13880 6328 13932
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 14924 13880 14976 13932
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 18236 14059 18288 14068
rect 18236 14025 18245 14059
rect 18245 14025 18279 14059
rect 18279 14025 18288 14059
rect 18236 14016 18288 14025
rect 16764 13948 16816 14000
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3608 13855 3660 13864
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 3608 13812 3660 13821
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 11612 13812 11664 13864
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 17868 13812 17920 13864
rect 1768 13744 1820 13796
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 7380 13744 7432 13796
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 2872 13472 2924 13524
rect 6000 13472 6052 13524
rect 7288 13472 7340 13524
rect 7472 13472 7524 13524
rect 11888 13472 11940 13524
rect 9772 13404 9824 13456
rect 15200 13404 15252 13456
rect 1768 13336 1820 13388
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 3332 13336 3384 13388
rect 5264 13336 5316 13388
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 1400 13268 1452 13320
rect 5908 13311 5960 13320
rect 2504 13200 2556 13252
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 6092 13311 6144 13320
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6092 13268 6144 13277
rect 6276 13268 6328 13320
rect 2044 13132 2096 13184
rect 3792 13132 3844 13184
rect 11152 13336 11204 13388
rect 6552 13268 6604 13320
rect 7104 13311 7156 13320
rect 7104 13277 7113 13311
rect 7113 13277 7147 13311
rect 7147 13277 7156 13311
rect 7104 13268 7156 13277
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 7748 13200 7800 13252
rect 14648 13336 14700 13388
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 11796 13200 11848 13252
rect 15292 13200 15344 13252
rect 7564 13132 7616 13184
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 10968 13175 11020 13184
rect 10968 13141 10977 13175
rect 10977 13141 11011 13175
rect 11011 13141 11020 13175
rect 10968 13132 11020 13141
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 2964 12928 3016 12980
rect 4712 12928 4764 12980
rect 5816 12928 5868 12980
rect 5540 12860 5592 12912
rect 6000 12860 6052 12912
rect 2688 12792 2740 12844
rect 3056 12792 3108 12844
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 2412 12724 2464 12776
rect 1492 12656 1544 12708
rect 1860 12588 1912 12640
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 4620 12792 4672 12844
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 7472 12928 7524 12980
rect 12808 12928 12860 12980
rect 16488 12928 16540 12980
rect 4344 12724 4396 12776
rect 4528 12656 4580 12708
rect 7104 12792 7156 12844
rect 7472 12792 7524 12844
rect 9312 12792 9364 12844
rect 7932 12724 7984 12776
rect 2136 12588 2188 12597
rect 3148 12631 3200 12640
rect 3148 12597 3157 12631
rect 3157 12597 3191 12631
rect 3191 12597 3200 12631
rect 3148 12588 3200 12597
rect 7380 12656 7432 12708
rect 5724 12588 5776 12640
rect 5816 12588 5868 12640
rect 6736 12588 6788 12640
rect 7748 12588 7800 12640
rect 8024 12656 8076 12708
rect 10692 12860 10744 12912
rect 11796 12860 11848 12912
rect 11888 12860 11940 12912
rect 10876 12792 10928 12844
rect 11612 12792 11664 12844
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12348 12724 12400 12776
rect 12808 12699 12860 12708
rect 12808 12665 12817 12699
rect 12817 12665 12851 12699
rect 12851 12665 12860 12699
rect 12808 12656 12860 12665
rect 17040 12656 17092 12708
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8668 12588 8720 12640
rect 9220 12588 9272 12640
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 13544 12631 13596 12640
rect 13544 12597 13553 12631
rect 13553 12597 13587 12631
rect 13587 12597 13596 12631
rect 13544 12588 13596 12597
rect 15016 12588 15068 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 2136 12384 2188 12436
rect 3148 12384 3200 12436
rect 4528 12384 4580 12436
rect 4896 12384 4948 12436
rect 5724 12384 5776 12436
rect 9680 12384 9732 12436
rect 14740 12384 14792 12436
rect 15200 12384 15252 12436
rect 3424 12316 3476 12368
rect 11520 12316 11572 12368
rect 2044 12248 2096 12300
rect 3332 12291 3384 12300
rect 3332 12257 3341 12291
rect 3341 12257 3375 12291
rect 3375 12257 3384 12291
rect 3332 12248 3384 12257
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 6644 12248 6696 12300
rect 7656 12248 7708 12300
rect 10508 12248 10560 12300
rect 11612 12248 11664 12300
rect 14280 12248 14332 12300
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 2780 12180 2832 12232
rect 4528 12223 4580 12232
rect 2228 12112 2280 12164
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 3792 12112 3844 12164
rect 6368 12180 6420 12232
rect 7288 12112 7340 12164
rect 8944 12180 8996 12232
rect 9312 12180 9364 12232
rect 9404 12180 9456 12232
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 8760 12112 8812 12164
rect 3608 12044 3660 12096
rect 6460 12044 6512 12096
rect 8116 12044 8168 12096
rect 10324 12044 10376 12096
rect 10784 12112 10836 12164
rect 12716 12180 12768 12232
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 17776 12223 17828 12232
rect 13820 12180 13872 12189
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 11428 12044 11480 12096
rect 11888 12044 11940 12096
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 15568 12112 15620 12164
rect 15108 12044 15160 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2688 11840 2740 11892
rect 3700 11840 3752 11892
rect 5908 11772 5960 11824
rect 9680 11772 9732 11824
rect 11612 11840 11664 11892
rect 16120 11840 16172 11892
rect 5540 11704 5592 11756
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 8576 11704 8628 11756
rect 9128 11704 9180 11756
rect 13176 11772 13228 11824
rect 1584 11636 1636 11688
rect 2504 11636 2556 11688
rect 2964 11500 3016 11552
rect 4252 11636 4304 11688
rect 4804 11636 4856 11688
rect 4344 11568 4396 11620
rect 6276 11636 6328 11688
rect 16580 11704 16632 11756
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 5816 11500 5868 11552
rect 8760 11636 8812 11688
rect 9404 11636 9456 11688
rect 10324 11636 10376 11688
rect 11060 11636 11112 11688
rect 11704 11636 11756 11688
rect 13268 11679 13320 11688
rect 13268 11645 13277 11679
rect 13277 11645 13311 11679
rect 13311 11645 13320 11679
rect 13268 11636 13320 11645
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 14004 11636 14056 11688
rect 15108 11636 15160 11688
rect 17132 11636 17184 11688
rect 17960 11636 18012 11688
rect 7656 11568 7708 11620
rect 8024 11568 8076 11620
rect 10600 11568 10652 11620
rect 7840 11500 7892 11552
rect 8300 11500 8352 11552
rect 8852 11500 8904 11552
rect 9496 11543 9548 11552
rect 9496 11509 9505 11543
rect 9505 11509 9539 11543
rect 9539 11509 9548 11543
rect 9496 11500 9548 11509
rect 9864 11500 9916 11552
rect 10968 11500 11020 11552
rect 14372 11568 14424 11620
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 14832 11500 14884 11552
rect 15016 11500 15068 11552
rect 15108 11500 15160 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 16672 11500 16724 11552
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 17500 11500 17552 11552
rect 18420 11500 18472 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2504 11296 2556 11348
rect 1952 11160 2004 11212
rect 4344 11228 4396 11280
rect 4160 11160 4212 11212
rect 5540 11228 5592 11280
rect 5908 11228 5960 11280
rect 6092 11228 6144 11280
rect 8208 11296 8260 11348
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 9128 11296 9180 11348
rect 14280 11339 14332 11348
rect 5724 11160 5776 11212
rect 4160 11024 4212 11076
rect 6092 11092 6144 11144
rect 4988 11024 5040 11076
rect 7656 11228 7708 11280
rect 7748 11228 7800 11280
rect 11520 11228 11572 11280
rect 11704 11271 11756 11280
rect 11704 11237 11713 11271
rect 11713 11237 11747 11271
rect 11747 11237 11756 11271
rect 11704 11228 11756 11237
rect 10968 11160 11020 11212
rect 7840 11092 7892 11144
rect 8576 11092 8628 11144
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 13820 11228 13872 11280
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 15016 11228 15068 11280
rect 17224 11271 17276 11280
rect 17224 11237 17258 11271
rect 17258 11237 17276 11271
rect 17224 11228 17276 11237
rect 13912 11160 13964 11212
rect 14096 11160 14148 11212
rect 15108 11160 15160 11212
rect 9036 11024 9088 11076
rect 12532 11024 12584 11076
rect 1584 10956 1636 11008
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 3424 10956 3476 11008
rect 4804 10956 4856 11008
rect 9588 10956 9640 11008
rect 10600 10956 10652 11008
rect 12624 10956 12676 11008
rect 14004 10999 14056 11008
rect 14004 10965 14013 10999
rect 14013 10965 14047 10999
rect 14047 10965 14056 10999
rect 14004 10956 14056 10965
rect 15292 10956 15344 11008
rect 16304 10956 16356 11008
rect 17592 10956 17644 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 1400 10795 1452 10804
rect 1400 10761 1409 10795
rect 1409 10761 1443 10795
rect 1443 10761 1452 10795
rect 1400 10752 1452 10761
rect 4252 10752 4304 10804
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 7748 10752 7800 10804
rect 8484 10752 8536 10804
rect 9128 10684 9180 10736
rect 10876 10752 10928 10804
rect 11796 10752 11848 10804
rect 13360 10752 13412 10804
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 2136 10616 2188 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 9496 10616 9548 10668
rect 12808 10684 12860 10736
rect 16120 10684 16172 10736
rect 11060 10616 11112 10668
rect 11428 10616 11480 10668
rect 12348 10616 12400 10668
rect 13820 10616 13872 10668
rect 14004 10616 14056 10668
rect 1584 10548 1636 10600
rect 2688 10591 2740 10600
rect 2688 10557 2722 10591
rect 2722 10557 2740 10591
rect 2688 10548 2740 10557
rect 4160 10548 4212 10600
rect 5908 10548 5960 10600
rect 7472 10548 7524 10600
rect 9036 10548 9088 10600
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 12532 10548 12584 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 3148 10480 3200 10532
rect 7656 10480 7708 10532
rect 3332 10412 3384 10464
rect 3700 10412 3752 10464
rect 4068 10412 4120 10464
rect 10508 10480 10560 10532
rect 10600 10480 10652 10532
rect 12808 10523 12860 10532
rect 12808 10489 12817 10523
rect 12817 10489 12851 10523
rect 12851 10489 12860 10523
rect 12808 10480 12860 10489
rect 13176 10480 13228 10532
rect 14648 10480 14700 10532
rect 15568 10616 15620 10668
rect 15752 10616 15804 10668
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 16580 10523 16632 10532
rect 16580 10489 16614 10523
rect 16614 10489 16632 10523
rect 16580 10480 16632 10489
rect 17592 10480 17644 10532
rect 8024 10412 8076 10464
rect 9404 10412 9456 10464
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 11612 10412 11664 10464
rect 13452 10412 13504 10464
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18328 10412 18380 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2412 10208 2464 10260
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3424 10140 3476 10192
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 2320 10072 2372 10124
rect 5356 10208 5408 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6000 10208 6052 10260
rect 6460 10208 6512 10260
rect 8392 10208 8444 10260
rect 10876 10208 10928 10260
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 12348 10208 12400 10260
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 13544 10208 13596 10260
rect 13728 10208 13780 10260
rect 16120 10208 16172 10260
rect 5448 10140 5500 10192
rect 7288 10140 7340 10192
rect 9404 10140 9456 10192
rect 6736 10072 6788 10124
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 4160 10047 4212 10056
rect 1584 9868 1636 9920
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 5172 10004 5224 10056
rect 5448 10004 5500 10056
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 5356 9936 5408 9988
rect 5724 9936 5776 9988
rect 3700 9868 3752 9920
rect 7104 10004 7156 10056
rect 8208 10072 8260 10124
rect 14096 10140 14148 10192
rect 14372 10183 14424 10192
rect 14372 10149 14381 10183
rect 14381 10149 14415 10183
rect 14415 10149 14424 10183
rect 14372 10140 14424 10149
rect 17868 10208 17920 10260
rect 7472 10004 7524 10056
rect 10508 10072 10560 10124
rect 11152 10072 11204 10124
rect 11980 10072 12032 10124
rect 12072 10072 12124 10124
rect 14556 10072 14608 10124
rect 6460 9936 6512 9988
rect 7564 9868 7616 9920
rect 8852 9868 8904 9920
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 13820 10004 13872 10056
rect 15108 10004 15160 10056
rect 16120 10004 16172 10056
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 10968 9868 11020 9920
rect 11060 9868 11112 9920
rect 13636 9936 13688 9988
rect 14924 9936 14976 9988
rect 15660 9936 15712 9988
rect 17684 10004 17736 10056
rect 18052 9979 18104 9988
rect 18052 9945 18061 9979
rect 18061 9945 18095 9979
rect 18095 9945 18104 9979
rect 18052 9936 18104 9945
rect 13452 9868 13504 9920
rect 14464 9868 14516 9920
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 17684 9868 17736 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3148 9664 3200 9716
rect 5080 9664 5132 9716
rect 5264 9664 5316 9716
rect 2044 9639 2096 9648
rect 2044 9605 2053 9639
rect 2053 9605 2087 9639
rect 2087 9605 2096 9639
rect 2044 9596 2096 9605
rect 4436 9596 4488 9648
rect 6368 9664 6420 9716
rect 14556 9664 14608 9716
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 11060 9596 11112 9648
rect 12072 9596 12124 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14096 9639 14148 9648
rect 14096 9605 14105 9639
rect 14105 9605 14139 9639
rect 14139 9605 14148 9639
rect 14096 9596 14148 9605
rect 2136 9528 2188 9580
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 4252 9528 4304 9580
rect 4344 9528 4396 9580
rect 4160 9460 4212 9512
rect 6736 9528 6788 9580
rect 3976 9392 4028 9444
rect 4712 9392 4764 9444
rect 9128 9503 9180 9512
rect 9128 9469 9162 9503
rect 9162 9469 9180 9503
rect 9128 9460 9180 9469
rect 9404 9460 9456 9512
rect 11336 9528 11388 9580
rect 12348 9528 12400 9580
rect 15292 9664 15344 9716
rect 16120 9664 16172 9716
rect 16580 9664 16632 9716
rect 17224 9664 17276 9716
rect 16028 9596 16080 9648
rect 16212 9596 16264 9648
rect 5172 9392 5224 9444
rect 5540 9392 5592 9444
rect 6368 9392 6420 9444
rect 7196 9392 7248 9444
rect 7380 9392 7432 9444
rect 1400 9324 1452 9376
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 3424 9367 3476 9376
rect 2504 9324 2556 9333
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 4344 9324 4396 9376
rect 4988 9324 5040 9376
rect 7472 9324 7524 9376
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 8576 9392 8628 9444
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11980 9460 12032 9512
rect 16396 9528 16448 9580
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 10968 9392 11020 9444
rect 13912 9460 13964 9512
rect 13268 9392 13320 9444
rect 15660 9460 15712 9512
rect 17776 9460 17828 9512
rect 11152 9324 11204 9376
rect 11428 9324 11480 9376
rect 11612 9324 11664 9376
rect 14832 9392 14884 9444
rect 15016 9392 15068 9444
rect 15292 9324 15344 9376
rect 17776 9324 17828 9376
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2596 9120 2648 9172
rect 3516 9120 3568 9172
rect 5264 9120 5316 9172
rect 5816 9120 5868 9172
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 6736 9120 6788 9172
rect 7564 9163 7616 9172
rect 7564 9129 7573 9163
rect 7573 9129 7607 9163
rect 7607 9129 7616 9163
rect 7564 9120 7616 9129
rect 7656 9120 7708 9172
rect 9220 9120 9272 9172
rect 10692 9120 10744 9172
rect 12348 9120 12400 9172
rect 14372 9120 14424 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 15200 9120 15252 9172
rect 17316 9120 17368 9172
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 2688 8984 2740 9036
rect 4712 9052 4764 9104
rect 6368 9052 6420 9104
rect 7840 9052 7892 9104
rect 8760 9052 8812 9104
rect 9036 9052 9088 9104
rect 7472 9027 7524 9036
rect 2412 8916 2464 8968
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 7380 8916 7432 8968
rect 8852 8984 8904 9036
rect 9680 9052 9732 9104
rect 13544 9095 13596 9104
rect 13544 9061 13553 9095
rect 13553 9061 13587 9095
rect 13587 9061 13596 9095
rect 13544 9052 13596 9061
rect 17684 9052 17736 9104
rect 3424 8848 3476 8900
rect 9128 8916 9180 8968
rect 10232 8984 10284 9036
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 11428 8984 11480 9036
rect 11612 9027 11664 9036
rect 11612 8993 11646 9027
rect 11646 8993 11664 9027
rect 11612 8984 11664 8993
rect 15384 8984 15436 9036
rect 16028 9027 16080 9036
rect 16028 8993 16062 9027
rect 16062 8993 16080 9027
rect 16028 8984 16080 8993
rect 10416 8916 10468 8968
rect 10876 8959 10928 8968
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 10968 8916 11020 8968
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 13820 8959 13872 8968
rect 13820 8925 13829 8959
rect 13829 8925 13863 8959
rect 13863 8925 13872 8959
rect 13820 8916 13872 8925
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 14924 8916 14976 8968
rect 17592 8916 17644 8968
rect 1584 8780 1636 8832
rect 3148 8780 3200 8832
rect 4804 8780 4856 8832
rect 4988 8780 5040 8832
rect 6368 8780 6420 8832
rect 6552 8780 6604 8832
rect 7288 8780 7340 8832
rect 8392 8780 8444 8832
rect 9312 8780 9364 8832
rect 10324 8780 10376 8832
rect 10876 8780 10928 8832
rect 13544 8780 13596 8832
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 14280 8780 14332 8832
rect 15384 8780 15436 8832
rect 16948 8780 17000 8832
rect 17132 8823 17184 8832
rect 17132 8789 17141 8823
rect 17141 8789 17175 8823
rect 17175 8789 17184 8823
rect 17132 8780 17184 8789
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2504 8576 2556 8628
rect 3792 8576 3844 8628
rect 4344 8576 4396 8628
rect 3700 8440 3752 8492
rect 7472 8576 7524 8628
rect 7932 8619 7984 8628
rect 7932 8585 7941 8619
rect 7941 8585 7975 8619
rect 7975 8585 7984 8619
rect 7932 8576 7984 8585
rect 5908 8508 5960 8560
rect 6368 8508 6420 8560
rect 8944 8508 8996 8560
rect 1584 8372 1636 8424
rect 1676 8304 1728 8356
rect 2596 8372 2648 8424
rect 8208 8440 8260 8492
rect 8484 8440 8536 8492
rect 5724 8372 5776 8424
rect 4252 8304 4304 8356
rect 4436 8347 4488 8356
rect 4436 8313 4470 8347
rect 4470 8313 4488 8347
rect 4436 8304 4488 8313
rect 5356 8304 5408 8356
rect 7748 8372 7800 8424
rect 7932 8372 7984 8424
rect 10048 8372 10100 8424
rect 10968 8576 11020 8628
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 15568 8576 15620 8628
rect 10324 8551 10376 8560
rect 10324 8517 10333 8551
rect 10333 8517 10367 8551
rect 10367 8517 10376 8551
rect 10324 8508 10376 8517
rect 13820 8508 13872 8560
rect 10232 8440 10284 8492
rect 13544 8440 13596 8492
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 15384 8440 15436 8492
rect 11704 8372 11756 8424
rect 14004 8372 14056 8424
rect 14280 8372 14332 8424
rect 4068 8236 4120 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 6092 8236 6144 8288
rect 8484 8236 8536 8288
rect 9404 8236 9456 8288
rect 9588 8304 9640 8356
rect 10876 8347 10928 8356
rect 10876 8313 10910 8347
rect 10910 8313 10928 8347
rect 10876 8304 10928 8313
rect 11060 8304 11112 8356
rect 12164 8304 12216 8356
rect 16212 8372 16264 8424
rect 16396 8372 16448 8424
rect 17500 8372 17552 8424
rect 10232 8236 10284 8288
rect 13728 8236 13780 8288
rect 14832 8304 14884 8356
rect 15200 8236 15252 8288
rect 15660 8236 15712 8288
rect 17224 8304 17276 8356
rect 17684 8279 17736 8288
rect 17684 8245 17693 8279
rect 17693 8245 17727 8279
rect 17727 8245 17736 8279
rect 17684 8236 17736 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 2688 8032 2740 8084
rect 4528 8032 4580 8084
rect 5724 8032 5776 8084
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 8944 8032 8996 8084
rect 10416 8032 10468 8084
rect 11428 8032 11480 8084
rect 12440 8032 12492 8084
rect 3792 7964 3844 8016
rect 6000 7964 6052 8016
rect 6644 7964 6696 8016
rect 11244 7964 11296 8016
rect 13360 8032 13412 8084
rect 14188 8032 14240 8084
rect 15568 7964 15620 8016
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4252 7896 4304 7948
rect 6552 7896 6604 7948
rect 7748 7896 7800 7948
rect 7932 7939 7984 7948
rect 7932 7905 7941 7939
rect 7941 7905 7975 7939
rect 7975 7905 7984 7939
rect 7932 7896 7984 7905
rect 4528 7828 4580 7880
rect 4712 7828 4764 7880
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 4988 7760 5040 7812
rect 7196 7828 7248 7880
rect 6828 7760 6880 7812
rect 9588 7828 9640 7880
rect 10784 7896 10836 7948
rect 10968 7828 11020 7880
rect 10600 7760 10652 7812
rect 11060 7760 11112 7812
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 4344 7692 4396 7744
rect 6000 7692 6052 7744
rect 7472 7692 7524 7744
rect 8484 7692 8536 7744
rect 9036 7692 9088 7744
rect 9588 7692 9640 7744
rect 13176 7896 13228 7948
rect 16672 7896 16724 7948
rect 12256 7828 12308 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15200 7828 15252 7880
rect 16304 7828 16356 7880
rect 13820 7760 13872 7812
rect 15016 7760 15068 7812
rect 13912 7692 13964 7744
rect 15108 7692 15160 7744
rect 15568 7760 15620 7812
rect 16212 7760 16264 7812
rect 16948 7964 17000 8016
rect 17316 7896 17368 7948
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 17224 7828 17276 7880
rect 16856 7760 16908 7812
rect 17684 7828 17736 7880
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 1952 7488 2004 7540
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 4252 7488 4304 7540
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 2872 7420 2924 7472
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 2596 7352 2648 7404
rect 4344 7420 4396 7472
rect 1860 7284 1912 7336
rect 2228 7284 2280 7336
rect 4436 7352 4488 7404
rect 6000 7420 6052 7472
rect 4896 7284 4948 7336
rect 10692 7488 10744 7540
rect 10784 7488 10836 7540
rect 11980 7488 12032 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 14004 7488 14056 7540
rect 6828 7420 6880 7472
rect 6552 7352 6604 7404
rect 12256 7420 12308 7472
rect 6736 7284 6788 7336
rect 10232 7352 10284 7404
rect 11612 7352 11664 7404
rect 11704 7352 11756 7404
rect 15016 7420 15068 7472
rect 15108 7352 15160 7404
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 8576 7284 8628 7336
rect 10784 7284 10836 7336
rect 2320 7216 2372 7268
rect 2228 7148 2280 7200
rect 2412 7148 2464 7200
rect 3332 7148 3384 7200
rect 4436 7148 4488 7200
rect 8116 7216 8168 7268
rect 8392 7216 8444 7268
rect 11612 7216 11664 7268
rect 12072 7216 12124 7268
rect 12716 7216 12768 7268
rect 6000 7148 6052 7200
rect 6644 7148 6696 7200
rect 8300 7148 8352 7200
rect 9496 7148 9548 7200
rect 9772 7148 9824 7200
rect 11060 7148 11112 7200
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 11888 7148 11940 7200
rect 12532 7148 12584 7200
rect 12624 7148 12676 7200
rect 13360 7148 13412 7200
rect 13544 7284 13596 7336
rect 15568 7352 15620 7404
rect 17224 7352 17276 7404
rect 16672 7284 16724 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 15200 7216 15252 7268
rect 16580 7216 16632 7268
rect 14924 7148 14976 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15292 7191 15344 7200
rect 15016 7148 15068 7157
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15292 7148 15344 7157
rect 15568 7148 15620 7200
rect 16488 7148 16540 7200
rect 17592 7148 17644 7200
rect 17868 7148 17920 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 4620 6944 4672 6996
rect 5080 6944 5132 6996
rect 6552 6944 6604 6996
rect 1308 6876 1360 6928
rect 7748 6944 7800 6996
rect 8852 6944 8904 6996
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 1860 6808 1912 6860
rect 2504 6851 2556 6860
rect 2504 6817 2538 6851
rect 2538 6817 2556 6851
rect 2504 6808 2556 6817
rect 3056 6808 3108 6860
rect 4620 6851 4672 6860
rect 1584 6740 1636 6792
rect 4620 6817 4629 6851
rect 4629 6817 4663 6851
rect 4663 6817 4672 6851
rect 4620 6808 4672 6817
rect 5172 6808 5224 6860
rect 6092 6808 6144 6860
rect 6920 6851 6972 6860
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 9588 6876 9640 6928
rect 11060 6944 11112 6996
rect 12256 6944 12308 6996
rect 15660 6944 15712 6996
rect 17224 6944 17276 6996
rect 17776 6944 17828 6996
rect 11888 6876 11940 6928
rect 11980 6876 12032 6928
rect 13176 6876 13228 6928
rect 14280 6876 14332 6928
rect 17500 6876 17552 6928
rect 8576 6808 8628 6860
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 6276 6740 6328 6792
rect 7472 6740 7524 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8944 6808 8996 6860
rect 9864 6808 9916 6860
rect 12900 6808 12952 6860
rect 9772 6740 9824 6792
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11704 6740 11756 6792
rect 3700 6672 3752 6724
rect 3792 6672 3844 6724
rect 2872 6604 2924 6656
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 7380 6604 7432 6656
rect 12256 6740 12308 6792
rect 13544 6808 13596 6860
rect 15568 6808 15620 6860
rect 15752 6808 15804 6860
rect 16212 6808 16264 6860
rect 17960 6808 18012 6860
rect 14832 6783 14884 6792
rect 9036 6604 9088 6656
rect 10232 6604 10284 6656
rect 11244 6604 11296 6656
rect 14004 6672 14056 6724
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 17500 6740 17552 6792
rect 13544 6604 13596 6656
rect 14372 6604 14424 6656
rect 15476 6672 15528 6724
rect 17132 6672 17184 6724
rect 15384 6604 15436 6656
rect 17408 6604 17460 6656
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 1676 6400 1728 6452
rect 2964 6400 3016 6452
rect 4896 6400 4948 6452
rect 6092 6443 6144 6452
rect 3056 6332 3108 6384
rect 6092 6409 6101 6443
rect 6101 6409 6135 6443
rect 6135 6409 6144 6443
rect 6092 6400 6144 6409
rect 6920 6400 6972 6452
rect 8576 6332 8628 6384
rect 11704 6400 11756 6452
rect 11980 6332 12032 6384
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 5724 6264 5776 6316
rect 6368 6264 6420 6316
rect 3516 6196 3568 6248
rect 8208 6264 8260 6316
rect 12716 6400 12768 6452
rect 12256 6332 12308 6384
rect 15108 6332 15160 6384
rect 15568 6332 15620 6384
rect 1584 6128 1636 6180
rect 1860 6128 1912 6180
rect 2228 6128 2280 6180
rect 3976 6128 4028 6180
rect 7380 6196 7432 6248
rect 7472 6196 7524 6248
rect 2688 6060 2740 6112
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3332 6060 3384 6112
rect 3516 6103 3568 6112
rect 3516 6069 3525 6103
rect 3525 6069 3559 6103
rect 3559 6069 3568 6103
rect 4252 6103 4304 6112
rect 3516 6060 3568 6069
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 5172 6128 5224 6180
rect 6276 6128 6328 6180
rect 6736 6128 6788 6180
rect 7840 6128 7892 6180
rect 8484 6128 8536 6180
rect 9036 6128 9088 6180
rect 10324 6196 10376 6248
rect 11980 6196 12032 6248
rect 12440 6196 12492 6248
rect 13176 6264 13228 6316
rect 13360 6196 13412 6248
rect 9312 6128 9364 6180
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 6460 6060 6512 6112
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 8300 6103 8352 6112
rect 7564 6060 7616 6069
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 8392 6060 8444 6112
rect 9128 6060 9180 6112
rect 9220 6060 9272 6112
rect 9772 6060 9824 6112
rect 11796 6128 11848 6180
rect 13636 6060 13688 6112
rect 14004 6196 14056 6248
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 15476 6264 15528 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 17132 6196 17184 6248
rect 14188 6060 14240 6112
rect 14648 6060 14700 6112
rect 16672 6060 16724 6112
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 17776 6060 17828 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 1492 5856 1544 5908
rect 3056 5856 3108 5908
rect 4620 5856 4672 5908
rect 2964 5788 3016 5840
rect 5632 5856 5684 5908
rect 6460 5856 6512 5908
rect 7472 5856 7524 5908
rect 8760 5856 8812 5908
rect 9220 5856 9272 5908
rect 11612 5856 11664 5908
rect 11796 5856 11848 5908
rect 12624 5856 12676 5908
rect 13176 5856 13228 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 14280 5856 14332 5908
rect 14740 5856 14792 5908
rect 15660 5856 15712 5908
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 2136 5720 2188 5772
rect 3700 5720 3752 5772
rect 5816 5763 5868 5772
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 2964 5652 3016 5704
rect 5448 5652 5500 5704
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 6184 5720 6236 5772
rect 6368 5720 6420 5772
rect 6920 5720 6972 5772
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 4344 5584 4396 5636
rect 8208 5627 8260 5636
rect 2504 5516 2556 5568
rect 2780 5516 2832 5568
rect 4712 5516 4764 5568
rect 5724 5516 5776 5568
rect 6276 5516 6328 5568
rect 6736 5516 6788 5568
rect 8208 5593 8217 5627
rect 8217 5593 8251 5627
rect 8251 5593 8260 5627
rect 8208 5584 8260 5593
rect 8392 5720 8444 5772
rect 8760 5652 8812 5704
rect 10324 5695 10376 5704
rect 8484 5584 8536 5636
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 9220 5584 9272 5636
rect 13912 5788 13964 5840
rect 14096 5788 14148 5840
rect 15476 5788 15528 5840
rect 16396 5788 16448 5840
rect 17316 5831 17368 5840
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 13176 5763 13228 5772
rect 13176 5729 13185 5763
rect 13185 5729 13219 5763
rect 13219 5729 13228 5763
rect 13176 5720 13228 5729
rect 17960 5763 18012 5772
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 14832 5695 14884 5704
rect 9588 5516 9640 5568
rect 12532 5584 12584 5636
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 13820 5584 13872 5636
rect 12256 5516 12308 5568
rect 12348 5516 12400 5568
rect 15016 5516 15068 5568
rect 17684 5652 17736 5704
rect 15568 5516 15620 5568
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 17868 5516 17920 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 5724 5312 5776 5364
rect 5816 5312 5868 5364
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 2596 5108 2648 5160
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 3884 5108 3936 5160
rect 1676 5040 1728 5092
rect 6276 5176 6328 5228
rect 6920 5176 6972 5228
rect 4068 5108 4120 5160
rect 5816 5108 5868 5160
rect 8208 5176 8260 5228
rect 11520 5312 11572 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 15200 5312 15252 5364
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 8852 5151 8904 5160
rect 5632 5040 5684 5092
rect 6092 5083 6144 5092
rect 6092 5049 6101 5083
rect 6101 5049 6135 5083
rect 6135 5049 6144 5083
rect 6092 5040 6144 5049
rect 7656 5040 7708 5092
rect 8208 5083 8260 5092
rect 8208 5049 8217 5083
rect 8217 5049 8251 5083
rect 8251 5049 8260 5083
rect 8208 5040 8260 5049
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 10324 5108 10376 5160
rect 12440 5244 12492 5296
rect 11796 5176 11848 5228
rect 13728 5176 13780 5228
rect 12348 5108 12400 5160
rect 12440 5151 12492 5160
rect 14832 5176 14884 5228
rect 12440 5117 12456 5151
rect 12456 5117 12490 5151
rect 12490 5117 12492 5151
rect 12440 5108 12492 5117
rect 15016 5151 15068 5160
rect 15016 5117 15025 5151
rect 15025 5117 15059 5151
rect 15059 5117 15068 5151
rect 15016 5108 15068 5117
rect 16672 5176 16724 5228
rect 16856 5176 16908 5228
rect 16948 5176 17000 5228
rect 17316 5108 17368 5160
rect 9772 5083 9824 5092
rect 9772 5049 9784 5083
rect 9784 5049 9824 5083
rect 9772 5040 9824 5049
rect 12072 5040 12124 5092
rect 14004 5040 14056 5092
rect 2412 4972 2464 5024
rect 3240 5015 3292 5024
rect 3240 4981 3249 5015
rect 3249 4981 3283 5015
rect 3283 4981 3292 5015
rect 3240 4972 3292 4981
rect 3884 4972 3936 5024
rect 4804 4972 4856 5024
rect 4896 4972 4948 5024
rect 8668 4972 8720 5024
rect 9128 4972 9180 5024
rect 10692 4972 10744 5024
rect 10876 5015 10928 5024
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 11612 4972 11664 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 11980 4972 12032 5024
rect 15752 4972 15804 5024
rect 16764 4972 16816 5024
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 3240 4768 3292 4820
rect 2688 4700 2740 4752
rect 6368 4768 6420 4820
rect 8484 4768 8536 4820
rect 9588 4768 9640 4820
rect 10416 4768 10468 4820
rect 11428 4768 11480 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 12164 4811 12216 4820
rect 12164 4777 12173 4811
rect 12173 4777 12207 4811
rect 12207 4777 12216 4811
rect 12164 4768 12216 4777
rect 12440 4768 12492 4820
rect 12716 4768 12768 4820
rect 13176 4768 13228 4820
rect 15384 4768 15436 4820
rect 5356 4700 5408 4752
rect 5632 4700 5684 4752
rect 4620 4632 4672 4684
rect 1584 4564 1636 4616
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 6552 4632 6604 4684
rect 8300 4700 8352 4752
rect 12900 4700 12952 4752
rect 13912 4743 13964 4752
rect 13912 4709 13921 4743
rect 13921 4709 13955 4743
rect 13955 4709 13964 4743
rect 16120 4768 16172 4820
rect 16764 4811 16816 4820
rect 16764 4777 16773 4811
rect 16773 4777 16807 4811
rect 16807 4777 16816 4811
rect 16764 4768 16816 4777
rect 18144 4768 18196 4820
rect 15752 4743 15804 4752
rect 13912 4700 13964 4709
rect 15752 4709 15761 4743
rect 15761 4709 15795 4743
rect 15795 4709 15804 4743
rect 15752 4700 15804 4709
rect 8208 4632 8260 4684
rect 8760 4632 8812 4684
rect 9496 4632 9548 4684
rect 10232 4607 10284 4616
rect 3148 4496 3200 4548
rect 3792 4496 3844 4548
rect 2596 4428 2648 4480
rect 6920 4496 6972 4548
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 11980 4564 12032 4616
rect 12440 4607 12492 4616
rect 8576 4496 8628 4548
rect 10692 4496 10744 4548
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 12624 4632 12676 4684
rect 14740 4632 14792 4684
rect 16120 4632 16172 4684
rect 17776 4675 17828 4684
rect 17776 4641 17785 4675
rect 17785 4641 17819 4675
rect 17819 4641 17828 4675
rect 17776 4632 17828 4641
rect 14004 4607 14056 4616
rect 6092 4428 6144 4480
rect 6552 4471 6604 4480
rect 6552 4437 6561 4471
rect 6561 4437 6595 4471
rect 6595 4437 6604 4471
rect 6552 4428 6604 4437
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 9772 4428 9824 4480
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 17684 4564 17736 4616
rect 18512 4564 18564 4616
rect 15200 4428 15252 4480
rect 15384 4428 15436 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 1216 4224 1268 4276
rect 1676 4156 1728 4208
rect 2044 4088 2096 4140
rect 2780 4156 2832 4208
rect 2596 4088 2648 4140
rect 1860 4020 1912 4072
rect 3148 4063 3200 4072
rect 3148 4029 3182 4063
rect 3182 4029 3200 4063
rect 3148 4020 3200 4029
rect 4436 4224 4488 4276
rect 7012 4224 7064 4276
rect 8208 4267 8260 4276
rect 8208 4233 8217 4267
rect 8217 4233 8251 4267
rect 8251 4233 8260 4267
rect 8208 4224 8260 4233
rect 12164 4224 12216 4276
rect 12900 4224 12952 4276
rect 15200 4224 15252 4276
rect 16856 4267 16908 4276
rect 16856 4233 16865 4267
rect 16865 4233 16899 4267
rect 16899 4233 16908 4267
rect 16856 4224 16908 4233
rect 5356 4088 5408 4140
rect 6000 4156 6052 4208
rect 14004 4156 14056 4208
rect 17776 4156 17828 4208
rect 6092 4131 6144 4140
rect 4896 4020 4948 4072
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 5724 4020 5776 4072
rect 6552 4088 6604 4140
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 6644 4020 6696 4072
rect 6920 4020 6972 4072
rect 2320 3952 2372 4004
rect 2688 3952 2740 4004
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 6736 3952 6788 4004
rect 7196 3952 7248 4004
rect 9404 4020 9456 4072
rect 9680 4020 9732 4072
rect 11152 4020 11204 4072
rect 12532 4088 12584 4140
rect 12716 4088 12768 4140
rect 9128 3995 9180 4004
rect 9128 3961 9162 3995
rect 9162 3961 9180 3995
rect 9128 3952 9180 3961
rect 9588 3952 9640 4004
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 10232 3927 10284 3936
rect 5632 3884 5684 3893
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 10416 3952 10468 4004
rect 13820 4020 13872 4072
rect 16948 4088 17000 4140
rect 17592 4088 17644 4140
rect 14556 4020 14608 4072
rect 15568 4020 15620 4072
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 17684 4020 17736 4072
rect 11980 3952 12032 4004
rect 11152 3884 11204 3936
rect 11336 3884 11388 3936
rect 17500 3952 17552 4004
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 16304 3927 16356 3936
rect 12440 3884 12492 3893
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 4344 3680 4396 3732
rect 388 3544 440 3596
rect 4712 3612 4764 3664
rect 6736 3680 6788 3732
rect 7564 3680 7616 3732
rect 9312 3680 9364 3732
rect 3608 3544 3660 3596
rect 4528 3544 4580 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 3792 3476 3844 3528
rect 4896 3476 4948 3528
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 6644 3612 6696 3664
rect 8392 3612 8444 3664
rect 5724 3544 5776 3596
rect 7840 3587 7892 3596
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 5356 3476 5408 3485
rect 8484 3476 8536 3528
rect 10232 3612 10284 3664
rect 10508 3612 10560 3664
rect 13268 3680 13320 3732
rect 13728 3680 13780 3732
rect 16120 3680 16172 3732
rect 16212 3680 16264 3732
rect 11520 3612 11572 3664
rect 10324 3587 10376 3596
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 11336 3544 11388 3596
rect 1768 3340 1820 3392
rect 2780 3340 2832 3392
rect 3608 3340 3660 3392
rect 4712 3340 4764 3392
rect 5172 3340 5224 3392
rect 8208 3408 8260 3460
rect 9404 3408 9456 3460
rect 16672 3612 16724 3664
rect 10232 3340 10284 3392
rect 11336 3340 11388 3392
rect 12716 3544 12768 3596
rect 13636 3544 13688 3596
rect 14004 3544 14056 3596
rect 11796 3476 11848 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 14280 3544 14332 3596
rect 17224 3612 17276 3664
rect 18052 3519 18104 3528
rect 16580 3408 16632 3460
rect 13820 3340 13872 3392
rect 16488 3340 16540 3392
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 3516 3136 3568 3188
rect 3700 3136 3752 3188
rect 5448 3136 5500 3188
rect 8576 3136 8628 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 10232 3136 10284 3188
rect 16212 3136 16264 3188
rect 18420 3136 18472 3188
rect 2320 3068 2372 3120
rect 1860 3000 1912 3052
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 3608 3000 3660 3052
rect 5632 3068 5684 3120
rect 10048 3068 10100 3120
rect 5172 3000 5224 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 7840 3000 7892 3052
rect 9128 3000 9180 3052
rect 9312 3000 9364 3052
rect 11336 3068 11388 3120
rect 11520 3068 11572 3120
rect 14096 3068 14148 3120
rect 16304 3111 16356 3120
rect 16304 3077 16313 3111
rect 16313 3077 16347 3111
rect 16347 3077 16356 3111
rect 16304 3068 16356 3077
rect 10508 3000 10560 3052
rect 11428 3000 11480 3052
rect 5540 2932 5592 2984
rect 7288 2932 7340 2984
rect 8024 2932 8076 2984
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 11704 2975 11756 2984
rect 2872 2864 2924 2916
rect 6184 2864 6236 2916
rect 6736 2864 6788 2916
rect 7564 2864 7616 2916
rect 8484 2864 8536 2916
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 11980 2932 12032 2984
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 14648 2932 14700 2984
rect 15292 2932 15344 2984
rect 16304 2932 16356 2984
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 2044 2796 2096 2848
rect 3332 2796 3384 2848
rect 4160 2839 4212 2848
rect 4160 2805 4169 2839
rect 4169 2805 4203 2839
rect 4203 2805 4212 2839
rect 4160 2796 4212 2805
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 5632 2796 5684 2848
rect 5816 2796 5868 2848
rect 6000 2796 6052 2848
rect 10140 2839 10192 2848
rect 10140 2805 10149 2839
rect 10149 2805 10183 2839
rect 10183 2805 10192 2839
rect 10140 2796 10192 2805
rect 10324 2796 10376 2848
rect 10508 2796 10560 2848
rect 11060 2839 11112 2848
rect 11060 2805 11069 2839
rect 11069 2805 11103 2839
rect 11103 2805 11112 2839
rect 11060 2796 11112 2805
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 12716 2796 12768 2848
rect 13176 2864 13228 2916
rect 14832 2864 14884 2916
rect 15660 2864 15712 2916
rect 16764 2907 16816 2916
rect 16764 2873 16773 2907
rect 16773 2873 16807 2907
rect 16807 2873 16816 2907
rect 16764 2864 16816 2873
rect 19432 2864 19484 2916
rect 13544 2796 13596 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2044 2592 2096 2644
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4160 2592 4212 2644
rect 4804 2592 4856 2644
rect 5080 2592 5132 2644
rect 5632 2592 5684 2644
rect 6184 2592 6236 2644
rect 5448 2524 5500 2576
rect 7840 2524 7892 2576
rect 9036 2592 9088 2644
rect 9772 2592 9824 2644
rect 10048 2592 10100 2644
rect 11060 2592 11112 2644
rect 11152 2592 11204 2644
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 2780 2456 2832 2508
rect 3608 2456 3660 2508
rect 4436 2456 4488 2508
rect 4712 2456 4764 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8852 2456 8904 2508
rect 9036 2499 9088 2508
rect 9036 2465 9045 2499
rect 9045 2465 9079 2499
rect 9079 2465 9088 2499
rect 9036 2456 9088 2465
rect 10876 2456 10928 2508
rect 12440 2592 12492 2644
rect 11612 2456 11664 2508
rect 12348 2456 12400 2508
rect 14464 2456 14516 2508
rect 16856 2592 16908 2644
rect 2412 2388 2464 2440
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 5724 2388 5776 2440
rect 6092 2388 6144 2440
rect 8760 2388 8812 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 11428 2388 11480 2440
rect 9404 2320 9456 2372
rect 10140 2320 10192 2372
rect 11244 2320 11296 2372
rect 12164 2388 12216 2440
rect 13912 2388 13964 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 16488 2320 16540 2372
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 3700 2048 3752 2100
rect 8392 2048 8444 2100
rect 1952 1980 2004 2032
rect 6920 1980 6972 2032
rect 3332 1300 3384 1352
rect 8668 1300 8720 1352
rect 4068 1164 4120 1216
rect 11888 1164 11940 1216
rect 3700 1028 3752 1080
rect 9220 1028 9272 1080
<< metal2 >>
rect 1674 16520 1730 17000
rect 3330 16824 3386 16833
rect 3330 16759 3386 16768
rect 3344 16590 3372 16759
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3790 16552 3846 16561
rect 1688 14074 1716 16520
rect 4986 16520 5042 17000
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 3790 16487 3846 16496
rect 3422 16144 3478 16153
rect 3422 16079 3478 16088
rect 3238 15464 3294 15473
rect 3238 15399 3294 15408
rect 2870 15192 2926 15201
rect 2870 15127 2926 15136
rect 2042 14784 2098 14793
rect 2042 14719 2098 14728
rect 2056 14550 2084 14719
rect 2044 14544 2096 14550
rect 2780 14544 2832 14550
rect 2044 14486 2096 14492
rect 2778 14512 2780 14521
rect 2832 14512 2834 14521
rect 2778 14447 2834 14456
rect 2778 14104 2834 14113
rect 1676 14068 1728 14074
rect 2778 14039 2834 14048
rect 1676 14010 1728 14016
rect 2792 13938 2820 14039
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 1860 13864 1912 13870
rect 1858 13832 1860 13841
rect 1912 13832 1914 13841
rect 1768 13796 1820 13802
rect 1858 13767 1914 13776
rect 1768 13738 1820 13744
rect 1780 13394 1808 13738
rect 2884 13530 2912 15127
rect 3252 14006 3280 15399
rect 3436 14618 3464 16079
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 14385 3372 14418
rect 3608 14408 3660 14414
rect 3330 14376 3386 14385
rect 3608 14350 3660 14356
rect 3330 14311 3386 14320
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3620 13870 3648 14350
rect 3804 14006 3832 16487
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 4080 14346 4108 15807
rect 5000 14618 5028 16520
rect 6472 14618 6500 16526
rect 8298 16520 8354 17000
rect 11610 16520 11666 17000
rect 14922 16520 14978 17000
rect 17866 16824 17922 16833
rect 17866 16759 17922 16768
rect 16118 16552 16174 16561
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3056 13864 3108 13870
rect 3054 13832 3056 13841
rect 3608 13864 3660 13870
rect 3108 13832 3110 13841
rect 3054 13767 3110 13776
rect 3606 13832 3608 13841
rect 3660 13832 3662 13841
rect 3606 13767 3662 13776
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3330 13424 3386 13433
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 2596 13388 2648 13394
rect 3330 13359 3332 13368
rect 2596 13330 2648 13336
rect 3384 13359 3386 13368
rect 3332 13330 3384 13336
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 10810 1440 13262
rect 1492 12708 1544 12714
rect 1492 12650 1544 12656
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1214 8664 1270 8673
rect 1214 8599 1270 8608
rect 1228 4282 1256 8599
rect 1308 6928 1360 6934
rect 1308 6870 1360 6876
rect 1320 4321 1348 6870
rect 1306 4312 1362 4321
rect 1216 4276 1268 4282
rect 1306 4247 1362 4256
rect 1216 4218 1268 4224
rect 1412 3913 1440 9318
rect 1504 5914 1532 12650
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1596 11014 1624 11630
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10606 1624 10950
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 9926 1624 10542
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 8838 1624 9862
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8430 1624 8774
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1674 8392 1730 8401
rect 1596 7954 1624 8366
rect 1674 8327 1676 8336
rect 1728 8327 1730 8336
rect 1676 8298 1728 8304
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6186 1624 6734
rect 1688 6458 1716 6802
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1584 6180 1636 6186
rect 1584 6122 1636 6128
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1596 5166 1624 6122
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1596 4622 1624 5102
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1584 4616 1636 4622
rect 1504 4576 1584 4604
rect 1398 3904 1454 3913
rect 1398 3839 1454 3848
rect 1504 3754 1532 4576
rect 1584 4558 1636 4564
rect 1688 4214 1716 5034
rect 1676 4208 1728 4214
rect 1676 4150 1728 4156
rect 1412 3726 1532 3754
rect 388 3596 440 3602
rect 388 3538 440 3544
rect 400 480 428 3538
rect 1412 3534 1440 3726
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1400 3528 1452 3534
rect 1214 3496 1270 3505
rect 1400 3470 1452 3476
rect 1214 3431 1270 3440
rect 1228 480 1256 3431
rect 1398 2680 1454 2689
rect 1596 2650 1624 3567
rect 1780 3398 1808 13330
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2056 12782 2084 13126
rect 2044 12776 2096 12782
rect 2412 12776 2464 12782
rect 2044 12718 2096 12724
rect 2332 12736 2412 12764
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1872 7426 1900 12582
rect 2148 12442 2176 12582
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1964 10674 1992 11154
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1964 7546 1992 10066
rect 2056 9654 2084 12242
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10062 2176 10610
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2148 9586 2176 9998
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2134 8120 2190 8129
rect 2134 8055 2190 8064
rect 2148 7721 2176 8055
rect 2134 7712 2190 7721
rect 2134 7647 2190 7656
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1872 7398 1992 7426
rect 2148 7410 2176 7647
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1872 6866 1900 7278
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1872 4078 1900 6122
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1872 3058 1900 3878
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1398 2615 1454 2624
rect 1584 2644 1636 2650
rect 1412 2514 1440 2615
rect 1584 2586 1636 2592
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1964 2038 1992 7398
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2042 7032 2098 7041
rect 2042 6967 2098 6976
rect 2056 4146 2084 6967
rect 2148 5896 2176 7346
rect 2240 7342 2268 12106
rect 2332 10130 2360 12736
rect 2412 12718 2464 12724
rect 2516 12238 2544 13194
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2424 10266 2452 12174
rect 2516 11694 2544 12174
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2516 11354 2544 11630
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2608 10266 2636 13330
rect 3792 13184 3844 13190
rect 2962 13152 3018 13161
rect 3792 13126 3844 13132
rect 2962 13087 3018 13096
rect 2976 12986 3004 13087
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2700 11898 2728 12786
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2700 10606 2728 11834
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2686 10296 2742 10305
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2596 10260 2648 10266
rect 2686 10231 2742 10240
rect 2596 10202 2648 10208
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 6186 2268 7142
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2332 6089 2360 7210
rect 2424 7206 2452 8910
rect 2516 8634 2544 9318
rect 2608 9178 2636 9522
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2700 9042 2728 10231
rect 2792 9489 2820 12174
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2870 11384 2926 11393
rect 2870 11319 2926 11328
rect 2778 9480 2834 9489
rect 2778 9415 2834 9424
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2596 8424 2648 8430
rect 2700 8378 2728 8978
rect 2648 8372 2728 8378
rect 2596 8366 2728 8372
rect 2608 8350 2728 8366
rect 2700 8090 2728 8350
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2700 7970 2728 8026
rect 2608 7942 2728 7970
rect 2608 7410 2636 7942
rect 2686 7848 2742 7857
rect 2686 7783 2742 7792
rect 2700 7546 2728 7783
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2594 7304 2650 7313
rect 2594 7239 2650 7248
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2504 6860 2556 6866
rect 2424 6820 2504 6848
rect 2318 6080 2374 6089
rect 2318 6015 2374 6024
rect 2148 5868 2268 5896
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2650 2084 2790
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 2148 480 2176 5714
rect 2240 3108 2268 5868
rect 2332 4010 2360 6015
rect 2424 5030 2452 6820
rect 2504 6802 2556 6808
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2320 3120 2372 3126
rect 2240 3080 2320 3108
rect 2320 3062 2372 3068
rect 2424 3058 2452 4966
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2424 2446 2452 2994
rect 2516 2938 2544 5510
rect 2608 5166 2636 7239
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5710 2728 6054
rect 2792 5817 2820 8327
rect 2884 7478 2912 11319
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2872 6656 2924 6662
rect 2976 6633 3004 11494
rect 3068 6866 3096 12786
rect 3804 12753 3832 13126
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4344 12776 4396 12782
rect 3790 12744 3846 12753
rect 3790 12679 3846 12688
rect 4264 12736 4344 12764
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3160 12442 3188 12582
rect 3330 12472 3386 12481
rect 3148 12436 3200 12442
rect 3330 12407 3386 12416
rect 3148 12378 3200 12384
rect 3344 12306 3372 12407
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3344 12209 3372 12242
rect 3330 12200 3386 12209
rect 3330 12135 3386 12144
rect 3146 11792 3202 11801
rect 3146 11727 3202 11736
rect 3160 10538 3188 11727
rect 3436 11121 3464 12310
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3698 12064 3754 12073
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3160 9722 3188 10474
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2872 6598 2924 6604
rect 2962 6624 3018 6633
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2700 4758 2728 5646
rect 2792 5574 2820 5743
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2608 4146 2636 4422
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2700 3108 2728 3946
rect 2792 3738 2820 4150
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2792 3398 2820 3674
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2884 3233 2912 6598
rect 2962 6559 3018 6568
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2976 5846 3004 6394
rect 3068 6390 3096 6802
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5914 3096 6054
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2870 3224 2926 3233
rect 2870 3159 2926 3168
rect 2700 3080 2912 3108
rect 2516 2910 2820 2938
rect 2884 2922 2912 3080
rect 2792 2514 2820 2910
rect 2872 2916 2924 2922
rect 2976 2904 3004 5646
rect 3160 4672 3188 8774
rect 3252 5953 3280 10950
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 7834 3372 10406
rect 3436 10198 3464 10950
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3436 8906 3464 9318
rect 3528 9178 3556 9318
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3344 7806 3556 7834
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3330 7304 3386 7313
rect 3330 7239 3386 7248
rect 3344 7206 3372 7239
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3238 5944 3294 5953
rect 3238 5879 3294 5888
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 4826 3280 4966
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3068 4644 3188 4672
rect 3068 3924 3096 4644
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3160 4078 3188 4490
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3068 3896 3188 3924
rect 2976 2876 3096 2904
rect 2872 2858 2924 2864
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 3068 480 3096 2876
rect 386 0 442 480
rect 1214 0 1270 480
rect 2134 0 2190 480
rect 3054 0 3110 480
rect 3160 241 3188 3896
rect 3344 2854 3372 6054
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3330 2680 3386 2689
rect 3330 2615 3332 2624
rect 3384 2615 3386 2624
rect 3332 2586 3384 2592
rect 3436 1873 3464 7686
rect 3528 6254 3556 7806
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 3194 3556 6054
rect 3620 3602 3648 12038
rect 3698 11999 3754 12008
rect 3712 11898 3740 11999
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 9926 3740 10406
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3698 9344 3754 9353
rect 3698 9279 3754 9288
rect 3712 8498 3740 9279
rect 3804 8634 3832 12106
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 4264 11778 4292 12736
rect 4344 12718 4396 12724
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12442 4568 12650
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4172 11750 4292 11778
rect 4172 11218 4200 11750
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4172 11082 4200 11154
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4264 10810 4292 11630
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4356 11286 4384 11562
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 4080 10470 4108 10639
rect 4160 10600 4212 10606
rect 4356 10588 4384 11222
rect 4212 10560 4384 10588
rect 4160 10542 4212 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4172 10062 4200 10542
rect 4342 10432 4398 10441
rect 4342 10367 4398 10376
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4356 9761 4384 10367
rect 4342 9752 4398 9761
rect 4342 9687 4398 9696
rect 4448 9654 4476 12242
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4436 9648 4488 9654
rect 3974 9616 4030 9625
rect 4436 9590 4488 9596
rect 3974 9551 4030 9560
rect 4252 9580 4304 9586
rect 3988 9450 4016 9551
rect 4252 9522 4304 9528
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 4172 9353 4200 9454
rect 4158 9344 4214 9353
rect 4158 9279 4214 9288
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3804 8022 3832 8570
rect 4066 8392 4122 8401
rect 4264 8362 4292 9522
rect 4356 9489 4384 9522
rect 4342 9480 4398 9489
rect 4342 9415 4398 9424
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 8634 4384 9318
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4066 8327 4122 8336
rect 4252 8356 4304 8362
rect 4080 8294 4108 8327
rect 4252 8298 4304 8304
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 4080 7954 4108 8230
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7546 4292 7890
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 7478 4384 7686
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4448 7410 4476 8298
rect 4540 8090 4568 12174
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3712 6322 3740 6666
rect 3804 6361 3832 6666
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 3790 6352 3846 6361
rect 3700 6316 3752 6322
rect 3790 6287 3846 6296
rect 3700 6258 3752 6264
rect 4264 6202 4292 6598
rect 3976 6180 4028 6186
rect 4264 6174 4384 6202
rect 3976 6122 4028 6128
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3620 3058 3648 3334
rect 3712 3194 3740 5714
rect 3988 5681 4016 6122
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4554 3832 5170
rect 3884 5160 3936 5166
rect 3882 5128 3884 5137
rect 4068 5160 4120 5166
rect 3936 5128 3938 5137
rect 4068 5102 4120 5108
rect 3882 5063 3938 5072
rect 3884 5024 3936 5030
rect 4080 5001 4108 5102
rect 3884 4966 3936 4972
rect 4066 4992 4122 5001
rect 3896 4593 3924 4966
rect 4066 4927 4122 4936
rect 3882 4584 3938 4593
rect 3792 4548 3844 4554
rect 3882 4519 3938 4528
rect 3792 4490 3844 4496
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3608 3052 3660 3058
rect 3528 3012 3608 3040
rect 3528 2446 3556 3012
rect 3608 2994 3660 3000
rect 3606 2544 3662 2553
rect 3606 2479 3608 2488
rect 3660 2479 3662 2488
rect 3608 2450 3660 2456
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3698 2272 3754 2281
rect 3698 2207 3754 2216
rect 3712 2106 3740 2207
rect 3700 2100 3752 2106
rect 3700 2042 3752 2048
rect 3422 1864 3478 1873
rect 3422 1799 3478 1808
rect 3804 1442 3832 3470
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4066 2952 4122 2961
rect 4264 2938 4292 6054
rect 4356 5642 4384 6174
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4448 5545 4476 7142
rect 4540 6633 4568 7822
rect 4632 7002 4660 12786
rect 4724 9450 4752 12922
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4816 11694 4844 12786
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4816 9330 4844 10950
rect 4724 9302 4844 9330
rect 4724 9110 4752 9302
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4724 8537 4752 9046
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4710 8528 4766 8537
rect 4710 8463 4766 8472
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7546 4752 7822
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4526 6624 4582 6633
rect 4526 6559 4582 6568
rect 4434 5536 4490 5545
rect 4434 5471 4490 5480
rect 4448 4434 4476 5471
rect 4356 4406 4476 4434
rect 4356 3738 4384 4406
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4122 2910 4292 2938
rect 4066 2887 4122 2896
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4172 2650 4200 2790
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4448 2514 4476 4218
rect 4540 3602 4568 6559
rect 4632 5914 4660 6802
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4724 6361 4752 6734
rect 4710 6352 4766 6361
rect 4710 6287 4766 6296
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4618 5400 4674 5409
rect 4618 5335 4674 5344
rect 4632 4690 4660 5335
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4632 2553 4660 4626
rect 4724 3670 4752 5510
rect 4816 5030 4844 8774
rect 4908 7449 4936 12378
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5000 10305 5028 11018
rect 4986 10296 5042 10305
rect 4986 10231 5042 10240
rect 5184 10062 5212 14418
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5276 9722 5304 13330
rect 5460 10810 5488 13874
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5552 11762 5580 12854
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11286 5580 11494
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5368 9994 5396 10202
rect 5460 10198 5488 10746
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8838 5028 9318
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4894 7440 4950 7449
rect 4894 7375 4950 7384
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4908 6798 4936 7278
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6458 4936 6734
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4894 5128 4950 5137
rect 4894 5063 4950 5072
rect 4908 5030 4936 5063
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4894 4584 4950 4593
rect 4894 4519 4950 4528
rect 4908 4078 4936 4519
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4618 2544 4674 2553
rect 4436 2508 4488 2514
rect 4724 2514 4752 3334
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4816 2650 4844 2790
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4618 2479 4674 2488
rect 4712 2508 4764 2514
rect 4436 2450 4488 2456
rect 4712 2450 4764 2456
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3804 1414 4016 1442
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 513 3372 1294
rect 3700 1080 3752 1086
rect 3700 1022 3752 1028
rect 3712 921 3740 1022
rect 3698 912 3754 921
rect 3698 847 3754 856
rect 3330 504 3386 513
rect 3988 480 4016 1414
rect 4068 1216 4120 1222
rect 4066 1184 4068 1193
rect 4120 1184 4122 1193
rect 4066 1119 4122 1128
rect 4908 480 4936 3470
rect 5000 1601 5028 7754
rect 5092 7585 5120 9658
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5078 7576 5134 7585
rect 5078 7511 5134 7520
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5092 2650 5120 6938
rect 5184 6866 5212 9386
rect 5276 9178 5304 9658
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5184 4622 5212 6122
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 3058 5212 3334
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5276 2961 5304 8910
rect 5368 8362 5396 8910
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5460 8242 5488 9998
rect 5552 9450 5580 10202
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5368 8214 5488 8242
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5368 4865 5396 8214
rect 5552 7886 5580 8230
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5644 7698 5672 13942
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13530 6040 13670
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5828 12986 5856 13330
rect 6288 13326 6316 13874
rect 8036 13870 8064 14418
rect 8312 13938 8340 16520
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 11624 13870 11652 16520
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 13450 13968 13506 13977
rect 14936 13938 14964 16520
rect 16118 16487 16174 16496
rect 15658 16144 15714 16153
rect 15658 16079 15714 16088
rect 15566 15464 15622 15473
rect 15566 15399 15622 15408
rect 15198 15192 15254 15201
rect 15198 15127 15254 15136
rect 13450 13903 13506 13912
rect 14924 13932 14976 13938
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7300 13530 7328 13670
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5736 12442 5764 12582
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5828 11642 5856 12582
rect 5920 11830 5948 13262
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5736 11614 5856 11642
rect 5736 11218 5764 11614
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5828 10146 5856 11494
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 5920 10606 5948 11222
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6012 10266 6040 12854
rect 6104 11286 6132 13262
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5828 10118 6040 10146
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5736 8514 5764 9930
rect 5828 9178 5856 9998
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5908 8560 5960 8566
rect 5736 8486 5856 8514
rect 5908 8502 5960 8508
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8090 5764 8366
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5552 7670 5672 7698
rect 5446 6216 5502 6225
rect 5446 6151 5502 6160
rect 5460 5710 5488 6151
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5354 4856 5410 4865
rect 5354 4791 5410 4800
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5368 4146 5396 4694
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5368 3534 5396 4082
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5368 3058 5396 3470
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5262 2952 5318 2961
rect 5262 2887 5318 2896
rect 5276 2854 5304 2887
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5460 2582 5488 3130
rect 5552 2990 5580 7670
rect 5828 6497 5856 8486
rect 5814 6488 5870 6497
rect 5814 6423 5870 6432
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 6202 5764 6258
rect 5644 6174 5764 6202
rect 5644 5914 5672 6174
rect 5632 5908 5684 5914
rect 5828 5896 5856 6423
rect 5632 5850 5684 5856
rect 5736 5868 5856 5896
rect 5736 5574 5764 5868
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5828 5370 5856 5714
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5644 4758 5672 5034
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5736 4321 5764 5306
rect 5920 5273 5948 8502
rect 6012 8022 6040 10118
rect 6104 8294 6132 11086
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6000 8016 6052 8022
rect 5998 7984 6000 7993
rect 6052 7984 6054 7993
rect 5998 7919 6054 7928
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7478 6040 7686
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5906 5264 5962 5273
rect 5906 5199 5962 5208
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5722 4312 5778 4321
rect 5722 4247 5778 4256
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3126 5672 3878
rect 5736 3602 5764 4014
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2650 5672 2790
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5736 2446 5764 3538
rect 5828 2854 5856 5102
rect 6012 4214 6040 7142
rect 6104 7041 6132 8230
rect 6090 7032 6146 7041
rect 6090 6967 6146 6976
rect 6196 6905 6224 10610
rect 6288 10033 6316 11630
rect 6380 10674 6408 12174
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6274 10024 6330 10033
rect 6274 9959 6330 9968
rect 6288 9178 6316 9959
rect 6380 9722 6408 10610
rect 6472 10266 6500 12038
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6380 9450 6408 9658
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6366 9344 6422 9353
rect 6366 9279 6422 9288
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6380 9110 6408 9279
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 8566 6408 8774
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6182 6896 6238 6905
rect 6092 6860 6144 6866
rect 6182 6831 6238 6840
rect 6092 6802 6144 6808
rect 6104 6458 6132 6802
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6104 5710 6132 6394
rect 6196 5778 6224 6831
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6186 6316 6734
rect 6380 6322 6408 8502
rect 6472 7834 6500 9930
rect 6564 8838 6592 13262
rect 7116 12850 7144 13262
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7392 12714 7420 13738
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7484 12986 7512 13466
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6552 8832 6604 8838
rect 6656 8809 6684 12242
rect 6748 10248 6776 12582
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6748 10220 6868 10248
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9586 6776 10066
rect 6840 9897 6868 10220
rect 7300 10198 7328 12106
rect 7484 11762 7512 12786
rect 7576 12458 7604 13126
rect 7760 12646 7788 13194
rect 8036 12866 8064 13806
rect 11624 13546 11652 13806
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 11532 13518 11652 13546
rect 11888 13524 11940 13530
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 7852 12838 8064 12866
rect 9312 12844 9364 12850
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7576 12430 7788 12458
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7668 12073 7696 12242
rect 7654 12064 7710 12073
rect 7654 11999 7710 12008
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 11286 7696 11562
rect 7760 11286 7788 12430
rect 7852 11558 7880 12838
rect 9312 12786 9364 12792
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 10282 7512 10542
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7392 10254 7512 10282
rect 7288 10192 7340 10198
rect 7102 10160 7158 10169
rect 7288 10134 7340 10140
rect 7102 10095 7158 10104
rect 7116 10062 7144 10095
rect 7104 10056 7156 10062
rect 7392 10044 7420 10254
rect 7472 10056 7524 10062
rect 7392 10016 7472 10044
rect 7104 9998 7156 10004
rect 7472 9998 7524 10004
rect 6826 9888 6882 9897
rect 6826 9823 6882 9832
rect 7194 9752 7250 9761
rect 7194 9687 7250 9696
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 9178 6776 9522
rect 7208 9450 7236 9687
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7392 9217 7420 9386
rect 7484 9382 7512 9998
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7378 9208 7434 9217
rect 6736 9172 6788 9178
rect 7576 9178 7604 9862
rect 7668 9178 7696 10474
rect 7378 9143 7434 9152
rect 7564 9172 7616 9178
rect 6736 9114 6788 9120
rect 7564 9114 7616 9120
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8832 7340 8838
rect 6552 8774 6604 8780
rect 6642 8800 6698 8809
rect 7288 8774 7340 8780
rect 6642 8735 6698 8744
rect 6656 8129 6684 8735
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6642 8120 6698 8129
rect 6886 8112 7182 8132
rect 6642 8055 6698 8064
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6564 7834 6592 7890
rect 6472 7806 6592 7834
rect 6472 6882 6500 7806
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6564 7002 6592 7346
rect 6656 7206 6684 7958
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 7478 6868 7754
rect 6828 7472 6880 7478
rect 7208 7449 7236 7822
rect 6828 7414 6880 7420
rect 7194 7440 7250 7449
rect 7194 7375 7250 7384
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6472 6854 6592 6882
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6380 5778 6408 6054
rect 6472 5914 6500 6054
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6090 5264 6146 5273
rect 6288 5234 6316 5510
rect 6090 5199 6146 5208
rect 6276 5228 6328 5234
rect 6104 5098 6132 5199
rect 6276 5170 6328 5176
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6380 4826 6408 5714
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6564 4690 6592 6854
rect 6656 5409 6684 7142
rect 6748 6186 6776 7278
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6932 6458 6960 6802
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6748 5692 6776 6122
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5704 6880 5710
rect 6748 5664 6828 5692
rect 6748 5574 6776 5664
rect 6828 5646 6880 5652
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6642 5400 6698 5409
rect 6642 5335 6698 5344
rect 6748 4808 6776 5510
rect 6932 5234 6960 5714
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6748 4780 6960 4808
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6932 4554 6960 4780
rect 7194 4720 7250 4729
rect 7194 4655 7250 4664
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 6012 2854 6040 4150
rect 6104 4146 6132 4422
rect 6564 4146 6592 4422
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6932 4078 6960 4490
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4282 7052 4422
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6656 3670 6684 4014
rect 7208 4010 7236 4655
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 6748 3738 6776 3946
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 7300 2990 7328 8774
rect 7392 6662 7420 8910
rect 7484 8634 7512 8978
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7760 8430 7788 10746
rect 7852 10577 7880 11086
rect 7838 10568 7894 10577
rect 7838 10503 7894 10512
rect 7852 9110 7880 10503
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7944 8634 7972 12718
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 11626 8064 12650
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7930 8528 7986 8537
rect 7930 8463 7986 8472
rect 7944 8430 7972 8463
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7930 7984 7986 7993
rect 7748 7948 7800 7954
rect 7930 7919 7932 7928
rect 7748 7890 7800 7896
rect 7984 7919 7986 7928
rect 7932 7890 7984 7896
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6798 7512 7686
rect 7654 7576 7710 7585
rect 7654 7511 7710 7520
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6254 7420 6598
rect 7470 6488 7526 6497
rect 7470 6423 7526 6432
rect 7484 6254 7512 6423
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7484 5914 7512 6054
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7576 3738 7604 6054
rect 7668 5098 7696 7511
rect 7760 7002 7788 7890
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7852 6186 7880 6734
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7852 3058 7880 3538
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6196 2650 6224 2858
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 5724 2440 5776 2446
rect 6092 2440 6144 2446
rect 5724 2382 5776 2388
rect 5828 2400 6092 2428
rect 4986 1592 5042 1601
rect 4986 1527 5042 1536
rect 5828 480 5856 2400
rect 6092 2382 6144 2388
rect 6748 480 6776 2858
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6932 2038 6960 2450
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 7576 480 7604 2858
rect 7944 2666 7972 7890
rect 8036 2990 8064 10406
rect 8128 7274 8156 12038
rect 8220 11354 8248 12582
rect 8482 12200 8538 12209
rect 8482 12135 8538 12144
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 9382 8248 10066
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 8498 8248 9318
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8312 7206 8340 11494
rect 8496 10810 8524 12135
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8588 11150 8616 11698
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8404 9897 8432 10202
rect 8390 9888 8446 9897
rect 8390 9823 8446 9832
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 7274 8432 8774
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 8294 8524 8434
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 7750 8524 8230
rect 8588 8090 8616 9386
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8574 7440 8630 7449
rect 8574 7375 8630 7384
rect 8588 7342 8616 7375
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8576 7336 8628 7342
rect 8680 7313 8708 12582
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8772 11694 8800 12106
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11354 8892 11494
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8956 9874 8984 12174
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9140 11354 9168 11698
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9036 11076 9088 11082
rect 9140 11064 9168 11290
rect 9088 11036 9168 11064
rect 9036 11018 9088 11024
rect 9048 10606 9076 11018
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8576 7278 8628 7284
rect 8666 7304 8722 7313
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8220 5642 8248 6258
rect 8404 6225 8432 7210
rect 8390 6216 8446 6225
rect 8496 6186 8524 7278
rect 8666 7239 8722 7248
rect 8772 7188 8800 9046
rect 8864 9042 8892 9862
rect 8956 9846 9076 9874
rect 9048 9353 9076 9846
rect 9140 9518 9168 10678
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9034 9344 9090 9353
rect 9034 9279 9090 9288
rect 9048 9110 9076 9279
rect 9232 9178 9260 12582
rect 9324 12238 9352 12786
rect 9692 12442 9720 13126
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 9128 8968 9180 8974
rect 8942 8936 8998 8945
rect 9128 8910 9180 8916
rect 8942 8871 8998 8880
rect 8956 8566 8984 8871
rect 9140 8809 9168 8910
rect 9324 8838 9352 12174
rect 9416 11694 9444 12174
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 10674 9536 11494
rect 9692 11150 9720 11766
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9600 10606 9628 10950
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10198 9444 10406
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9692 10062 9720 11086
rect 9784 10169 9812 13398
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11257 9904 11494
rect 9862 11248 9918 11257
rect 9862 11183 9918 11192
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9770 10160 9826 10169
rect 9770 10095 9826 10104
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10244 9654 10272 13262
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11694 10364 12038
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10520 10996 10548 12242
rect 10612 11626 10640 12582
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10600 11008 10652 11014
rect 10520 10968 10600 10996
rect 10520 10538 10548 10968
rect 10600 10950 10652 10956
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10232 9648 10284 9654
rect 10520 9625 10548 10066
rect 10232 9590 10284 9596
rect 10506 9616 10562 9625
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9081 9444 9454
rect 9680 9104 9732 9110
rect 9402 9072 9458 9081
rect 9680 9046 9732 9052
rect 9402 9007 9458 9016
rect 9312 8832 9364 8838
rect 9126 8800 9182 8809
rect 9312 8774 9364 8780
rect 9126 8735 9182 8744
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7857 8984 8026
rect 8942 7848 8998 7857
rect 8942 7783 8998 7792
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8680 7160 8800 7188
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 6390 8616 6802
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8574 6216 8630 6225
rect 8390 6151 8446 6160
rect 8484 6180 8536 6186
rect 8404 6118 8432 6151
rect 8574 6151 8630 6160
rect 8484 6122 8536 6128
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8220 5234 8248 5578
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8220 4865 8248 5034
rect 8206 4856 8262 4865
rect 8206 4791 8262 4800
rect 8312 4758 8340 6054
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8404 5273 8432 5714
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8390 5264 8446 5273
rect 8496 5234 8524 5578
rect 8588 5545 8616 6151
rect 8680 5794 8708 7160
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8758 5944 8814 5953
rect 8758 5879 8760 5888
rect 8812 5879 8814 5888
rect 8760 5850 8812 5856
rect 8758 5808 8814 5817
rect 8680 5766 8758 5794
rect 8758 5743 8814 5752
rect 8772 5710 8800 5743
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8574 5536 8630 5545
rect 8574 5471 8630 5480
rect 8574 5400 8630 5409
rect 8574 5335 8630 5344
rect 8390 5199 8446 5208
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4826 8524 5170
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8220 4282 8248 4626
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8220 3466 8248 4218
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7852 2638 7972 2666
rect 7852 2582 7880 2638
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8404 2106 8432 3606
rect 8496 3534 8524 4762
rect 8588 4554 8616 5335
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8588 3194 8616 4490
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8496 480 8524 2858
rect 8680 1358 8708 4966
rect 8772 4690 8800 5646
rect 8864 5166 8892 6938
rect 8942 6896 8998 6905
rect 8942 6831 8944 6840
rect 8996 6831 8998 6840
rect 8944 6802 8996 6808
rect 9048 6746 9076 7686
rect 8956 6718 9076 6746
rect 8852 5160 8904 5166
rect 8850 5128 8852 5137
rect 8904 5128 8906 5137
rect 8850 5063 8906 5072
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8758 4312 8814 4321
rect 8758 4247 8814 4256
rect 8772 2446 8800 4247
rect 8956 3602 8984 6718
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9310 6624 9366 6633
rect 9048 6186 9076 6598
rect 9310 6559 9366 6568
rect 9324 6186 9352 6559
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9140 5030 9168 6054
rect 9232 5914 9260 6054
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9232 4593 9260 5578
rect 9416 5273 9444 8230
rect 9600 7886 9628 8298
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9402 5264 9458 5273
rect 9402 5199 9458 5208
rect 9034 4584 9090 4593
rect 9034 4519 9090 4528
rect 9218 4584 9274 4593
rect 9218 4519 9274 4528
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9048 2990 9076 4519
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 9140 3058 9168 3946
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9036 2644 9088 2650
rect 8864 2604 9036 2632
rect 8864 2514 8892 2604
rect 9036 2586 9088 2592
rect 9034 2544 9090 2553
rect 8852 2508 8904 2514
rect 9034 2479 9036 2488
rect 8852 2450 8904 2456
rect 9088 2479 9090 2488
rect 9036 2450 9088 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 9232 1086 9260 4422
rect 9416 4162 9444 5199
rect 9508 4690 9536 7142
rect 9600 6934 9628 7686
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9692 6769 9720 9046
rect 10244 9042 10272 9590
rect 10506 9551 10562 9560
rect 10414 9208 10470 9217
rect 10414 9143 10470 9152
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10244 8616 10272 8978
rect 10428 8974 10456 9143
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10060 8588 10272 8616
rect 10060 8430 10088 8588
rect 10336 8566 10364 8774
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10244 8294 10272 8434
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10244 7410 10272 8230
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6798 9812 7142
rect 9862 6896 9918 6905
rect 9862 6831 9864 6840
rect 9916 6831 9918 6840
rect 9864 6802 9916 6808
rect 9772 6792 9824 6798
rect 9678 6760 9734 6769
rect 9772 6734 9824 6740
rect 9678 6695 9734 6704
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 4826 9628 5510
rect 9784 5098 9812 6054
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 10244 4622 10272 6598
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10336 5710 10364 6190
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10336 5166 10364 5646
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9324 4134 9444 4162
rect 9324 3738 9352 4134
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3466 9444 4014
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9324 2446 9352 2994
rect 9600 2961 9628 3946
rect 9692 3194 9720 4014
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9586 2952 9642 2961
rect 9586 2887 9642 2896
rect 9784 2650 9812 4422
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3670 10272 3878
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10336 3602 10364 5102
rect 10428 4826 10456 8026
rect 10520 5545 10548 9551
rect 10612 7818 10640 10474
rect 10704 10470 10732 12854
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10888 12594 10916 12786
rect 10980 12782 11008 13126
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10888 12566 11008 12594
rect 10980 12238 11008 12566
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9178 10732 9318
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10704 7546 10732 8978
rect 10796 7954 10824 12106
rect 10888 10810 10916 12174
rect 10980 11558 11008 12174
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10980 11218 11008 11494
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 11072 10674 11100 11630
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11072 10266 11100 10610
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10888 10010 10916 10202
rect 11164 10130 11192 13330
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12102 11468 13262
rect 11532 12730 11560 13518
rect 11888 13466 11940 13472
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12850 11652 13262
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12918 11836 13194
rect 11900 12918 11928 13466
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11612 12844 11664 12850
rect 11664 12804 11744 12832
rect 11612 12786 11664 12792
rect 11532 12702 11652 12730
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11532 11286 11560 12310
rect 11624 12306 11652 12702
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 10888 9982 11100 10010
rect 11072 9926 11100 9982
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10980 9450 11008 9862
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10980 8974 11008 9386
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10888 8838 10916 8910
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 8362 10916 8774
rect 10980 8634 11008 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11072 8362 11100 9590
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11058 7848 11114 7857
rect 10980 7721 11008 7822
rect 11058 7783 11060 7792
rect 11112 7783 11114 7792
rect 11060 7754 11112 7760
rect 10966 7712 11022 7721
rect 10966 7647 11022 7656
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10796 7342 10824 7482
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10796 6798 10824 7278
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 7002 11100 7142
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10506 5536 10562 5545
rect 10506 5471 10562 5480
rect 10690 5128 10746 5137
rect 10690 5063 10746 5072
rect 10704 5030 10732 5063
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10704 4457 10732 4490
rect 10690 4448 10746 4457
rect 10690 4383 10746 4392
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10336 3505 10364 3538
rect 10322 3496 10378 3505
rect 10322 3431 10378 3440
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 10244 3194 10272 3334
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10060 2650 10088 3062
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 10152 2378 10180 2790
rect 10336 2446 10364 2790
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 9220 1080 9272 1086
rect 9220 1022 9272 1028
rect 9416 480 9444 2314
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10428 1442 10456 3946
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10520 3058 10548 3606
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10520 2854 10548 2994
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10888 2514 10916 4966
rect 11164 4078 11192 9318
rect 11348 9217 11376 9522
rect 11440 9382 11468 10610
rect 11624 10470 11652 11834
rect 11716 11694 11744 12804
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11612 10464 11664 10470
rect 11532 10424 11612 10452
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11334 9208 11390 9217
rect 11334 9143 11390 9152
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11256 6662 11284 7958
rect 11348 6984 11376 9143
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8090 11468 8978
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11348 6956 11468 6984
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11440 5953 11468 6956
rect 11426 5944 11482 5953
rect 11426 5879 11482 5888
rect 11440 4826 11468 5879
rect 11532 5370 11560 10424
rect 11612 10406 11664 10412
rect 11612 9376 11664 9382
rect 11610 9344 11612 9353
rect 11664 9344 11666 9353
rect 11610 9279 11666 9288
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11624 7410 11652 8978
rect 11716 8430 11744 11222
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10810 11836 11086
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11704 7404 11756 7410
rect 11900 7392 11928 12038
rect 12360 10674 12388 12718
rect 12820 12714 12848 12922
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12360 10266 12388 10610
rect 12544 10606 12572 11018
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12532 10600 12584 10606
rect 12438 10568 12494 10577
rect 12532 10542 12584 10548
rect 12438 10503 12494 10512
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11992 9518 12020 10066
rect 12084 9654 12112 10066
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12360 9586 12388 10202
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11992 8634 12020 9454
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12360 8401 12388 9114
rect 12346 8392 12402 8401
rect 12164 8356 12216 8362
rect 12346 8327 12402 8336
rect 12164 8298 12216 8304
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11704 7346 11756 7352
rect 11808 7364 11928 7392
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11624 6168 11652 7210
rect 11716 6798 11744 7346
rect 11808 7206 11836 7364
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 6934 11928 7142
rect 11992 6934 12020 7482
rect 12070 7440 12126 7449
rect 12070 7375 12126 7384
rect 12084 7274 12112 7375
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6458 11744 6734
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11992 6254 12020 6326
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11796 6180 11848 6186
rect 11624 6140 11744 6168
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11624 5409 11652 5850
rect 11610 5400 11666 5409
rect 11520 5364 11572 5370
rect 11610 5335 11666 5344
rect 11520 5306 11572 5312
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11164 2961 11192 3878
rect 11348 3602 11376 3878
rect 11532 3670 11560 5306
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11348 3126 11376 3334
rect 11532 3126 11560 3606
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 2650 11100 2790
rect 11164 2650 11192 2887
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 11440 2446 11468 2994
rect 11624 2514 11652 4966
rect 11716 2990 11744 6140
rect 11796 6122 11848 6128
rect 11808 5914 11836 6122
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11808 5234 11836 5850
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11992 5030 12020 6190
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11808 4826 11836 4966
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11980 4616 12032 4622
rect 12084 4604 12112 5034
rect 12176 5012 12204 8298
rect 12452 8090 12480 10503
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7478 12296 7822
rect 12438 7712 12494 7721
rect 12438 7647 12494 7656
rect 12452 7546 12480 7647
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12268 7002 12296 7414
rect 12544 7392 12572 9687
rect 12452 7364 12572 7392
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 6798 12296 6938
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12268 5574 12296 6326
rect 12452 6254 12480 7364
rect 12530 7304 12586 7313
rect 12530 7239 12586 7248
rect 12544 7206 12572 7239
rect 12636 7206 12664 10950
rect 12728 7993 12756 12174
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12806 11112 12862 11121
rect 12806 11047 12862 11056
rect 12820 10742 12848 11047
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12820 10538 12848 10678
rect 13188 10656 13216 11766
rect 13280 11694 13308 12038
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10810 13400 11494
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13188 10628 13308 10656
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 13188 10266 13216 10474
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13280 10169 13308 10628
rect 13464 10470 13492 13903
rect 14924 13874 14976 13880
rect 15212 13546 15240 15127
rect 15382 13832 15438 13841
rect 15382 13767 15438 13776
rect 14752 13518 15240 13546
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13266 10160 13322 10169
rect 13266 10095 13322 10104
rect 13280 9602 13308 10095
rect 13464 10010 13492 10406
rect 13556 10266 13584 12582
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11286 13860 12174
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13832 10674 13860 11222
rect 13924 11218 13952 11630
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14016 11014 14044 11630
rect 14292 11354 14320 12242
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10674 14044 10950
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13832 10062 13860 10610
rect 14108 10198 14136 11154
rect 14384 10198 14412 11562
rect 14660 10713 14688 13330
rect 14752 12442 14780 13518
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15212 12889 15240 13398
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15198 12880 15254 12889
rect 15198 12815 15254 12824
rect 15016 12640 15068 12646
rect 15304 12617 15332 13194
rect 15016 12582 15068 12588
rect 15290 12608 15346 12617
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 15028 11558 15056 12582
rect 15290 12543 15346 12552
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 11694 15148 12038
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14646 10704 14702 10713
rect 14646 10639 14702 10648
rect 14660 10538 14688 10639
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14844 10441 14872 11494
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14830 10432 14886 10441
rect 14660 10390 14830 10418
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 13820 10056 13872 10062
rect 13464 9982 13584 10010
rect 13820 9998 13872 10004
rect 13452 9920 13504 9926
rect 13358 9888 13414 9897
rect 13452 9862 13504 9868
rect 13358 9823 13414 9832
rect 13188 9574 13308 9602
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12714 7984 12770 7993
rect 13188 7954 13216 9574
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 12714 7919 12770 7928
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12728 6458 12756 7210
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13176 6928 13228 6934
rect 12898 6896 12954 6905
rect 12898 6831 12900 6840
rect 12952 6831 12954 6840
rect 13174 6896 13176 6905
rect 13228 6896 13230 6905
rect 13174 6831 13230 6840
rect 12900 6802 12952 6808
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13188 5914 13216 6258
rect 13280 6225 13308 9386
rect 13372 8090 13400 9823
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6254 13400 7142
rect 13360 6248 13412 6254
rect 13266 6216 13322 6225
rect 13360 6190 13412 6196
rect 13266 6151 13322 6160
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 5166 12388 5510
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12452 5166 12480 5238
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12176 4984 12388 5012
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12032 4576 12112 4604
rect 11980 4558 12032 4564
rect 11992 4146 12020 4558
rect 12176 4282 12204 4762
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11796 3528 11848 3534
rect 11794 3496 11796 3505
rect 11848 3496 11850 3505
rect 11794 3431 11850 3440
rect 11992 2990 12020 3946
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 10336 1414 10456 1442
rect 10336 480 10364 1414
rect 11256 480 11284 2314
rect 11900 1222 11928 2790
rect 12360 2514 12388 4984
rect 12452 4826 12480 5102
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12440 4616 12492 4622
rect 12544 4604 12572 5578
rect 12636 4690 12664 5850
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 13188 4826 13216 5714
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12492 4576 12572 4604
rect 12440 4558 12492 4564
rect 12530 4176 12586 4185
rect 12728 4146 12756 4762
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12912 4282 12940 4694
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12530 4111 12532 4120
rect 12584 4111 12586 4120
rect 12716 4140 12768 4146
rect 12532 4082 12584 4088
rect 12716 4082 12768 4088
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 2650 12480 3878
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 13280 3738 13308 5646
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12728 2854 12756 3538
rect 13464 2990 13492 9862
rect 13556 9761 13584 9982
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 8945 13584 9046
rect 13648 8974 13676 9930
rect 13832 9654 13860 9998
rect 14108 9654 14136 10134
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14094 9480 14150 9489
rect 13636 8968 13688 8974
rect 13542 8936 13598 8945
rect 13820 8968 13872 8974
rect 13636 8910 13688 8916
rect 13818 8936 13820 8945
rect 13872 8936 13874 8945
rect 13542 8871 13598 8880
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8498 13584 8774
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13648 7698 13676 8910
rect 13818 8871 13874 8880
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 8294 13768 8434
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 7886 13768 8230
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13832 7818 13860 8502
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13924 7750 13952 9454
rect 14094 9415 14150 9424
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 7744 13964 7750
rect 13648 7670 13768 7698
rect 13912 7686 13964 7692
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 6866 13584 7278
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 6662 13584 6802
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 12176 480 12204 2382
rect 13188 1442 13216 2858
rect 13556 2854 13584 6151
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 3602 13676 6054
rect 13740 5234 13768 7670
rect 13924 5846 13952 7686
rect 14016 7546 14044 8366
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6254 14044 6666
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14108 5846 14136 9415
rect 14370 9208 14426 9217
rect 14370 9143 14372 9152
rect 14424 9143 14426 9152
rect 14372 9114 14424 9120
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14200 8090 14228 8774
rect 14292 8430 14320 8774
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14292 6769 14320 6870
rect 14278 6760 14334 6769
rect 14278 6695 14334 6704
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5914 14228 6054
rect 14292 5914 14320 6695
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6254 14412 6598
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5370 13860 5578
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 13910 5400 13966 5409
rect 13820 5364 13872 5370
rect 13910 5335 13966 5344
rect 13820 5306 13872 5312
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13924 4758 13952 5335
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 13912 4752 13964 4758
rect 13726 4720 13782 4729
rect 13912 4694 13964 4700
rect 13726 4655 13782 4664
rect 13740 3738 13768 4655
rect 14016 4622 14044 5034
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14016 4214 14044 4558
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13832 3398 13860 4014
rect 14016 3602 14044 4150
rect 14292 3602 14320 5471
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 14108 3126 14136 3470
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 14476 2514 14504 9862
rect 14568 9722 14596 10066
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14568 9178 14596 9658
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14660 6202 14688 10390
rect 14830 10367 14886 10376
rect 14830 10296 14886 10305
rect 14830 10231 14886 10240
rect 14844 9450 14872 10231
rect 14936 9994 14964 10542
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 15028 9450 15056 11222
rect 15120 11218 15148 11494
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15120 10062 15148 11154
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15212 9178 15240 12378
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 9722 15332 10950
rect 15396 10577 15424 13767
rect 15580 12170 15608 15399
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15474 11656 15530 11665
rect 15474 11591 15530 11600
rect 15382 10568 15438 10577
rect 15382 10503 15438 10512
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 9466 15332 9658
rect 15304 9438 15424 9466
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14844 8362 14872 8910
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14936 7206 14964 8910
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 7886 15240 8230
rect 15304 7993 15332 9318
rect 15396 9042 15424 9438
rect 15488 9217 15516 11591
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 10674 15608 11494
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15672 10554 15700 16079
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 16132 12322 16160 16487
rect 16302 15872 16358 15881
rect 16302 15807 16358 15816
rect 16132 12294 16252 12322
rect 16118 12200 16174 12209
rect 16118 12135 16174 12144
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16132 11898 16160 12135
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 15752 10668 15804 10674
rect 15844 10668 15896 10674
rect 15804 10628 15844 10656
rect 15752 10610 15804 10616
rect 16028 10668 16080 10674
rect 15844 10610 15896 10616
rect 15948 10628 16028 10656
rect 15580 10526 15700 10554
rect 15474 9208 15530 9217
rect 15474 9143 15530 9152
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15396 8838 15424 8978
rect 15384 8832 15436 8838
rect 15580 8786 15608 10526
rect 15948 10520 15976 10628
rect 16028 10610 16080 10616
rect 15764 10492 15976 10520
rect 15764 10180 15792 10492
rect 16132 10266 16160 10678
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 15672 10152 15792 10180
rect 15672 9994 15700 10152
rect 16120 10056 16172 10062
rect 16224 10033 16252 12294
rect 16316 11676 16344 15807
rect 16394 14920 16450 14929
rect 16394 14855 16450 14864
rect 16408 11812 16436 14855
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 14074 17632 14282
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16500 11880 16528 12922
rect 16500 11852 16712 11880
rect 16408 11784 16528 11812
rect 16316 11648 16436 11676
rect 16408 11257 16436 11648
rect 16394 11248 16450 11257
rect 16394 11183 16450 11192
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10606 16344 10950
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16302 10160 16358 10169
rect 16302 10095 16304 10104
rect 16356 10095 16358 10104
rect 16304 10066 16356 10072
rect 16120 9998 16172 10004
rect 16210 10024 16266 10033
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15672 9518 15700 9930
rect 16132 9874 16160 9998
rect 16210 9959 16266 9968
rect 16132 9846 16252 9874
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 16040 9042 16068 9590
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15384 8774 15436 8780
rect 15396 8498 15424 8774
rect 15488 8758 15608 8786
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15382 8392 15438 8401
rect 15382 8327 15438 8336
rect 15290 7984 15346 7993
rect 15290 7919 15346 7928
rect 15200 7880 15252 7886
rect 15014 7848 15070 7857
rect 15200 7822 15252 7828
rect 15014 7783 15016 7792
rect 15068 7783 15070 7792
rect 15016 7754 15068 7760
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 15028 7206 15056 7414
rect 15120 7410 15148 7686
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15106 7304 15162 7313
rect 15212 7274 15240 7822
rect 15106 7239 15162 7248
rect 15200 7268 15252 7274
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14568 6174 14688 6202
rect 14568 5273 14596 6174
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14554 5264 14610 5273
rect 14554 5199 14610 5208
rect 14568 4078 14596 5199
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14660 2990 14688 6054
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14752 4690 14780 5850
rect 14844 5710 14872 6734
rect 15028 6066 15056 7142
rect 15120 6390 15148 7239
rect 15200 7210 15252 7216
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15198 6760 15254 6769
rect 15198 6695 15254 6704
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14936 6038 15056 6066
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14844 5234 14872 5646
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14936 3641 14964 6038
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15028 5166 15056 5510
rect 15212 5370 15240 6695
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4282 15240 4422
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 14922 3632 14978 3641
rect 14922 3567 14978 3576
rect 15304 2990 15332 7142
rect 15396 6662 15424 8327
rect 15488 6730 15516 8758
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15580 8022 15608 8570
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7410 15608 7754
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15568 7200 15620 7206
rect 15566 7168 15568 7177
rect 15620 7168 15622 7177
rect 15566 7103 15622 7112
rect 15672 7002 15700 8230
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15568 6860 15620 6866
rect 15752 6860 15804 6866
rect 15568 6802 15620 6808
rect 15672 6820 15752 6848
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15580 6390 15608 6802
rect 15568 6384 15620 6390
rect 15382 6352 15438 6361
rect 15568 6326 15620 6332
rect 15382 6287 15438 6296
rect 15476 6316 15528 6322
rect 15396 4826 15424 6287
rect 15476 6258 15528 6264
rect 15488 5846 15516 6258
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15580 5574 15608 6326
rect 15672 6322 15700 6820
rect 15752 6802 15804 6808
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 5914 15700 6258
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15842 5128 15898 5137
rect 15842 5063 15898 5072
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15764 4758 15792 4966
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15856 4622 15884 5063
rect 16132 4826 16160 9658
rect 16224 9654 16252 9846
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16224 7818 16252 8366
rect 16316 7886 16344 10066
rect 16408 9586 16436 11183
rect 16500 10010 16528 11784
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16592 10538 16620 11698
rect 16684 11558 16712 11852
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16684 10577 16712 11494
rect 16670 10568 16726 10577
rect 16580 10532 16632 10538
rect 16670 10503 16726 10512
rect 16580 10474 16632 10480
rect 16500 9982 16620 10010
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16394 8936 16450 8945
rect 16394 8871 16450 8880
rect 16408 8430 16436 8871
rect 16500 8673 16528 9862
rect 16592 9722 16620 9982
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16486 8664 16542 8673
rect 16486 8599 16542 8608
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16684 8242 16712 10503
rect 16500 8214 16712 8242
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16500 7206 16528 8214
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 7342 16712 7890
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16302 7032 16358 7041
rect 16302 6967 16358 6976
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15566 4448 15622 4457
rect 15396 4185 15424 4422
rect 15566 4383 15622 4392
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 15580 4078 15608 4383
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 16132 4078 16160 4626
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16224 3890 16252 6802
rect 16316 3942 16344 6967
rect 16592 6905 16620 7210
rect 16578 6896 16634 6905
rect 16578 6831 16634 6840
rect 16486 6352 16542 6361
rect 16486 6287 16542 6296
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16408 5370 16436 5782
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16132 3862 16252 3890
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16132 3738 16160 3862
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16224 3194 16252 3674
rect 16500 3482 16528 6287
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 5370 16712 6054
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16684 4078 16712 5170
rect 16776 5114 16804 13942
rect 17880 13870 17908 16759
rect 18234 16520 18290 17000
rect 18248 14074 18276 16520
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 17052 11558 17080 12650
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16854 11248 16910 11257
rect 16854 11183 16910 11192
rect 16868 10713 16896 11183
rect 16854 10704 16910 10713
rect 16854 10639 16910 10648
rect 16868 7818 16896 10639
rect 17144 8922 17172 11630
rect 17236 11286 17264 11698
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9722 17264 10066
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17328 9178 17356 9998
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17144 8894 17356 8922
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 16960 8022 16988 8774
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 7449 16896 7754
rect 16854 7440 16910 7449
rect 16854 7375 16910 7384
rect 16960 7188 16988 7822
rect 16868 7160 16988 7188
rect 16868 5234 16896 7160
rect 17144 6730 17172 8774
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17236 7886 17264 8298
rect 17328 7954 17356 8894
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17236 7410 17264 7822
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17236 7002 17264 7346
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17420 6746 17448 13806
rect 17866 13288 17922 13297
rect 17866 13223 17922 13232
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 8786 17540 11494
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10538 17632 10950
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17604 9586 17632 10474
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10062 17724 10406
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17604 8974 17632 9522
rect 17696 9110 17724 9862
rect 17788 9518 17816 12174
rect 17880 10266 17908 13223
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17866 10160 17922 10169
rect 17866 10095 17922 10104
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9178 17816 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17512 8758 17632 8786
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17512 6934 17540 8366
rect 17604 7206 17632 8758
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 7886 17724 8230
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17880 7290 17908 10095
rect 17788 7262 17908 7290
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 17236 6718 17448 6746
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17144 6254 17172 6666
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16960 5234 16988 5510
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16776 5086 16988 5114
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4826 16804 4966
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16854 4720 16910 4729
rect 16854 4655 16910 4664
rect 16868 4282 16896 4655
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16960 4146 16988 5086
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16500 3466 16620 3482
rect 16500 3460 16632 3466
rect 16500 3454 16580 3460
rect 16580 3402 16632 3408
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 13096 1414 13216 1442
rect 13096 480 13124 1414
rect 13924 480 13952 2382
rect 14844 480 14872 2858
rect 15672 1442 15700 2858
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16224 1873 16252 3130
rect 16304 3120 16356 3126
rect 16302 3088 16304 3097
rect 16356 3088 16358 3097
rect 16302 3023 16358 3032
rect 16316 2990 16344 3023
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16500 2496 16528 3334
rect 16500 2468 16620 2496
rect 16486 2408 16542 2417
rect 16486 2343 16488 2352
rect 16540 2343 16542 2352
rect 16488 2314 16540 2320
rect 16500 2145 16528 2314
rect 16486 2136 16542 2145
rect 16486 2071 16542 2080
rect 16592 1986 16620 2468
rect 16500 1958 16620 1986
rect 16210 1864 16266 1873
rect 16210 1799 16266 1808
rect 15672 1414 15792 1442
rect 15764 480 15792 1414
rect 3330 439 3386 448
rect 3146 232 3202 241
rect 3146 167 3202 176
rect 3974 0 4030 480
rect 4894 0 4950 480
rect 5814 0 5870 480
rect 6734 0 6790 480
rect 7562 0 7618 480
rect 8482 0 8538 480
rect 9402 0 9458 480
rect 10322 0 10378 480
rect 11242 0 11298 480
rect 12162 0 12218 480
rect 13082 0 13138 480
rect 13910 0 13966 480
rect 14830 0 14886 480
rect 15750 0 15806 480
rect 16500 241 16528 1958
rect 16684 480 16712 3606
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16776 1465 16804 2858
rect 16868 2825 16896 3975
rect 17236 3670 17264 6718
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 5914 17448 6598
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5840 17368 5846
rect 17314 5808 17316 5817
rect 17368 5808 17370 5817
rect 17314 5743 17370 5752
rect 17328 5166 17356 5743
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17406 4040 17462 4049
rect 17512 4010 17540 6734
rect 17604 4434 17632 7142
rect 17788 7002 17816 7262
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17776 6112 17828 6118
rect 17880 6089 17908 7142
rect 17972 6866 18000 11630
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18050 11112 18106 11121
rect 18050 11047 18106 11056
rect 18064 10606 18092 11047
rect 18142 10976 18198 10985
rect 18142 10911 18198 10920
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18156 10305 18184 10911
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18142 10296 18198 10305
rect 18142 10231 18198 10240
rect 18050 10024 18106 10033
rect 18050 9959 18052 9968
rect 18104 9959 18106 9968
rect 18052 9930 18104 9936
rect 18050 8120 18106 8129
rect 18050 8055 18106 8064
rect 18064 7342 18092 8055
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17776 6054 17828 6060
rect 17866 6080 17922 6089
rect 17696 5710 17724 6054
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17696 4622 17724 5646
rect 17788 5409 17816 6054
rect 17866 6015 17922 6024
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17972 5681 18000 5714
rect 17958 5672 18014 5681
rect 17958 5607 18014 5616
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17774 5400 17830 5409
rect 17774 5335 17830 5344
rect 17880 5137 17908 5510
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 18156 4826 18184 10231
rect 18236 9376 18288 9382
rect 18234 9344 18236 9353
rect 18288 9344 18290 9353
rect 18234 9279 18290 9288
rect 18340 8945 18368 10406
rect 18326 8936 18382 8945
rect 18326 8871 18382 8880
rect 18432 8401 18460 11494
rect 18970 9616 19026 9625
rect 18970 9551 18972 9560
rect 19024 9551 19026 9560
rect 18972 9522 19024 9528
rect 18418 8392 18474 8401
rect 18418 8327 18474 8336
rect 18418 5672 18474 5681
rect 18418 5607 18474 5616
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17604 4406 17724 4434
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17406 3975 17462 3984
rect 17500 4004 17552 4010
rect 17420 3942 17448 3975
rect 17500 3946 17552 3952
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17236 2990 17264 3606
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 16854 2816 16910 2825
rect 16854 2751 16910 2760
rect 16868 2650 16896 2751
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17040 2440 17092 2446
rect 17236 2417 17264 2926
rect 17040 2382 17092 2388
rect 17222 2408 17278 2417
rect 16762 1456 16818 1465
rect 16762 1391 16818 1400
rect 17052 1193 17080 2382
rect 17222 2343 17278 2352
rect 17038 1184 17094 1193
rect 17038 1119 17094 1128
rect 17604 480 17632 4082
rect 17696 4078 17724 4406
rect 17788 4214 17816 4626
rect 18248 4457 18276 4966
rect 18234 4448 18290 4457
rect 18234 4383 18290 4392
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17788 3505 17816 4150
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3777 18276 3878
rect 18234 3768 18290 3777
rect 18234 3703 18290 3712
rect 18052 3528 18104 3534
rect 17774 3496 17830 3505
rect 18052 3470 18104 3476
rect 17774 3431 17830 3440
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17788 513 17816 2382
rect 18064 785 18092 3470
rect 18432 3194 18460 5607
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18050 776 18106 785
rect 18050 711 18106 720
rect 17774 504 17830 513
rect 16486 232 16542 241
rect 16486 167 16542 176
rect 16670 0 16726 480
rect 17590 0 17646 480
rect 18524 480 18552 4558
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19444 480 19472 2858
rect 17774 439 17830 448
rect 18510 0 18566 480
rect 19430 0 19486 480
<< via2 >>
rect 3330 16768 3386 16824
rect 3790 16496 3846 16552
rect 3422 16088 3478 16144
rect 3238 15408 3294 15464
rect 2870 15136 2926 15192
rect 2042 14728 2098 14784
rect 2778 14492 2780 14512
rect 2780 14492 2832 14512
rect 2832 14492 2834 14512
rect 2778 14456 2834 14492
rect 2778 14048 2834 14104
rect 1858 13812 1860 13832
rect 1860 13812 1912 13832
rect 1912 13812 1914 13832
rect 1858 13776 1914 13812
rect 3330 14320 3386 14376
rect 4066 15816 4122 15872
rect 17866 16768 17922 16824
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3054 13812 3056 13832
rect 3056 13812 3108 13832
rect 3108 13812 3110 13832
rect 3054 13776 3110 13812
rect 3606 13812 3608 13832
rect 3608 13812 3660 13832
rect 3660 13812 3662 13832
rect 3606 13776 3662 13812
rect 3330 13388 3386 13424
rect 3330 13368 3332 13388
rect 3332 13368 3384 13388
rect 3384 13368 3386 13388
rect 1214 8608 1270 8664
rect 1306 4256 1362 4312
rect 1674 8356 1730 8392
rect 1674 8336 1676 8356
rect 1676 8336 1728 8356
rect 1728 8336 1730 8356
rect 1398 3848 1454 3904
rect 1582 3576 1638 3632
rect 1214 3440 1270 3496
rect 1398 2624 1454 2680
rect 2134 8064 2190 8120
rect 2134 7656 2190 7712
rect 2042 6976 2098 7032
rect 2962 13096 3018 13152
rect 2686 10240 2742 10296
rect 2870 11328 2926 11384
rect 2778 9424 2834 9480
rect 2778 8336 2834 8392
rect 2686 7792 2742 7848
rect 2594 7248 2650 7304
rect 2318 6024 2374 6080
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3790 12688 3846 12744
rect 3330 12416 3386 12472
rect 3330 12144 3386 12200
rect 3146 11736 3202 11792
rect 3422 11056 3478 11112
rect 2778 5752 2834 5808
rect 2962 6568 3018 6624
rect 2870 3168 2926 3224
rect 3330 7248 3386 7304
rect 3238 5888 3294 5944
rect 3330 2644 3386 2680
rect 3330 2624 3332 2644
rect 3332 2624 3384 2644
rect 3384 2624 3386 2644
rect 3698 12008 3754 12064
rect 3698 9288 3754 9344
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 4066 10648 4122 10704
rect 4342 10376 4398 10432
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4342 9696 4398 9752
rect 3974 9560 4030 9616
rect 4158 9288 4214 9344
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 4066 8336 4122 8392
rect 4342 9424 4398 9480
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3790 6296 3846 6352
rect 3974 5616 4030 5672
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3882 5108 3884 5128
rect 3884 5108 3936 5128
rect 3936 5108 3938 5128
rect 3882 5072 3938 5108
rect 4066 4936 4122 4992
rect 3882 4528 3938 4584
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3606 2508 3662 2544
rect 3606 2488 3608 2508
rect 3608 2488 3660 2508
rect 3660 2488 3662 2508
rect 3698 2216 3754 2272
rect 3422 1808 3478 1864
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 4066 2896 4122 2952
rect 4710 8472 4766 8528
rect 4526 6568 4582 6624
rect 4434 5480 4490 5536
rect 4710 6296 4766 6352
rect 4618 5344 4674 5400
rect 4986 10240 5042 10296
rect 4894 7384 4950 7440
rect 4894 5072 4950 5128
rect 4894 4528 4950 4584
rect 4618 2488 4674 2544
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 3698 856 3754 912
rect 3330 448 3386 504
rect 4066 1164 4068 1184
rect 4068 1164 4120 1184
rect 4120 1164 4122 1184
rect 4066 1128 4122 1164
rect 5078 7520 5134 7576
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 13450 13912 13506 13968
rect 16118 16496 16174 16552
rect 15658 16088 15714 16144
rect 15566 15408 15622 15464
rect 15198 15136 15254 15192
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 5446 6160 5502 6216
rect 5354 4800 5410 4856
rect 5262 2896 5318 2952
rect 5814 6432 5870 6488
rect 5998 7964 6000 7984
rect 6000 7964 6052 7984
rect 6052 7964 6054 7984
rect 5998 7928 6054 7964
rect 5906 5208 5962 5264
rect 5722 4256 5778 4312
rect 6090 6976 6146 7032
rect 6274 9968 6330 10024
rect 6366 9288 6422 9344
rect 6182 6840 6238 6896
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 7654 12008 7710 12064
rect 7102 10104 7158 10160
rect 6826 9832 6882 9888
rect 7194 9696 7250 9752
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7378 9152 7434 9208
rect 6642 8744 6698 8800
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6642 8064 6698 8120
rect 7194 7384 7250 7440
rect 6090 5208 6146 5264
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6642 5344 6698 5400
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 7194 4664 7250 4720
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 7838 10512 7894 10568
rect 7930 8472 7986 8528
rect 7930 7948 7986 7984
rect 7930 7928 7932 7948
rect 7932 7928 7984 7948
rect 7984 7928 7986 7948
rect 7654 7520 7710 7576
rect 7470 6432 7526 6488
rect 4986 1536 5042 1592
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 8482 12144 8538 12200
rect 8390 9832 8446 9888
rect 8574 7384 8630 7440
rect 8390 6160 8446 6216
rect 8666 7248 8722 7304
rect 9034 9288 9090 9344
rect 8942 8880 8998 8936
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9862 11192 9918 11248
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9770 10104 9826 10160
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9402 9016 9458 9072
rect 9126 8744 9182 8800
rect 8942 7792 8998 7848
rect 8574 6160 8630 6216
rect 8206 4800 8262 4856
rect 8390 5208 8446 5264
rect 8758 5908 8814 5944
rect 8758 5888 8760 5908
rect 8760 5888 8812 5908
rect 8812 5888 8814 5908
rect 8758 5752 8814 5808
rect 8574 5480 8630 5536
rect 8574 5344 8630 5400
rect 8942 6860 8998 6896
rect 8942 6840 8944 6860
rect 8944 6840 8996 6860
rect 8996 6840 8998 6860
rect 8850 5108 8852 5128
rect 8852 5108 8904 5128
rect 8904 5108 8906 5128
rect 8850 5072 8906 5108
rect 8758 4256 8814 4312
rect 9310 6568 9366 6624
rect 9402 5208 9458 5264
rect 9034 4528 9090 4584
rect 9218 4528 9274 4584
rect 9034 2508 9090 2544
rect 9034 2488 9036 2508
rect 9036 2488 9088 2508
rect 9088 2488 9090 2508
rect 10506 9560 10562 9616
rect 10414 9152 10470 9208
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9862 6860 9918 6896
rect 9862 6840 9864 6860
rect 9864 6840 9916 6860
rect 9916 6840 9918 6860
rect 9678 6704 9734 6760
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9586 2896 9642 2952
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 11058 7812 11114 7848
rect 11058 7792 11060 7812
rect 11060 7792 11112 7812
rect 11112 7792 11114 7812
rect 10966 7656 11022 7712
rect 10506 5480 10562 5536
rect 10690 5072 10746 5128
rect 10690 4392 10746 4448
rect 10322 3440 10378 3496
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 11334 9152 11390 9208
rect 11426 5888 11482 5944
rect 11610 9324 11612 9344
rect 11612 9324 11664 9344
rect 11664 9324 11666 9344
rect 11610 9288 11666 9324
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12438 10512 12494 10568
rect 12346 8336 12402 8392
rect 12070 7384 12126 7440
rect 11610 5344 11666 5400
rect 11150 2896 11206 2952
rect 12530 9696 12586 9752
rect 12438 7656 12494 7712
rect 12530 7248 12586 7304
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12806 11056 12862 11112
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 15382 13776 15438 13832
rect 13266 10104 13322 10160
rect 15198 12824 15254 12880
rect 15290 12552 15346 12608
rect 14646 10648 14702 10704
rect 13358 9832 13414 9888
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12714 7928 12770 7984
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12898 6860 12954 6896
rect 12898 6840 12900 6860
rect 12900 6840 12952 6860
rect 12952 6840 12954 6860
rect 13174 6876 13176 6896
rect 13176 6876 13228 6896
rect 13228 6876 13230 6896
rect 13174 6840 13230 6876
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 13266 6160 13322 6216
rect 11794 3476 11796 3496
rect 11796 3476 11848 3496
rect 11848 3476 11850 3496
rect 11794 3440 11850 3476
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12530 4140 12586 4176
rect 12530 4120 12532 4140
rect 12532 4120 12584 4140
rect 12584 4120 12586 4140
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 13542 9696 13598 9752
rect 13542 8880 13598 8936
rect 13818 8916 13820 8936
rect 13820 8916 13872 8936
rect 13872 8916 13874 8936
rect 13818 8880 13874 8916
rect 14094 9424 14150 9480
rect 13542 6160 13598 6216
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 14370 9172 14426 9208
rect 14370 9152 14372 9172
rect 14372 9152 14424 9172
rect 14424 9152 14426 9172
rect 14278 6704 14334 6760
rect 14278 5480 14334 5536
rect 13910 5344 13966 5400
rect 13726 4664 13782 4720
rect 14830 10376 14886 10432
rect 14830 10240 14886 10296
rect 15474 11600 15530 11656
rect 15382 10512 15438 10568
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 16302 15816 16358 15872
rect 16118 12144 16174 12200
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15474 9152 15530 9208
rect 16394 14864 16450 14920
rect 16394 11192 16450 11248
rect 16302 10124 16358 10160
rect 16302 10104 16304 10124
rect 16304 10104 16356 10124
rect 16356 10104 16358 10124
rect 16210 9968 16266 10024
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15382 8336 15438 8392
rect 15290 7928 15346 7984
rect 15014 7812 15070 7848
rect 15014 7792 15016 7812
rect 15016 7792 15068 7812
rect 15068 7792 15070 7812
rect 15106 7248 15162 7304
rect 14554 5208 14610 5264
rect 15198 6704 15254 6760
rect 14922 3576 14978 3632
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15566 7148 15568 7168
rect 15568 7148 15620 7168
rect 15620 7148 15622 7168
rect 15566 7112 15622 7148
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15382 6296 15438 6352
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15842 5072 15898 5128
rect 16670 10512 16726 10568
rect 16394 8880 16450 8936
rect 16486 8608 16542 8664
rect 16302 6976 16358 7032
rect 15566 4392 15622 4448
rect 15382 4120 15438 4176
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 16578 6840 16634 6896
rect 16486 6296 16542 6352
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 16854 11192 16910 11248
rect 16854 10648 16910 10704
rect 16854 7384 16910 7440
rect 17866 13232 17922 13288
rect 17866 10104 17922 10160
rect 16854 4664 16910 4720
rect 16854 3984 16910 4040
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16302 3068 16304 3088
rect 16304 3068 16356 3088
rect 16356 3068 16358 3088
rect 16302 3032 16358 3068
rect 16486 2372 16542 2408
rect 16486 2352 16488 2372
rect 16488 2352 16540 2372
rect 16540 2352 16542 2372
rect 16486 2080 16542 2136
rect 16210 1808 16266 1864
rect 3146 176 3202 232
rect 17314 5788 17316 5808
rect 17316 5788 17368 5808
rect 17368 5788 17370 5808
rect 17314 5752 17370 5788
rect 17406 3984 17462 4040
rect 18050 11056 18106 11112
rect 18142 10920 18198 10976
rect 18142 10240 18198 10296
rect 18050 9988 18106 10024
rect 18050 9968 18052 9988
rect 18052 9968 18104 9988
rect 18104 9968 18106 9988
rect 18050 8064 18106 8120
rect 17866 6024 17922 6080
rect 17958 5616 18014 5672
rect 17774 5344 17830 5400
rect 17866 5072 17922 5128
rect 18234 9324 18236 9344
rect 18236 9324 18288 9344
rect 18288 9324 18290 9344
rect 18234 9288 18290 9324
rect 18326 8880 18382 8936
rect 18970 9580 19026 9616
rect 18970 9560 18972 9580
rect 18972 9560 19024 9580
rect 19024 9560 19026 9580
rect 18418 8336 18474 8392
rect 18418 5616 18474 5672
rect 16854 2760 16910 2816
rect 16762 1400 16818 1456
rect 17222 2352 17278 2408
rect 17038 1128 17094 1184
rect 18234 4392 18290 4448
rect 18234 3712 18290 3768
rect 17774 3440 17830 3496
rect 18050 720 18106 776
rect 16486 176 16542 232
rect 17774 448 17830 504
<< metal3 >>
rect 0 16826 480 16856
rect 3325 16826 3391 16829
rect 0 16824 3391 16826
rect 0 16768 3330 16824
rect 3386 16768 3391 16824
rect 0 16766 3391 16768
rect 0 16736 480 16766
rect 3325 16763 3391 16766
rect 17861 16826 17927 16829
rect 19520 16826 20000 16856
rect 17861 16824 20000 16826
rect 17861 16768 17866 16824
rect 17922 16768 20000 16824
rect 17861 16766 20000 16768
rect 17861 16763 17927 16766
rect 19520 16736 20000 16766
rect 0 16554 480 16584
rect 3785 16554 3851 16557
rect 0 16552 3851 16554
rect 0 16496 3790 16552
rect 3846 16496 3851 16552
rect 0 16494 3851 16496
rect 0 16464 480 16494
rect 3785 16491 3851 16494
rect 16113 16554 16179 16557
rect 19520 16554 20000 16584
rect 16113 16552 20000 16554
rect 16113 16496 16118 16552
rect 16174 16496 20000 16552
rect 16113 16494 20000 16496
rect 16113 16491 16179 16494
rect 19520 16464 20000 16494
rect 0 16146 480 16176
rect 3417 16146 3483 16149
rect 0 16144 3483 16146
rect 0 16088 3422 16144
rect 3478 16088 3483 16144
rect 0 16086 3483 16088
rect 0 16056 480 16086
rect 3417 16083 3483 16086
rect 15653 16146 15719 16149
rect 19520 16146 20000 16176
rect 15653 16144 20000 16146
rect 15653 16088 15658 16144
rect 15714 16088 20000 16144
rect 15653 16086 20000 16088
rect 15653 16083 15719 16086
rect 19520 16056 20000 16086
rect 0 15874 480 15904
rect 4061 15874 4127 15877
rect 0 15872 4127 15874
rect 0 15816 4066 15872
rect 4122 15816 4127 15872
rect 0 15814 4127 15816
rect 0 15784 480 15814
rect 4061 15811 4127 15814
rect 16297 15874 16363 15877
rect 19520 15874 20000 15904
rect 16297 15872 20000 15874
rect 16297 15816 16302 15872
rect 16358 15816 20000 15872
rect 16297 15814 20000 15816
rect 16297 15811 16363 15814
rect 19520 15784 20000 15814
rect 0 15466 480 15496
rect 3233 15466 3299 15469
rect 0 15464 3299 15466
rect 0 15408 3238 15464
rect 3294 15408 3299 15464
rect 0 15406 3299 15408
rect 0 15376 480 15406
rect 3233 15403 3299 15406
rect 15561 15466 15627 15469
rect 19520 15466 20000 15496
rect 15561 15464 20000 15466
rect 15561 15408 15566 15464
rect 15622 15408 20000 15464
rect 15561 15406 20000 15408
rect 15561 15403 15627 15406
rect 19520 15376 20000 15406
rect 0 15194 480 15224
rect 2865 15194 2931 15197
rect 0 15192 2931 15194
rect 0 15136 2870 15192
rect 2926 15136 2931 15192
rect 0 15134 2931 15136
rect 0 15104 480 15134
rect 2865 15131 2931 15134
rect 15193 15194 15259 15197
rect 19520 15194 20000 15224
rect 15193 15192 20000 15194
rect 15193 15136 15198 15192
rect 15254 15136 20000 15192
rect 15193 15134 20000 15136
rect 15193 15131 15259 15134
rect 19520 15104 20000 15134
rect 16389 14922 16455 14925
rect 19520 14922 20000 14952
rect 16389 14920 20000 14922
rect 16389 14864 16394 14920
rect 16450 14864 20000 14920
rect 16389 14862 20000 14864
rect 16389 14859 16455 14862
rect 19520 14832 20000 14862
rect 0 14786 480 14816
rect 2037 14786 2103 14789
rect 0 14784 2103 14786
rect 0 14728 2042 14784
rect 2098 14728 2103 14784
rect 0 14726 2103 14728
rect 0 14696 480 14726
rect 2037 14723 2103 14726
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 0 14514 480 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 480 14454
rect 2773 14451 2839 14454
rect 16246 14452 16252 14516
rect 16316 14514 16322 14516
rect 19520 14514 20000 14544
rect 16316 14454 20000 14514
rect 16316 14452 16322 14454
rect 19520 14424 20000 14454
rect 3325 14380 3391 14381
rect 3325 14378 3372 14380
rect 3280 14376 3372 14378
rect 3280 14320 3330 14376
rect 3280 14318 3372 14320
rect 3325 14316 3372 14318
rect 3436 14316 3442 14380
rect 3325 14315 3391 14316
rect 19520 14242 20000 14272
rect 16208 14182 20000 14242
rect 3909 14176 4229 14177
rect 0 14106 480 14136
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 14111 16090 14112
rect 2773 14106 2839 14109
rect 0 14104 2839 14106
rect 0 14048 2778 14104
rect 2834 14048 2839 14104
rect 0 14046 2839 14048
rect 0 14016 480 14046
rect 2773 14043 2839 14046
rect 13445 13970 13511 13973
rect 16208 13970 16268 14182
rect 19520 14152 20000 14182
rect 13445 13968 16268 13970
rect 13445 13912 13450 13968
rect 13506 13912 16268 13968
rect 13445 13910 16268 13912
rect 13445 13907 13511 13910
rect 0 13834 480 13864
rect 1853 13834 1919 13837
rect 0 13832 1919 13834
rect 0 13776 1858 13832
rect 1914 13776 1919 13832
rect 0 13774 1919 13776
rect 0 13744 480 13774
rect 1853 13771 1919 13774
rect 3049 13834 3115 13837
rect 3182 13834 3188 13836
rect 3049 13832 3188 13834
rect 3049 13776 3054 13832
rect 3110 13776 3188 13832
rect 3049 13774 3188 13776
rect 3049 13771 3115 13774
rect 3182 13772 3188 13774
rect 3252 13772 3258 13836
rect 3601 13834 3667 13837
rect 3734 13834 3740 13836
rect 3601 13832 3740 13834
rect 3601 13776 3606 13832
rect 3662 13776 3740 13832
rect 3601 13774 3740 13776
rect 3601 13771 3667 13774
rect 3734 13772 3740 13774
rect 3804 13772 3810 13836
rect 15377 13834 15443 13837
rect 19520 13834 20000 13864
rect 15377 13832 20000 13834
rect 15377 13776 15382 13832
rect 15438 13776 20000 13832
rect 15377 13774 20000 13776
rect 15377 13771 15443 13774
rect 19520 13744 20000 13774
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 15142 13500 15148 13564
rect 15212 13562 15218 13564
rect 19520 13562 20000 13592
rect 15212 13502 20000 13562
rect 15212 13500 15218 13502
rect 19520 13472 20000 13502
rect 0 13426 480 13456
rect 3325 13426 3391 13429
rect 0 13424 3391 13426
rect 0 13368 3330 13424
rect 3386 13368 3391 13424
rect 0 13366 3391 13368
rect 0 13336 480 13366
rect 3325 13363 3391 13366
rect 17861 13290 17927 13293
rect 19520 13290 20000 13320
rect 17861 13288 20000 13290
rect 17861 13232 17866 13288
rect 17922 13232 20000 13288
rect 17861 13230 20000 13232
rect 17861 13227 17927 13230
rect 19520 13200 20000 13230
rect 0 13154 480 13184
rect 2957 13154 3023 13157
rect 0 13152 3023 13154
rect 0 13096 2962 13152
rect 3018 13096 3023 13152
rect 0 13094 3023 13096
rect 0 13064 480 13094
rect 2957 13091 3023 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 15193 12882 15259 12885
rect 19520 12882 20000 12912
rect 15193 12880 20000 12882
rect 15193 12824 15198 12880
rect 15254 12824 20000 12880
rect 15193 12822 20000 12824
rect 15193 12819 15259 12822
rect 19520 12792 20000 12822
rect 0 12746 480 12776
rect 3785 12746 3851 12749
rect 0 12744 3851 12746
rect 0 12688 3790 12744
rect 3846 12688 3851 12744
rect 0 12686 3851 12688
rect 0 12656 480 12686
rect 3785 12683 3851 12686
rect 15285 12610 15351 12613
rect 19520 12610 20000 12640
rect 15285 12608 20000 12610
rect 15285 12552 15290 12608
rect 15346 12552 20000 12608
rect 15285 12550 20000 12552
rect 15285 12547 15351 12550
rect 6874 12544 7194 12545
rect 0 12474 480 12504
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 19520 12520 20000 12550
rect 12805 12479 13125 12480
rect 3325 12474 3391 12477
rect 0 12472 3391 12474
rect 0 12416 3330 12472
rect 3386 12416 3391 12472
rect 0 12414 3391 12416
rect 0 12384 480 12414
rect 3325 12411 3391 12414
rect 3325 12202 3391 12205
rect 8477 12202 8543 12205
rect 3325 12200 8543 12202
rect 3325 12144 3330 12200
rect 3386 12144 8482 12200
rect 8538 12144 8543 12200
rect 3325 12142 8543 12144
rect 3325 12139 3391 12142
rect 8477 12139 8543 12142
rect 16113 12202 16179 12205
rect 19520 12202 20000 12232
rect 16113 12200 20000 12202
rect 16113 12144 16118 12200
rect 16174 12144 20000 12200
rect 16113 12142 20000 12144
rect 16113 12139 16179 12142
rect 19520 12112 20000 12142
rect 0 12066 480 12096
rect 3693 12066 3759 12069
rect 7649 12068 7715 12069
rect 0 12064 3759 12066
rect 0 12008 3698 12064
rect 3754 12008 3759 12064
rect 0 12006 3759 12008
rect 0 11976 480 12006
rect 3693 12003 3759 12006
rect 7598 12004 7604 12068
rect 7668 12066 7715 12068
rect 7668 12064 7760 12066
rect 7710 12008 7760 12064
rect 7668 12006 7760 12008
rect 7668 12004 7715 12006
rect 7649 12003 7715 12004
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 19520 11930 20000 11960
rect 16254 11870 20000 11930
rect 0 11794 480 11824
rect 3141 11794 3207 11797
rect 0 11792 3207 11794
rect 0 11736 3146 11792
rect 3202 11736 3207 11792
rect 0 11734 3207 11736
rect 0 11704 480 11734
rect 3141 11731 3207 11734
rect 15510 11732 15516 11796
rect 15580 11794 15586 11796
rect 16254 11794 16314 11870
rect 19520 11840 20000 11870
rect 15580 11734 16314 11794
rect 15580 11732 15586 11734
rect 15469 11658 15535 11661
rect 19520 11658 20000 11688
rect 15469 11656 20000 11658
rect 15469 11600 15474 11656
rect 15530 11600 20000 11656
rect 15469 11598 20000 11600
rect 15469 11595 15535 11598
rect 19520 11568 20000 11598
rect 6874 11456 7194 11457
rect 0 11386 480 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 2865 11386 2931 11389
rect 0 11384 2931 11386
rect 0 11328 2870 11384
rect 2926 11328 2931 11384
rect 0 11326 2931 11328
rect 0 11296 480 11326
rect 2865 11323 2931 11326
rect 9857 11250 9923 11253
rect 16389 11250 16455 11253
rect 9857 11248 16455 11250
rect 9857 11192 9862 11248
rect 9918 11192 16394 11248
rect 16450 11192 16455 11248
rect 9857 11190 16455 11192
rect 9857 11187 9923 11190
rect 16389 11187 16455 11190
rect 16849 11250 16915 11253
rect 19520 11250 20000 11280
rect 16849 11248 20000 11250
rect 16849 11192 16854 11248
rect 16910 11192 20000 11248
rect 16849 11190 20000 11192
rect 16849 11187 16915 11190
rect 19520 11160 20000 11190
rect 0 11114 480 11144
rect 3417 11114 3483 11117
rect 0 11112 3483 11114
rect 0 11056 3422 11112
rect 3478 11056 3483 11112
rect 0 11054 3483 11056
rect 0 11024 480 11054
rect 3417 11051 3483 11054
rect 12801 11114 12867 11117
rect 18045 11114 18111 11117
rect 12801 11112 18111 11114
rect 12801 11056 12806 11112
rect 12862 11056 18050 11112
rect 18106 11056 18111 11112
rect 12801 11054 18111 11056
rect 12801 11051 12867 11054
rect 18045 11051 18111 11054
rect 18137 10978 18203 10981
rect 19520 10978 20000 11008
rect 18137 10976 20000 10978
rect 18137 10920 18142 10976
rect 18198 10920 20000 10976
rect 18137 10918 20000 10920
rect 18137 10915 18203 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 19520 10888 20000 10918
rect 15770 10847 16090 10848
rect 0 10706 480 10736
rect 4061 10706 4127 10709
rect 0 10704 4127 10706
rect 0 10648 4066 10704
rect 4122 10648 4127 10704
rect 0 10646 4127 10648
rect 0 10616 480 10646
rect 4061 10643 4127 10646
rect 14641 10706 14707 10709
rect 16849 10706 16915 10709
rect 14641 10704 16915 10706
rect 14641 10648 14646 10704
rect 14702 10648 16854 10704
rect 16910 10648 16915 10704
rect 14641 10646 16915 10648
rect 14641 10643 14707 10646
rect 16849 10643 16915 10646
rect 7833 10570 7899 10573
rect 12433 10570 12499 10573
rect 15377 10570 15443 10573
rect 7833 10568 15443 10570
rect 7833 10512 7838 10568
rect 7894 10512 12438 10568
rect 12494 10512 15382 10568
rect 15438 10512 15443 10568
rect 7833 10510 15443 10512
rect 7833 10507 7899 10510
rect 12433 10507 12499 10510
rect 15377 10507 15443 10510
rect 16665 10570 16731 10573
rect 19520 10570 20000 10600
rect 16665 10568 20000 10570
rect 16665 10512 16670 10568
rect 16726 10512 20000 10568
rect 16665 10510 20000 10512
rect 16665 10507 16731 10510
rect 19520 10480 20000 10510
rect 0 10434 480 10464
rect 4337 10434 4403 10437
rect 0 10432 4403 10434
rect 0 10376 4342 10432
rect 4398 10376 4403 10432
rect 0 10374 4403 10376
rect 0 10344 480 10374
rect 4337 10371 4403 10374
rect 14825 10434 14891 10437
rect 14825 10432 18338 10434
rect 14825 10376 14830 10432
rect 14886 10376 18338 10432
rect 14825 10374 18338 10376
rect 14825 10371 14891 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 10303 13125 10304
rect 2681 10298 2747 10301
rect 4981 10298 5047 10301
rect 2681 10296 5047 10298
rect 2681 10240 2686 10296
rect 2742 10240 4986 10296
rect 5042 10240 5047 10296
rect 2681 10238 5047 10240
rect 2681 10235 2747 10238
rect 4981 10235 5047 10238
rect 14825 10298 14891 10301
rect 18137 10298 18203 10301
rect 14825 10296 18203 10298
rect 14825 10240 14830 10296
rect 14886 10240 18142 10296
rect 18198 10240 18203 10296
rect 14825 10238 18203 10240
rect 14825 10235 14891 10238
rect 18137 10235 18203 10238
rect 18278 10298 18338 10374
rect 19520 10298 20000 10328
rect 18278 10238 20000 10298
rect 7097 10162 7163 10165
rect 9765 10162 9831 10165
rect 7097 10160 9831 10162
rect 7097 10104 7102 10160
rect 7158 10104 9770 10160
rect 9826 10104 9831 10160
rect 7097 10102 9831 10104
rect 7097 10099 7163 10102
rect 9765 10099 9831 10102
rect 13261 10162 13327 10165
rect 16297 10162 16363 10165
rect 13261 10160 16363 10162
rect 13261 10104 13266 10160
rect 13322 10104 16302 10160
rect 16358 10104 16363 10160
rect 13261 10102 16363 10104
rect 13261 10099 13327 10102
rect 16297 10099 16363 10102
rect 17861 10162 17927 10165
rect 18278 10162 18338 10238
rect 19520 10208 20000 10238
rect 17861 10160 18338 10162
rect 17861 10104 17866 10160
rect 17922 10104 18338 10160
rect 17861 10102 18338 10104
rect 17861 10099 17927 10102
rect 0 10026 480 10056
rect 6269 10026 6335 10029
rect 16205 10026 16271 10029
rect 0 9966 6194 10026
rect 0 9936 480 9966
rect 6134 9890 6194 9966
rect 6269 10024 16271 10026
rect 6269 9968 6274 10024
rect 6330 9968 16210 10024
rect 16266 9968 16271 10024
rect 6269 9966 16271 9968
rect 6269 9963 6335 9966
rect 13310 9893 13370 9966
rect 16205 9963 16271 9966
rect 18045 10026 18111 10029
rect 19520 10026 20000 10056
rect 18045 10024 20000 10026
rect 18045 9968 18050 10024
rect 18106 9968 20000 10024
rect 18045 9966 20000 9968
rect 18045 9963 18111 9966
rect 19520 9936 20000 9966
rect 6821 9890 6887 9893
rect 8385 9890 8451 9893
rect 6134 9888 8451 9890
rect 6134 9832 6826 9888
rect 6882 9832 8390 9888
rect 8446 9832 8451 9888
rect 6134 9830 8451 9832
rect 13310 9888 13419 9893
rect 13310 9832 13358 9888
rect 13414 9832 13419 9888
rect 13310 9830 13419 9832
rect 6821 9827 6887 9830
rect 8385 9827 8451 9830
rect 13353 9827 13419 9830
rect 3909 9824 4229 9825
rect 0 9754 480 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 4337 9754 4403 9757
rect 7189 9754 7255 9757
rect 7598 9754 7604 9756
rect 0 9694 3848 9754
rect 0 9664 480 9694
rect 3788 9618 3848 9694
rect 4337 9752 7604 9754
rect 4337 9696 4342 9752
rect 4398 9696 7194 9752
rect 7250 9696 7604 9752
rect 4337 9694 7604 9696
rect 4337 9691 4403 9694
rect 7189 9691 7255 9694
rect 7598 9692 7604 9694
rect 7668 9692 7674 9756
rect 12525 9754 12591 9757
rect 13537 9754 13603 9757
rect 12525 9752 13603 9754
rect 12525 9696 12530 9752
rect 12586 9696 13542 9752
rect 13598 9696 13603 9752
rect 12525 9694 13603 9696
rect 12525 9691 12591 9694
rect 13537 9691 13603 9694
rect 3969 9618 4035 9621
rect 10501 9618 10567 9621
rect 3788 9616 10567 9618
rect 3788 9560 3974 9616
rect 4030 9560 10506 9616
rect 10562 9560 10567 9616
rect 3788 9558 10567 9560
rect 3969 9555 4035 9558
rect 10501 9555 10567 9558
rect 18965 9618 19031 9621
rect 19520 9618 20000 9648
rect 18965 9616 20000 9618
rect 18965 9560 18970 9616
rect 19026 9560 20000 9616
rect 18965 9558 20000 9560
rect 18965 9555 19031 9558
rect 19520 9528 20000 9558
rect 2773 9482 2839 9485
rect 2998 9482 3004 9484
rect 2773 9480 3004 9482
rect 2773 9424 2778 9480
rect 2834 9424 3004 9480
rect 2773 9422 3004 9424
rect 2773 9419 2839 9422
rect 2998 9420 3004 9422
rect 3068 9482 3074 9484
rect 4337 9482 4403 9485
rect 14089 9482 14155 9485
rect 15142 9482 15148 9484
rect 3068 9480 15148 9482
rect 3068 9424 4342 9480
rect 4398 9424 14094 9480
rect 14150 9424 15148 9480
rect 3068 9422 15148 9424
rect 3068 9420 3074 9422
rect 4337 9419 4403 9422
rect 14089 9419 14155 9422
rect 15142 9420 15148 9422
rect 15212 9420 15218 9484
rect 0 9346 480 9376
rect 3693 9346 3759 9349
rect 0 9344 3759 9346
rect 0 9288 3698 9344
rect 3754 9288 3759 9344
rect 0 9286 3759 9288
rect 0 9256 480 9286
rect 3693 9283 3759 9286
rect 4153 9346 4219 9349
rect 6361 9346 6427 9349
rect 4153 9344 6427 9346
rect 4153 9288 4158 9344
rect 4214 9288 6366 9344
rect 6422 9288 6427 9344
rect 4153 9286 6427 9288
rect 4153 9283 4219 9286
rect 6361 9283 6427 9286
rect 9029 9346 9095 9349
rect 11605 9346 11671 9349
rect 9029 9344 11671 9346
rect 9029 9288 9034 9344
rect 9090 9288 11610 9344
rect 11666 9288 11671 9344
rect 9029 9286 11671 9288
rect 9029 9283 9095 9286
rect 11605 9283 11671 9286
rect 18229 9346 18295 9349
rect 19520 9346 20000 9376
rect 18229 9344 20000 9346
rect 18229 9288 18234 9344
rect 18290 9288 20000 9344
rect 18229 9286 20000 9288
rect 18229 9283 18295 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 19520 9256 20000 9286
rect 12805 9215 13125 9216
rect 7373 9212 7439 9213
rect 7373 9210 7420 9212
rect 7328 9208 7420 9210
rect 7328 9152 7378 9208
rect 7328 9150 7420 9152
rect 7373 9148 7420 9150
rect 7484 9148 7490 9212
rect 10409 9210 10475 9213
rect 11329 9210 11395 9213
rect 10409 9208 11395 9210
rect 10409 9152 10414 9208
rect 10470 9152 11334 9208
rect 11390 9152 11395 9208
rect 10409 9150 11395 9152
rect 7373 9147 7439 9148
rect 10409 9147 10475 9150
rect 11329 9147 11395 9150
rect 14365 9210 14431 9213
rect 15469 9210 15535 9213
rect 14365 9208 15535 9210
rect 14365 9152 14370 9208
rect 14426 9152 15474 9208
rect 15530 9152 15535 9208
rect 14365 9150 15535 9152
rect 14365 9147 14431 9150
rect 15469 9147 15535 9150
rect 0 9074 480 9104
rect 8702 9074 8708 9076
rect 0 9014 8708 9074
rect 0 8984 480 9014
rect 8702 9012 8708 9014
rect 8772 9074 8778 9076
rect 9397 9074 9463 9077
rect 8772 9072 9463 9074
rect 8772 9016 9402 9072
rect 9458 9016 9463 9072
rect 8772 9014 9463 9016
rect 8772 9012 8778 9014
rect 9397 9011 9463 9014
rect 8937 8938 9003 8941
rect 13537 8938 13603 8941
rect 8937 8936 13603 8938
rect 8937 8880 8942 8936
rect 8998 8880 13542 8936
rect 13598 8880 13603 8936
rect 8937 8878 13603 8880
rect 8937 8875 9003 8878
rect 13537 8875 13603 8878
rect 13813 8938 13879 8941
rect 16389 8938 16455 8941
rect 13813 8936 16455 8938
rect 13813 8880 13818 8936
rect 13874 8880 16394 8936
rect 16450 8880 16455 8936
rect 13813 8878 16455 8880
rect 13813 8875 13879 8878
rect 16389 8875 16455 8878
rect 18321 8938 18387 8941
rect 19520 8938 20000 8968
rect 18321 8936 20000 8938
rect 18321 8880 18326 8936
rect 18382 8880 20000 8936
rect 18321 8878 20000 8880
rect 18321 8875 18387 8878
rect 19520 8848 20000 8878
rect 6637 8802 6703 8805
rect 9121 8802 9187 8805
rect 6637 8800 9187 8802
rect 6637 8744 6642 8800
rect 6698 8744 9126 8800
rect 9182 8744 9187 8800
rect 6637 8742 9187 8744
rect 6637 8739 6703 8742
rect 9121 8739 9187 8742
rect 3909 8736 4229 8737
rect 0 8666 480 8696
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 1209 8666 1275 8669
rect 0 8664 1275 8666
rect 0 8608 1214 8664
rect 1270 8608 1275 8664
rect 0 8606 1275 8608
rect 0 8576 480 8606
rect 1209 8603 1275 8606
rect 16481 8666 16547 8669
rect 19520 8666 20000 8696
rect 16481 8664 20000 8666
rect 16481 8608 16486 8664
rect 16542 8608 20000 8664
rect 16481 8606 20000 8608
rect 16481 8603 16547 8606
rect 19520 8576 20000 8606
rect 4705 8530 4771 8533
rect 7925 8530 7991 8533
rect 4705 8528 7991 8530
rect 4705 8472 4710 8528
rect 4766 8472 7930 8528
rect 7986 8472 7991 8528
rect 4705 8470 7991 8472
rect 4705 8467 4771 8470
rect 7925 8467 7991 8470
rect 0 8394 480 8424
rect 1669 8394 1735 8397
rect 2773 8394 2839 8397
rect 0 8392 2839 8394
rect 0 8336 1674 8392
rect 1730 8336 2778 8392
rect 2834 8336 2839 8392
rect 0 8334 2839 8336
rect 0 8304 480 8334
rect 1669 8331 1735 8334
rect 2773 8331 2839 8334
rect 3550 8332 3556 8396
rect 3620 8394 3626 8396
rect 4061 8394 4127 8397
rect 12341 8394 12407 8397
rect 3620 8392 12407 8394
rect 3620 8336 4066 8392
rect 4122 8336 12346 8392
rect 12402 8336 12407 8392
rect 3620 8334 12407 8336
rect 3620 8332 3626 8334
rect 4061 8331 4127 8334
rect 12341 8331 12407 8334
rect 15377 8394 15443 8397
rect 15510 8394 15516 8396
rect 15377 8392 15516 8394
rect 15377 8336 15382 8392
rect 15438 8336 15516 8392
rect 15377 8334 15516 8336
rect 15377 8331 15443 8334
rect 15510 8332 15516 8334
rect 15580 8332 15586 8396
rect 18413 8394 18479 8397
rect 19520 8394 20000 8424
rect 18413 8392 20000 8394
rect 18413 8336 18418 8392
rect 18474 8336 20000 8392
rect 18413 8334 20000 8336
rect 18413 8331 18479 8334
rect 19520 8304 20000 8334
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 2129 8122 2195 8125
rect 6637 8122 6703 8125
rect 18045 8122 18111 8125
rect 2129 8120 6703 8122
rect 2129 8064 2134 8120
rect 2190 8064 6642 8120
rect 6698 8064 6703 8120
rect 2129 8062 6703 8064
rect 2129 8059 2195 8062
rect 6637 8059 6703 8062
rect 13264 8120 18111 8122
rect 13264 8064 18050 8120
rect 18106 8064 18111 8120
rect 13264 8062 18111 8064
rect 0 7986 480 8016
rect 5993 7986 6059 7989
rect 0 7984 6059 7986
rect 0 7928 5998 7984
rect 6054 7928 6059 7984
rect 0 7926 6059 7928
rect 0 7896 480 7926
rect 5993 7923 6059 7926
rect 7925 7986 7991 7989
rect 12709 7986 12775 7989
rect 7925 7984 12775 7986
rect 7925 7928 7930 7984
rect 7986 7928 12714 7984
rect 12770 7928 12775 7984
rect 7925 7926 12775 7928
rect 7925 7923 7991 7926
rect 12709 7923 12775 7926
rect 2681 7850 2747 7853
rect 8937 7850 9003 7853
rect 2681 7848 9003 7850
rect 2681 7792 2686 7848
rect 2742 7792 8942 7848
rect 8998 7792 9003 7848
rect 2681 7790 9003 7792
rect 2681 7787 2747 7790
rect 8937 7787 9003 7790
rect 11053 7850 11119 7853
rect 13264 7850 13324 8062
rect 18045 8059 18111 8062
rect 15285 7986 15351 7989
rect 19520 7986 20000 8016
rect 15285 7984 20000 7986
rect 15285 7928 15290 7984
rect 15346 7928 20000 7984
rect 15285 7926 20000 7928
rect 15285 7923 15351 7926
rect 19520 7896 20000 7926
rect 11053 7848 13324 7850
rect 11053 7792 11058 7848
rect 11114 7792 13324 7848
rect 11053 7790 13324 7792
rect 15009 7850 15075 7853
rect 15009 7848 16314 7850
rect 15009 7792 15014 7848
rect 15070 7792 16314 7848
rect 15009 7790 16314 7792
rect 11053 7787 11119 7790
rect 15009 7787 15075 7790
rect 0 7714 480 7744
rect 2129 7714 2195 7717
rect 0 7712 2195 7714
rect 0 7656 2134 7712
rect 2190 7656 2195 7712
rect 0 7654 2195 7656
rect 0 7624 480 7654
rect 2129 7651 2195 7654
rect 10961 7714 11027 7717
rect 12433 7714 12499 7717
rect 10961 7712 12499 7714
rect 10961 7656 10966 7712
rect 11022 7656 12438 7712
rect 12494 7656 12499 7712
rect 10961 7654 12499 7656
rect 16254 7714 16314 7790
rect 19520 7714 20000 7744
rect 16254 7654 20000 7714
rect 10961 7651 11027 7654
rect 12433 7651 12499 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 19520 7624 20000 7654
rect 15770 7583 16090 7584
rect 5073 7578 5139 7581
rect 7649 7578 7715 7581
rect 5073 7576 7715 7578
rect 5073 7520 5078 7576
rect 5134 7520 7654 7576
rect 7710 7520 7715 7576
rect 5073 7518 7715 7520
rect 5073 7515 5139 7518
rect 7649 7515 7715 7518
rect 4889 7442 4955 7445
rect 7189 7442 7255 7445
rect 8569 7442 8635 7445
rect 2592 7440 8635 7442
rect 2592 7384 4894 7440
rect 4950 7384 7194 7440
rect 7250 7384 8574 7440
rect 8630 7384 8635 7440
rect 2592 7382 8635 7384
rect 0 7306 480 7336
rect 2592 7309 2652 7382
rect 4889 7379 4955 7382
rect 7189 7379 7255 7382
rect 8569 7379 8635 7382
rect 12065 7442 12131 7445
rect 16849 7442 16915 7445
rect 12065 7440 16915 7442
rect 12065 7384 12070 7440
rect 12126 7384 16854 7440
rect 16910 7384 16915 7440
rect 12065 7382 16915 7384
rect 12065 7379 12131 7382
rect 16849 7379 16915 7382
rect 2589 7306 2655 7309
rect 0 7304 2655 7306
rect 0 7248 2594 7304
rect 2650 7248 2655 7304
rect 0 7246 2655 7248
rect 0 7216 480 7246
rect 2589 7243 2655 7246
rect 3325 7306 3391 7309
rect 8661 7306 8727 7309
rect 3325 7304 8727 7306
rect 3325 7248 3330 7304
rect 3386 7248 8666 7304
rect 8722 7248 8727 7304
rect 3325 7246 8727 7248
rect 3325 7243 3391 7246
rect 8661 7243 8727 7246
rect 12525 7306 12591 7309
rect 15101 7306 15167 7309
rect 19520 7306 20000 7336
rect 12525 7304 14842 7306
rect 12525 7248 12530 7304
rect 12586 7248 14842 7304
rect 12525 7246 14842 7248
rect 12525 7243 12591 7246
rect 14782 7170 14842 7246
rect 15101 7304 20000 7306
rect 15101 7248 15106 7304
rect 15162 7248 20000 7304
rect 15101 7246 20000 7248
rect 15101 7243 15167 7246
rect 19520 7216 20000 7246
rect 15561 7170 15627 7173
rect 14782 7168 15627 7170
rect 14782 7112 15566 7168
rect 15622 7112 15627 7168
rect 14782 7110 15627 7112
rect 15561 7107 15627 7110
rect 6874 7104 7194 7105
rect 0 7034 480 7064
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 2037 7034 2103 7037
rect 6085 7034 6151 7037
rect 0 7032 6151 7034
rect 0 6976 2042 7032
rect 2098 6976 6090 7032
rect 6146 6976 6151 7032
rect 0 6974 6151 6976
rect 0 6944 480 6974
rect 2037 6971 2103 6974
rect 6085 6971 6151 6974
rect 16297 7034 16363 7037
rect 19520 7034 20000 7064
rect 16297 7032 20000 7034
rect 16297 6976 16302 7032
rect 16358 6976 20000 7032
rect 16297 6974 20000 6976
rect 16297 6971 16363 6974
rect 19520 6944 20000 6974
rect 6177 6898 6243 6901
rect 8937 6898 9003 6901
rect 6177 6896 9003 6898
rect 6177 6840 6182 6896
rect 6238 6840 8942 6896
rect 8998 6840 9003 6896
rect 6177 6838 9003 6840
rect 6177 6835 6243 6838
rect 8937 6835 9003 6838
rect 9857 6898 9923 6901
rect 12893 6898 12959 6901
rect 9857 6896 12959 6898
rect 9857 6840 9862 6896
rect 9918 6840 12898 6896
rect 12954 6840 12959 6896
rect 9857 6838 12959 6840
rect 9857 6835 9923 6838
rect 12893 6835 12959 6838
rect 13169 6898 13235 6901
rect 16573 6898 16639 6901
rect 13169 6896 16639 6898
rect 13169 6840 13174 6896
rect 13230 6840 16578 6896
rect 16634 6840 16639 6896
rect 13169 6838 16639 6840
rect 13169 6835 13235 6838
rect 16573 6835 16639 6838
rect 9673 6762 9739 6765
rect 14273 6762 14339 6765
rect 9673 6760 14339 6762
rect 9673 6704 9678 6760
rect 9734 6704 14278 6760
rect 14334 6704 14339 6760
rect 9673 6702 14339 6704
rect 9673 6699 9739 6702
rect 14273 6699 14339 6702
rect 15193 6762 15259 6765
rect 19520 6762 20000 6792
rect 15193 6760 20000 6762
rect 15193 6704 15198 6760
rect 15254 6704 20000 6760
rect 15193 6702 20000 6704
rect 15193 6699 15259 6702
rect 19520 6672 20000 6702
rect 0 6626 480 6656
rect 2957 6626 3023 6629
rect 0 6624 3023 6626
rect 0 6568 2962 6624
rect 3018 6568 3023 6624
rect 0 6566 3023 6568
rect 0 6536 480 6566
rect 2957 6563 3023 6566
rect 4521 6626 4587 6629
rect 9305 6626 9371 6629
rect 4521 6624 9371 6626
rect 4521 6568 4526 6624
rect 4582 6568 9310 6624
rect 9366 6568 9371 6624
rect 4521 6566 9371 6568
rect 4521 6563 4587 6566
rect 9305 6563 9371 6566
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 5809 6490 5875 6493
rect 7465 6490 7531 6493
rect 5809 6488 7531 6490
rect 5809 6432 5814 6488
rect 5870 6432 7470 6488
rect 7526 6432 7531 6488
rect 5809 6430 7531 6432
rect 5809 6427 5875 6430
rect 7465 6427 7531 6430
rect 0 6354 480 6384
rect 3785 6354 3851 6357
rect 0 6352 3851 6354
rect 0 6296 3790 6352
rect 3846 6296 3851 6352
rect 0 6294 3851 6296
rect 0 6264 480 6294
rect 3785 6291 3851 6294
rect 4705 6354 4771 6357
rect 15377 6354 15443 6357
rect 4705 6352 15443 6354
rect 4705 6296 4710 6352
rect 4766 6296 15382 6352
rect 15438 6296 15443 6352
rect 4705 6294 15443 6296
rect 4705 6291 4771 6294
rect 15377 6291 15443 6294
rect 16481 6354 16547 6357
rect 19520 6354 20000 6384
rect 16481 6352 20000 6354
rect 16481 6296 16486 6352
rect 16542 6296 20000 6352
rect 16481 6294 20000 6296
rect 16481 6291 16547 6294
rect 19520 6264 20000 6294
rect 5441 6218 5507 6221
rect 8385 6218 8451 6221
rect 5441 6216 8451 6218
rect 5441 6160 5446 6216
rect 5502 6160 8390 6216
rect 8446 6160 8451 6216
rect 5441 6158 8451 6160
rect 5441 6155 5507 6158
rect 8385 6155 8451 6158
rect 8569 6218 8635 6221
rect 13261 6218 13327 6221
rect 13537 6218 13603 6221
rect 8569 6216 13603 6218
rect 8569 6160 8574 6216
rect 8630 6160 13266 6216
rect 13322 6160 13542 6216
rect 13598 6160 13603 6216
rect 8569 6158 13603 6160
rect 8569 6155 8635 6158
rect 13261 6155 13327 6158
rect 13537 6155 13603 6158
rect 2313 6082 2379 6085
rect 17861 6082 17927 6085
rect 19520 6082 20000 6112
rect 2313 6080 6746 6082
rect 2313 6024 2318 6080
rect 2374 6024 6746 6080
rect 2313 6022 6746 6024
rect 2313 6019 2379 6022
rect 0 5946 480 5976
rect 3233 5946 3299 5949
rect 0 5944 3299 5946
rect 0 5888 3238 5944
rect 3294 5888 3299 5944
rect 0 5886 3299 5888
rect 0 5856 480 5886
rect 3233 5883 3299 5886
rect 2773 5810 2839 5813
rect 6686 5810 6746 6022
rect 17861 6080 20000 6082
rect 17861 6024 17866 6080
rect 17922 6024 20000 6080
rect 17861 6022 20000 6024
rect 17861 6019 17927 6022
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19520 5992 20000 6022
rect 12805 5951 13125 5952
rect 8753 5948 8819 5949
rect 8702 5884 8708 5948
rect 8772 5946 8819 5948
rect 11421 5946 11487 5949
rect 8772 5944 8864 5946
rect 8814 5888 8864 5944
rect 8772 5886 8864 5888
rect 11421 5944 12680 5946
rect 11421 5888 11426 5944
rect 11482 5888 12680 5944
rect 11421 5886 12680 5888
rect 8772 5884 8819 5886
rect 8753 5883 8819 5884
rect 11421 5883 11487 5886
rect 8753 5810 8819 5813
rect 2773 5808 4170 5810
rect 2773 5752 2778 5808
rect 2834 5752 4170 5808
rect 2773 5750 4170 5752
rect 6686 5808 8819 5810
rect 6686 5752 8758 5808
rect 8814 5752 8819 5808
rect 6686 5750 8819 5752
rect 12620 5810 12680 5886
rect 17309 5810 17375 5813
rect 12620 5808 17375 5810
rect 12620 5752 17314 5808
rect 17370 5752 17375 5808
rect 12620 5750 17375 5752
rect 2773 5747 2839 5750
rect 0 5674 480 5704
rect 3969 5674 4035 5677
rect 0 5672 4035 5674
rect 0 5616 3974 5672
rect 4030 5616 4035 5672
rect 0 5614 4035 5616
rect 4110 5674 4170 5750
rect 8753 5747 8819 5750
rect 17309 5747 17375 5750
rect 17953 5674 18019 5677
rect 4110 5672 18019 5674
rect 4110 5616 17958 5672
rect 18014 5616 18019 5672
rect 4110 5614 18019 5616
rect 0 5584 480 5614
rect 3969 5611 4035 5614
rect 17953 5611 18019 5614
rect 18413 5674 18479 5677
rect 19520 5674 20000 5704
rect 18413 5672 20000 5674
rect 18413 5616 18418 5672
rect 18474 5616 20000 5672
rect 18413 5614 20000 5616
rect 18413 5611 18479 5614
rect 19520 5584 20000 5614
rect 4429 5538 4495 5541
rect 8569 5538 8635 5541
rect 4429 5536 8635 5538
rect 4429 5480 4434 5536
rect 4490 5480 8574 5536
rect 8630 5480 8635 5536
rect 4429 5478 8635 5480
rect 4429 5475 4495 5478
rect 8569 5475 8635 5478
rect 10501 5538 10567 5541
rect 14273 5538 14339 5541
rect 10501 5536 14339 5538
rect 10501 5480 10506 5536
rect 10562 5480 14278 5536
rect 14334 5480 14339 5536
rect 10501 5478 14339 5480
rect 10501 5475 10567 5478
rect 14273 5475 14339 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 4613 5402 4679 5405
rect 6637 5402 6703 5405
rect 4613 5400 6703 5402
rect 4613 5344 4618 5400
rect 4674 5344 6642 5400
rect 6698 5344 6703 5400
rect 4613 5342 6703 5344
rect 4613 5339 4679 5342
rect 6637 5339 6703 5342
rect 7414 5340 7420 5404
rect 7484 5402 7490 5404
rect 8569 5402 8635 5405
rect 7484 5400 8635 5402
rect 7484 5344 8574 5400
rect 8630 5344 8635 5400
rect 7484 5342 8635 5344
rect 7484 5340 7490 5342
rect 8569 5339 8635 5342
rect 11605 5402 11671 5405
rect 13905 5402 13971 5405
rect 11605 5400 13971 5402
rect 11605 5344 11610 5400
rect 11666 5344 13910 5400
rect 13966 5344 13971 5400
rect 11605 5342 13971 5344
rect 11605 5339 11671 5342
rect 13905 5339 13971 5342
rect 17769 5402 17835 5405
rect 19520 5402 20000 5432
rect 17769 5400 20000 5402
rect 17769 5344 17774 5400
rect 17830 5344 20000 5400
rect 17769 5342 20000 5344
rect 17769 5339 17835 5342
rect 19520 5312 20000 5342
rect 0 5266 480 5296
rect 5901 5266 5967 5269
rect 0 5264 5967 5266
rect 0 5208 5906 5264
rect 5962 5208 5967 5264
rect 0 5206 5967 5208
rect 0 5176 480 5206
rect 5901 5203 5967 5206
rect 6085 5266 6151 5269
rect 8385 5266 8451 5269
rect 6085 5264 8451 5266
rect 6085 5208 6090 5264
rect 6146 5208 8390 5264
rect 8446 5208 8451 5264
rect 6085 5206 8451 5208
rect 6085 5203 6151 5206
rect 8385 5203 8451 5206
rect 9397 5266 9463 5269
rect 14549 5266 14615 5269
rect 9397 5264 14615 5266
rect 9397 5208 9402 5264
rect 9458 5208 14554 5264
rect 14610 5208 14615 5264
rect 9397 5206 14615 5208
rect 9397 5203 9463 5206
rect 14549 5203 14615 5206
rect 3877 5130 3943 5133
rect 4889 5130 4955 5133
rect 8845 5130 8911 5133
rect 3877 5128 8911 5130
rect 3877 5072 3882 5128
rect 3938 5072 4894 5128
rect 4950 5072 8850 5128
rect 8906 5072 8911 5128
rect 3877 5070 8911 5072
rect 3877 5067 3943 5070
rect 4889 5067 4955 5070
rect 8845 5067 8911 5070
rect 10685 5130 10751 5133
rect 15837 5130 15903 5133
rect 10685 5128 15903 5130
rect 10685 5072 10690 5128
rect 10746 5072 15842 5128
rect 15898 5072 15903 5128
rect 10685 5070 15903 5072
rect 10685 5067 10751 5070
rect 15837 5067 15903 5070
rect 17861 5130 17927 5133
rect 19520 5130 20000 5160
rect 17861 5128 20000 5130
rect 17861 5072 17866 5128
rect 17922 5072 20000 5128
rect 17861 5070 20000 5072
rect 17861 5067 17927 5070
rect 19520 5040 20000 5070
rect 0 4994 480 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 0 4904 480 4934
rect 4061 4931 4127 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 5349 4858 5415 4861
rect 8201 4858 8267 4861
rect 5349 4856 5458 4858
rect 5349 4800 5354 4856
rect 5410 4800 5458 4856
rect 5349 4795 5458 4800
rect 8201 4856 12680 4858
rect 8201 4800 8206 4856
rect 8262 4800 12680 4856
rect 8201 4798 12680 4800
rect 8201 4795 8267 4798
rect 5398 4722 5458 4795
rect 7189 4722 7255 4725
rect 5398 4720 7255 4722
rect 5398 4664 7194 4720
rect 7250 4664 7255 4720
rect 5398 4662 7255 4664
rect 12620 4722 12680 4798
rect 13721 4722 13787 4725
rect 12620 4720 13787 4722
rect 12620 4664 13726 4720
rect 13782 4664 13787 4720
rect 12620 4662 13787 4664
rect 7189 4659 7255 4662
rect 13721 4659 13787 4662
rect 16849 4722 16915 4725
rect 19520 4722 20000 4752
rect 16849 4720 20000 4722
rect 16849 4664 16854 4720
rect 16910 4664 20000 4720
rect 16849 4662 20000 4664
rect 16849 4659 16915 4662
rect 19520 4632 20000 4662
rect 0 4586 480 4616
rect 3877 4586 3943 4589
rect 0 4584 3943 4586
rect 0 4528 3882 4584
rect 3938 4528 3943 4584
rect 0 4526 3943 4528
rect 0 4496 480 4526
rect 3877 4523 3943 4526
rect 4889 4586 4955 4589
rect 9029 4586 9095 4589
rect 9213 4586 9279 4589
rect 4889 4584 9279 4586
rect 4889 4528 4894 4584
rect 4950 4528 9034 4584
rect 9090 4528 9218 4584
rect 9274 4528 9279 4584
rect 4889 4526 9279 4528
rect 4889 4523 4955 4526
rect 9029 4523 9095 4526
rect 9213 4523 9279 4526
rect 10685 4450 10751 4453
rect 15561 4450 15627 4453
rect 10685 4448 15627 4450
rect 10685 4392 10690 4448
rect 10746 4392 15566 4448
rect 15622 4392 15627 4448
rect 10685 4390 15627 4392
rect 10685 4387 10751 4390
rect 15561 4387 15627 4390
rect 18229 4450 18295 4453
rect 19520 4450 20000 4480
rect 18229 4448 20000 4450
rect 18229 4392 18234 4448
rect 18290 4392 20000 4448
rect 18229 4390 20000 4392
rect 18229 4387 18295 4390
rect 3909 4384 4229 4385
rect 0 4314 480 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19520 4360 20000 4390
rect 15770 4319 16090 4320
rect 1301 4314 1367 4317
rect 0 4312 1367 4314
rect 0 4256 1306 4312
rect 1362 4256 1367 4312
rect 0 4254 1367 4256
rect 0 4224 480 4254
rect 1301 4251 1367 4254
rect 5717 4314 5783 4317
rect 8753 4314 8819 4317
rect 5717 4312 8819 4314
rect 5717 4256 5722 4312
rect 5778 4256 8758 4312
rect 8814 4256 8819 4312
rect 5717 4254 8819 4256
rect 5717 4251 5783 4254
rect 8753 4251 8819 4254
rect 12525 4178 12591 4181
rect 15377 4178 15443 4181
rect 12525 4176 15443 4178
rect 12525 4120 12530 4176
rect 12586 4120 15382 4176
rect 15438 4120 15443 4176
rect 12525 4118 15443 4120
rect 12525 4115 12591 4118
rect 15377 4115 15443 4118
rect 3366 3980 3372 4044
rect 3436 4042 3442 4044
rect 16849 4042 16915 4045
rect 3436 4040 16915 4042
rect 3436 3984 16854 4040
rect 16910 3984 16915 4040
rect 3436 3982 16915 3984
rect 3436 3980 3442 3982
rect 16849 3979 16915 3982
rect 17401 4042 17467 4045
rect 19520 4042 20000 4072
rect 17401 4040 20000 4042
rect 17401 3984 17406 4040
rect 17462 3984 20000 4040
rect 17401 3982 20000 3984
rect 17401 3979 17467 3982
rect 19520 3952 20000 3982
rect 0 3906 480 3936
rect 1393 3906 1459 3909
rect 0 3904 1459 3906
rect 0 3848 1398 3904
rect 1454 3848 1459 3904
rect 0 3846 1459 3848
rect 0 3816 480 3846
rect 1393 3843 1459 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 18229 3770 18295 3773
rect 19520 3770 20000 3800
rect 18229 3768 20000 3770
rect 18229 3712 18234 3768
rect 18290 3712 20000 3768
rect 18229 3710 20000 3712
rect 18229 3707 18295 3710
rect 19520 3680 20000 3710
rect 0 3634 480 3664
rect 1577 3634 1643 3637
rect 14917 3634 14983 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 480 3574
rect 1577 3571 1643 3574
rect 1718 3632 14983 3634
rect 1718 3576 14922 3632
rect 14978 3576 14983 3632
rect 1718 3574 14983 3576
rect 1209 3498 1275 3501
rect 1718 3498 1778 3574
rect 14917 3571 14983 3574
rect 1209 3496 1778 3498
rect 1209 3440 1214 3496
rect 1270 3440 1778 3496
rect 1209 3438 1778 3440
rect 10317 3498 10383 3501
rect 11789 3498 11855 3501
rect 10317 3496 11855 3498
rect 10317 3440 10322 3496
rect 10378 3440 11794 3496
rect 11850 3440 11855 3496
rect 10317 3438 11855 3440
rect 1209 3435 1275 3438
rect 10317 3435 10383 3438
rect 11789 3435 11855 3438
rect 17769 3498 17835 3501
rect 19520 3498 20000 3528
rect 17769 3496 20000 3498
rect 17769 3440 17774 3496
rect 17830 3440 20000 3496
rect 17769 3438 20000 3440
rect 17769 3435 17835 3438
rect 19520 3408 20000 3438
rect 3909 3296 4229 3297
rect 0 3226 480 3256
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 2865 3226 2931 3229
rect 0 3224 2931 3226
rect 0 3168 2870 3224
rect 2926 3168 2931 3224
rect 0 3166 2931 3168
rect 0 3136 480 3166
rect 2865 3163 2931 3166
rect 3734 3028 3740 3092
rect 3804 3090 3810 3092
rect 16297 3090 16363 3093
rect 19520 3090 20000 3120
rect 3804 3088 20000 3090
rect 3804 3032 16302 3088
rect 16358 3032 20000 3088
rect 3804 3030 20000 3032
rect 3804 3028 3810 3030
rect 16297 3027 16363 3030
rect 19520 3000 20000 3030
rect 0 2954 480 2984
rect 4061 2954 4127 2957
rect 0 2952 4127 2954
rect 0 2896 4066 2952
rect 4122 2896 4127 2952
rect 0 2894 4127 2896
rect 0 2864 480 2894
rect 4061 2891 4127 2894
rect 5257 2954 5323 2957
rect 9581 2954 9647 2957
rect 5257 2952 9647 2954
rect 5257 2896 5262 2952
rect 5318 2896 9586 2952
rect 9642 2896 9647 2952
rect 5257 2894 9647 2896
rect 5257 2891 5323 2894
rect 9581 2891 9647 2894
rect 11145 2954 11211 2957
rect 16246 2954 16252 2956
rect 11145 2952 16252 2954
rect 11145 2896 11150 2952
rect 11206 2896 16252 2952
rect 11145 2894 16252 2896
rect 11145 2891 11211 2894
rect 16246 2892 16252 2894
rect 16316 2892 16322 2956
rect 16849 2818 16915 2821
rect 19520 2818 20000 2848
rect 16849 2816 20000 2818
rect 16849 2760 16854 2816
rect 16910 2760 20000 2816
rect 16849 2758 20000 2760
rect 16849 2755 16915 2758
rect 6874 2752 7194 2753
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 19520 2728 20000 2758
rect 12805 2687 13125 2688
rect 1393 2682 1459 2685
rect 2998 2682 3004 2684
rect 1393 2680 3004 2682
rect 1393 2624 1398 2680
rect 1454 2624 3004 2680
rect 1393 2622 3004 2624
rect 1393 2619 1459 2622
rect 2998 2620 3004 2622
rect 3068 2620 3074 2684
rect 3325 2682 3391 2685
rect 3550 2682 3556 2684
rect 3325 2680 3556 2682
rect 3325 2624 3330 2680
rect 3386 2624 3556 2680
rect 3325 2622 3556 2624
rect 3325 2619 3391 2622
rect 3550 2620 3556 2622
rect 3620 2620 3626 2684
rect 0 2546 480 2576
rect 3601 2546 3667 2549
rect 0 2544 3667 2546
rect 0 2488 3606 2544
rect 3662 2488 3667 2544
rect 0 2486 3667 2488
rect 0 2456 480 2486
rect 3601 2483 3667 2486
rect 4613 2546 4679 2549
rect 9029 2546 9095 2549
rect 4613 2544 9095 2546
rect 4613 2488 4618 2544
rect 4674 2488 9034 2544
rect 9090 2488 9095 2544
rect 4613 2486 9095 2488
rect 4613 2483 4679 2486
rect 9029 2483 9095 2486
rect 3182 2348 3188 2412
rect 3252 2410 3258 2412
rect 16481 2410 16547 2413
rect 3252 2408 16547 2410
rect 3252 2352 16486 2408
rect 16542 2352 16547 2408
rect 3252 2350 16547 2352
rect 3252 2348 3258 2350
rect 16481 2347 16547 2350
rect 17217 2410 17283 2413
rect 19520 2410 20000 2440
rect 17217 2408 20000 2410
rect 17217 2352 17222 2408
rect 17278 2352 20000 2408
rect 17217 2350 20000 2352
rect 17217 2347 17283 2350
rect 19520 2320 20000 2350
rect 0 2274 480 2304
rect 3693 2274 3759 2277
rect 0 2272 3759 2274
rect 0 2216 3698 2272
rect 3754 2216 3759 2272
rect 0 2214 3759 2216
rect 0 2184 480 2214
rect 3693 2211 3759 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2143 16090 2144
rect 16481 2138 16547 2141
rect 19520 2138 20000 2168
rect 16481 2136 20000 2138
rect 16481 2080 16486 2136
rect 16542 2080 20000 2136
rect 16481 2078 20000 2080
rect 16481 2075 16547 2078
rect 19520 2048 20000 2078
rect 0 1866 480 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 480 1806
rect 3417 1803 3483 1806
rect 16205 1866 16271 1869
rect 19520 1866 20000 1896
rect 16205 1864 20000 1866
rect 16205 1808 16210 1864
rect 16266 1808 20000 1864
rect 16205 1806 20000 1808
rect 16205 1803 16271 1806
rect 19520 1776 20000 1806
rect 0 1594 480 1624
rect 4981 1594 5047 1597
rect 0 1592 5047 1594
rect 0 1536 4986 1592
rect 5042 1536 5047 1592
rect 0 1534 5047 1536
rect 0 1504 480 1534
rect 4981 1531 5047 1534
rect 16757 1458 16823 1461
rect 19520 1458 20000 1488
rect 16757 1456 20000 1458
rect 16757 1400 16762 1456
rect 16818 1400 20000 1456
rect 16757 1398 20000 1400
rect 16757 1395 16823 1398
rect 19520 1368 20000 1398
rect 0 1186 480 1216
rect 4061 1186 4127 1189
rect 0 1184 4127 1186
rect 0 1128 4066 1184
rect 4122 1128 4127 1184
rect 0 1126 4127 1128
rect 0 1096 480 1126
rect 4061 1123 4127 1126
rect 17033 1186 17099 1189
rect 19520 1186 20000 1216
rect 17033 1184 20000 1186
rect 17033 1128 17038 1184
rect 17094 1128 20000 1184
rect 17033 1126 20000 1128
rect 17033 1123 17099 1126
rect 19520 1096 20000 1126
rect 0 914 480 944
rect 3693 914 3759 917
rect 0 912 3759 914
rect 0 856 3698 912
rect 3754 856 3759 912
rect 0 854 3759 856
rect 0 824 480 854
rect 3693 851 3759 854
rect 18045 778 18111 781
rect 19520 778 20000 808
rect 18045 776 20000 778
rect 18045 720 18050 776
rect 18106 720 20000 776
rect 18045 718 20000 720
rect 18045 715 18111 718
rect 19520 688 20000 718
rect 0 506 480 536
rect 3325 506 3391 509
rect 0 504 3391 506
rect 0 448 3330 504
rect 3386 448 3391 504
rect 0 446 3391 448
rect 0 416 480 446
rect 3325 443 3391 446
rect 17769 506 17835 509
rect 19520 506 20000 536
rect 17769 504 20000 506
rect 17769 448 17774 504
rect 17830 448 20000 504
rect 17769 446 20000 448
rect 17769 443 17835 446
rect 19520 416 20000 446
rect 0 234 480 264
rect 3141 234 3207 237
rect 0 232 3207 234
rect 0 176 3146 232
rect 3202 176 3207 232
rect 0 174 3207 176
rect 0 144 480 174
rect 3141 171 3207 174
rect 16481 234 16547 237
rect 19520 234 20000 264
rect 16481 232 20000 234
rect 16481 176 16486 232
rect 16542 176 20000 232
rect 16481 174 20000 176
rect 16481 171 16547 174
rect 19520 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 16252 14452 16316 14516
rect 3372 14376 3436 14380
rect 3372 14320 3386 14376
rect 3386 14320 3436 14376
rect 3372 14316 3436 14320
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 3188 13772 3252 13836
rect 3740 13772 3804 13836
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 15148 13500 15212 13564
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 7604 12064 7668 12068
rect 7604 12008 7654 12064
rect 7654 12008 7668 12064
rect 7604 12004 7668 12008
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 15516 11732 15580 11796
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 7604 9692 7668 9756
rect 3004 9420 3068 9484
rect 15148 9420 15212 9484
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 7420 9208 7484 9212
rect 7420 9152 7434 9208
rect 7434 9152 7484 9208
rect 7420 9148 7484 9152
rect 8708 9012 8772 9076
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 3556 8332 3620 8396
rect 15516 8332 15580 8396
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 8708 5944 8772 5948
rect 8708 5888 8758 5944
rect 8758 5888 8772 5944
rect 8708 5884 8772 5888
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 7420 5340 7484 5404
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 3372 3980 3436 4044
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 3740 3028 3804 3092
rect 16252 2892 16316 2956
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 3004 2620 3068 2684
rect 3556 2620 3620 2684
rect 3188 2348 3252 2412
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3371 14380 3437 14381
rect 3371 14316 3372 14380
rect 3436 14316 3437 14380
rect 3371 14315 3437 14316
rect 3187 13836 3253 13837
rect 3187 13772 3188 13836
rect 3252 13772 3253 13836
rect 3187 13771 3253 13772
rect 3003 9484 3069 9485
rect 3003 9420 3004 9484
rect 3068 9420 3069 9484
rect 3003 9419 3069 9420
rect 3006 2685 3066 9419
rect 3003 2684 3069 2685
rect 3003 2620 3004 2684
rect 3068 2620 3069 2684
rect 3003 2619 3069 2620
rect 3190 2413 3250 13771
rect 3374 4045 3434 14315
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3739 13836 3805 13837
rect 3739 13772 3740 13836
rect 3804 13772 3805 13836
rect 3739 13771 3805 13772
rect 3555 8396 3621 8397
rect 3555 8332 3556 8396
rect 3620 8332 3621 8396
rect 3555 8331 3621 8332
rect 3371 4044 3437 4045
rect 3371 3980 3372 4044
rect 3436 3980 3437 4044
rect 3371 3979 3437 3980
rect 3558 2685 3618 8331
rect 3742 3093 3802 13771
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3739 3092 3805 3093
rect 3739 3028 3740 3092
rect 3804 3028 3805 3092
rect 3739 3027 3805 3028
rect 3555 2684 3621 2685
rect 3555 2620 3556 2684
rect 3620 2620 3621 2684
rect 3555 2619 3621 2620
rect 3187 2412 3253 2413
rect 3187 2348 3188 2412
rect 3252 2348 3253 2412
rect 3187 2347 3253 2348
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 7603 12068 7669 12069
rect 7603 12004 7604 12068
rect 7668 12004 7669 12068
rect 7603 12003 7669 12004
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 7606 9757 7666 12003
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 7603 9756 7669 9757
rect 7603 9692 7604 9756
rect 7668 9692 7669 9756
rect 7603 9691 7669 9692
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 7419 9212 7485 9213
rect 7419 9148 7420 9212
rect 7484 9148 7485 9212
rect 7419 9147 7485 9148
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 7422 5405 7482 9147
rect 8707 9076 8773 9077
rect 8707 9012 8708 9076
rect 8772 9012 8773 9076
rect 8707 9011 8773 9012
rect 8710 5949 8770 9011
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 8707 5948 8773 5949
rect 8707 5884 8708 5948
rect 8772 5884 8773 5948
rect 8707 5883 8773 5884
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 7419 5404 7485 5405
rect 7419 5340 7420 5404
rect 7484 5340 7485 5404
rect 7419 5339 7485 5340
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 15770 14176 16090 14736
rect 16251 14516 16317 14517
rect 16251 14452 16252 14516
rect 16316 14452 16317 14516
rect 16251 14451 16317 14452
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15147 13564 15213 13565
rect 15147 13500 15148 13564
rect 15212 13500 15213 13564
rect 15147 13499 15213 13500
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 15150 9485 15210 13499
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15515 11796 15581 11797
rect 15515 11732 15516 11796
rect 15580 11732 15581 11796
rect 15515 11731 15581 11732
rect 15147 9484 15213 9485
rect 15147 9420 15148 9484
rect 15212 9420 15213 9484
rect 15147 9419 15213 9420
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 15518 8397 15578 11731
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15515 8396 15581 8397
rect 15515 8332 15516 8396
rect 15580 8332 15581 8396
rect 15515 8331 15581 8332
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 2208 16090 3232
rect 16254 2957 16314 14451
rect 16251 2956 16317 2957
rect 16251 2892 16252 2956
rect 16316 2892 16317 2956
rect 16251 2891 16317 2892
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1748 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _44_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1606256979
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1606256979
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2760 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4784 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4324 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 3772 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606256979
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_38
timestamp 1606256979
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_49
timestamp 1606256979
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1606256979
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55
timestamp 1606256979
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5980 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _20_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1606256979
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1606256979
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7176 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1606256979
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1606256979
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7820 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7912 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9660 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606256979
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606256979
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1606256979
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1606256979
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1606256979
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1606256979
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1606256979
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606256979
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13432 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14352 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14168 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_131 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143
timestamp 1606256979
transform 1 0 14260 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1606256979
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1606256979
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1606256979
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1606256979
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15456 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_164
timestamp 1606256979
transform 1 0 16192 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1606256979
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1606256979
transform 1 0 16744 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1606256979
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1606256979
transform 1 0 17480 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_S_FTB01
timestamp 1606256979
transform 1 0 17204 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606256979
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606256979
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1606256979
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1606256979
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4784 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1606256979
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_38
timestamp 1606256979
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5796 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1606256979
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7452 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1606256979
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_78
timestamp 1606256979
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10304 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1606256979
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp 1606256979
transform 1 0 10028 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11960 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1606256979
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1606256979
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1606256979
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1606256979
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_N_FTB01
timestamp 1606256979
transform 1 0 17756 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1606256979
transform 1 0 17020 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1606256979
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_179
timestamp 1606256979
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1606256979
transform 1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2852 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1606256979
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1606256979
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4600 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_35
timestamp 1606256979
transform 1 0 4324 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5612 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1606256979
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1606256979
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_78 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8280 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8832 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10488 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1606256979
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_108
timestamp 1606256979
transform 1 0 11040 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1606256979
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12972 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_126
timestamp 1606256979
transform 1 0 12696 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1606256979
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 16100 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14628 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_156
timestamp 1606256979
transform 1 0 15456 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp 1606256979
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 16652 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 17204 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_167
timestamp 1606256979
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1606256979
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1606256979
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1606256979
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1840 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1606256979
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4140 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_top_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp 1606256979
transform 1 0 3312 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1606256979
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606256979
transform 1 0 6808 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5152 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1606256979
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1606256979
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1606256979
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 9016 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1606256979
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606256979
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_102
timestamp 1606256979
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10764 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1606256979
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1606256979
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1606256979
transform 1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 12788 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1606256979
transform 1 0 13064 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1606256979
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1606256979
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606256979
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_163
timestamp 1606256979
transform 1 0 16100 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_1_S_FTB01
timestamp 1606256979
transform 1 0 17756 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16744 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_169
timestamp 1606256979
transform 1 0 16652 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_179
timestamp 1606256979
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_187
timestamp 1606256979
transform 1 0 18308 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1564 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606256979
transform 1 0 4232 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3220 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1606256979
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp 1606256979
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_37
timestamp 1606256979
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1606256979
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1606256979
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606256979
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9476 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_88
timestamp 1606256979
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1606256979
transform 1 0 10948 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606256979
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_139
timestamp 1606256979
transform 1 0 13892 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14996 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1606256979
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16652 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_167
timestamp 1606256979
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1606256979
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606256979
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1606256979
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2116 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_9
timestamp 1606256979
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_20
timestamp 1606256979
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1606256979
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1606256979
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1606256979
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3220 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 3036 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp 1606256979
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4416 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606256979
transform 1 0 4048 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1606256979
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 5428 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1606256979
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1606256979
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp 1606256979
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 6348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606256979
transform 1 0 8096 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8464 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp 1606256979
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1606256979
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_80
timestamp 1606256979
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606256979
transform 1 0 9844 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10304 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10672 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1606256979
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_98
timestamp 1606256979
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606256979
transform 1 0 11960 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 12420 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 1606256979
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1606256979
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606256979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 13432 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12788 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1606256979
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1606256979
transform 1 0 12696 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_136
timestamp 1606256979
transform 1 0 13616 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1606256979
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1606256979
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16284 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1606256979
transform 1 0 14996 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606256979
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1606256979
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1606256979
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 17940 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1606256979
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_181
timestamp 1606256979
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_187
timestamp 1606256979
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1606256979
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606256979
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2208 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_10
timestamp 1606256979
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4232 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1606256979
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5244 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_43
timestamp 1606256979
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1606256979
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606256979
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7820 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 7452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1606256979
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_72
timestamp 1606256979
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10304 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1606256979
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp 1606256979
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12328 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11316 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1606256979
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1606256979
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_138
timestamp 1606256979
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15640 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17296 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1606256979
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_185
timestamp 1606256979
transform 1 0 18124 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1606256979
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 1656 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2668 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1606256979
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1606256979
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1606256979
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606256979
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1606256979
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_96
timestamp 1606256979
transform 1 0 9936 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606256979
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 13616 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606256979
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15272 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1606256979
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1606256979
transform 1 0 16100 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606256979
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16468 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_176
timestamp 1606256979
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606256979
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1606256979
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1564 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606256979
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_21
timestamp 1606256979
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1606256979
transform 1 0 4416 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_40
timestamp 1606256979
transform 1 0 4784 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5888 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1606256979
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1606256979
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606256979
transform 1 0 7912 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1606256979
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_78
timestamp 1606256979
transform 1 0 8280 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_top_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9844 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 11868 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp 1606256979
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1606256979
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1606256979
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1606256979
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16468 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1606256979
transform 1 0 17480 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_176
timestamp 1606256979
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_187
timestamp 1606256979
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2484 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1606256979
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4140 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 1606256979
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606256979
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_49
timestamp 1606256979
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_55
timestamp 1606256979
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6900 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7912 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 1606256979
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_83
timestamp 1606256979
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10580 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8924 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1606256979
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 12604 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1606256979
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14168 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1606256979
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1606256979
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606256979
transform 1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16284 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1606256979
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_163
timestamp 1606256979
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606256979
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1606256979
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1606256979
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4784 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_25
timestamp 1606256979
transform 1 0 3404 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 1606256979
transform 1 0 4416 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 6808 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1606256979
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1606256979
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606256979
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_74
timestamp 1606256979
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1606256979
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10304 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606256979
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1606256979
transform 1 0 10212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11316 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1606256979
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1606256979
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1606256979
transform 1 0 12788 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1606256979
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15732 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606256979
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1606256979
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1606256979
transform 1 0 17388 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1606256979
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1606256979
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1606256979
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606256979
transform 1 0 1472 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_14
timestamp 1606256979
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1606256979
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2576 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1606256979
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_25
timestamp 1606256979
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1606256979
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_41
timestamp 1606256979
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4140 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606256979
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1606256979
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1606256979
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1606256979
transform 1 0 6440 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 8464 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1606256979
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_83
timestamp 1606256979
transform 1 0 8740 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1606256979
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8832 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_86
timestamp 1606256979
transform 1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11408 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11132 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1606256979
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 14352 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13156 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1606256979
transform 1 0 13984 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1606256979
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_128
timestamp 1606256979
transform 1 0 12880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 16284 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 14904 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_148
timestamp 1606256979
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_166
timestamp 1606256979
transform 1 0 16376 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1606256979
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1606256979
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 17848 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1606256979
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606256979
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1606256979
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_180
timestamp 1606256979
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1606256979
transform 1 0 18216 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1606256979
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2392 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1606256979
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4048 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1606256979
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7544 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1606256979
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_97
timestamp 1606256979
transform 1 0 10028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1606256979
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13708 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_136
timestamp 1606256979
transform 1 0 13616 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14536 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1606256979
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606256979
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1606256979
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1606256979
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606256979
transform 1 0 3036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1606256979
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1606256979
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5060 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1606256979
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606256979
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1606256979
transform 1 0 8464 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_66
timestamp 1606256979
transform 1 0 7176 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1606256979
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1606256979
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12604 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11316 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1606256979
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1606256979
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_124
timestamp 1606256979
transform 1 0 12512 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606256979
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1606256979
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_top_ipin_0.prog_clk
timestamp 1606256979
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1606256979
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1606256979
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16928 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606256979
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1606256979
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1748 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606256979
transform 1 0 3404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4140 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_23
timestamp 1606256979
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1606256979
transform 1 0 3772 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1606256979
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8464 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_71
timestamp 1606256979
transform 1 0 7636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp 1606256979
transform 1 0 8372 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10488 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9476 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1606256979
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_100
timestamp 1606256979
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606256979
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 13892 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12880 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1606256979
transform 1 0 12788 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1606256979
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15548 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1606256979
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1606256979
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16560 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_177
timestamp 1606256979
transform 1 0 17388 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1606256979
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1606256979
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606256979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 1606256979
transform 1 0 4876 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1606256979
transform 1 0 6440 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1606256979
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1606256979
transform 1 0 8188 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10396 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606256979
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1606256979
transform 1 0 9936 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_100
timestamp 1606256979
transform 1 0 10304 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11960 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_110
timestamp 1606256979
transform 1 0 11224 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1606256979
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1606256979
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1606256979
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606256979
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_178
timestamp 1606256979
transform 1 0 17480 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_184
timestamp 1606256979
transform 1 0 18032 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606256979
transform 1 0 1656 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1606256979
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1606256979
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2668 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606256979
transform 1 0 3680 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4232 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1606256979
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_31
timestamp 1606256979
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_21
timestamp 1606256979
transform 1 0 3036 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606256979
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_44
timestamp 1606256979
transform 1 0 5152 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_43
timestamp 1606256979
transform 1 0 5060 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5428 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5428 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1606256979
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1606256979
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1606256979
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1606256979
transform 1 0 8648 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_67
timestamp 1606256979
transform 1 0 7268 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_79
timestamp 1606256979
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9108 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1606256979
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_96
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_102
timestamp 1606256979
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606256979
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1606256979
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10948 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_112
timestamp 1606256979
transform 1 0 11408 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_106
timestamp 1606256979
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_116
timestamp 1606256979
transform 1 0 11776 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_132
timestamp 1606256979
transform 1 0 13248 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_144
timestamp 1606256979
transform 1 0 14352 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 1606256979
transform 1 0 12880 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_140
timestamp 1606256979
transform 1 0 13984 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_156
timestamp 1606256979
transform 1 0 15456 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606256979
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606256979
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_168
timestamp 1606256979
transform 1 0 16560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1606256979
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606256979
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1606256979
transform 1 0 2300 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1606256979
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1606256979
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1606256979
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606256979
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1606256979
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1606256979
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_43
timestamp 1606256979
transform 1 0 5060 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_47
timestamp 1606256979
transform 1 0 5428 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606256979
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_N_FTB01
timestamp 1606256979
transform 1 0 8004 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1606256979
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1606256979
transform 1 0 8556 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1606256979
transform 1 0 9660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_105
timestamp 1606256979
transform 1 0 10764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1606256979
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606256979
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1606256979
transform 1 0 14168 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_135
timestamp 1606256979
transform 1 0 13524 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_141
timestamp 1606256979
transform 1 0 14076 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_148
timestamp 1606256979
transform 1 0 14720 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1606256979
transform 1 0 15824 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606256979
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606256979
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_168
timestamp 1606256979
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1606256979
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606256979
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1606256979
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1606256979
transform 1 0 1748 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 1606256979
transform 1 0 2300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606256979
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_21
timestamp 1606256979
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606256979
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 6256 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1606256979
transform 1 0 5152 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_49
timestamp 1606256979
transform 1 0 5612 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1606256979
transform 1 0 6164 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1606256979
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1606256979
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606256979
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1606256979
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1606256979
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1606256979
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1606256979
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1606256979
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606256979
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1606256979
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1606256979
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1606256979
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_180
timestamp 1606256979
transform 1 0 17664 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606256979
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal3 s 19520 16736 20000 16856 6 REGIN_FEEDTHROUGH
port 0 nsew default input
rlabel metal2 s 18234 16520 18290 17000 6 REGOUT_FEEDTHROUGH
port 1 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 SC_IN_BOT
port 2 nsew default input
rlabel metal2 s 1674 16520 1730 17000 6 SC_IN_TOP
port 3 nsew default input
rlabel metal2 s 17590 0 17646 480 6 SC_OUT_BOT
port 4 nsew default tristate
rlabel metal2 s 4986 16520 5042 17000 6 SC_OUT_TOP
port 5 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal2 s 11242 0 11298 480 6 bottom_grid_pin_10_
port 7 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 bottom_grid_pin_11_
port 8 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 bottom_grid_pin_13_
port 10 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 bottom_grid_pin_14_
port 11 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 bottom_grid_pin_15_
port 12 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 bottom_grid_pin_1_
port 13 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 bottom_grid_pin_2_
port 14 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_3_
port 15 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 bottom_grid_pin_4_
port 16 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 bottom_grid_pin_5_
port 17 nsew default tristate
rlabel metal2 s 7562 0 7618 480 6 bottom_grid_pin_6_
port 18 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 bottom_grid_pin_7_
port 19 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 bottom_grid_pin_8_
port 20 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 bottom_grid_pin_9_
port 21 nsew default tristate
rlabel metal2 s 386 0 442 480 6 ccff_head
port 22 nsew default input
rlabel metal2 s 1214 0 1270 480 6 ccff_tail
port 23 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[0]
port 24 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[10]
port 25 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 26 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[12]
port 27 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[13]
port 28 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[14]
port 29 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[15]
port 30 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[16]
port 31 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[17]
port 32 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[18]
port 33 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[19]
port 34 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[1]
port 35 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[2]
port 36 nsew default input
rlabel metal3 s 0 7896 480 8016 6 chanx_left_in[3]
port 37 nsew default input
rlabel metal3 s 0 8304 480 8424 6 chanx_left_in[4]
port 38 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[5]
port 39 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[6]
port 40 nsew default input
rlabel metal3 s 0 9256 480 9376 6 chanx_left_in[7]
port 41 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[8]
port 42 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[9]
port 43 nsew default input
rlabel metal3 s 0 144 480 264 6 chanx_left_out[0]
port 44 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 chanx_left_out[10]
port 45 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[11]
port 46 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_out[12]
port 47 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chanx_left_out[13]
port 48 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_out[14]
port 49 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 chanx_left_out[15]
port 50 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[16]
port 51 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 chanx_left_out[17]
port 52 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[18]
port 53 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[19]
port 54 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_out[1]
port 55 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[2]
port 56 nsew default tristate
rlabel metal3 s 0 1096 480 1216 6 chanx_left_out[3]
port 57 nsew default tristate
rlabel metal3 s 0 1504 480 1624 6 chanx_left_out[4]
port 58 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[5]
port 59 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[6]
port 60 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 chanx_left_out[7]
port 61 nsew default tristate
rlabel metal3 s 0 2864 480 2984 6 chanx_left_out[8]
port 62 nsew default tristate
rlabel metal3 s 0 3136 480 3256 6 chanx_left_out[9]
port 63 nsew default tristate
rlabel metal3 s 19520 10208 20000 10328 6 chanx_right_in[0]
port 64 nsew default input
rlabel metal3 s 19520 13472 20000 13592 6 chanx_right_in[10]
port 65 nsew default input
rlabel metal3 s 19520 13744 20000 13864 6 chanx_right_in[11]
port 66 nsew default input
rlabel metal3 s 19520 14152 20000 14272 6 chanx_right_in[12]
port 67 nsew default input
rlabel metal3 s 19520 14424 20000 14544 6 chanx_right_in[13]
port 68 nsew default input
rlabel metal3 s 19520 14832 20000 14952 6 chanx_right_in[14]
port 69 nsew default input
rlabel metal3 s 19520 15104 20000 15224 6 chanx_right_in[15]
port 70 nsew default input
rlabel metal3 s 19520 15376 20000 15496 6 chanx_right_in[16]
port 71 nsew default input
rlabel metal3 s 19520 15784 20000 15904 6 chanx_right_in[17]
port 72 nsew default input
rlabel metal3 s 19520 16056 20000 16176 6 chanx_right_in[18]
port 73 nsew default input
rlabel metal3 s 19520 16464 20000 16584 6 chanx_right_in[19]
port 74 nsew default input
rlabel metal3 s 19520 10480 20000 10600 6 chanx_right_in[1]
port 75 nsew default input
rlabel metal3 s 19520 10888 20000 11008 6 chanx_right_in[2]
port 76 nsew default input
rlabel metal3 s 19520 11160 20000 11280 6 chanx_right_in[3]
port 77 nsew default input
rlabel metal3 s 19520 11568 20000 11688 6 chanx_right_in[4]
port 78 nsew default input
rlabel metal3 s 19520 11840 20000 11960 6 chanx_right_in[5]
port 79 nsew default input
rlabel metal3 s 19520 12112 20000 12232 6 chanx_right_in[6]
port 80 nsew default input
rlabel metal3 s 19520 12520 20000 12640 6 chanx_right_in[7]
port 81 nsew default input
rlabel metal3 s 19520 12792 20000 12912 6 chanx_right_in[8]
port 82 nsew default input
rlabel metal3 s 19520 13200 20000 13320 6 chanx_right_in[9]
port 83 nsew default input
rlabel metal3 s 19520 3680 20000 3800 6 chanx_right_out[0]
port 84 nsew default tristate
rlabel metal3 s 19520 6944 20000 7064 6 chanx_right_out[10]
port 85 nsew default tristate
rlabel metal3 s 19520 7216 20000 7336 6 chanx_right_out[11]
port 86 nsew default tristate
rlabel metal3 s 19520 7624 20000 7744 6 chanx_right_out[12]
port 87 nsew default tristate
rlabel metal3 s 19520 7896 20000 8016 6 chanx_right_out[13]
port 88 nsew default tristate
rlabel metal3 s 19520 8304 20000 8424 6 chanx_right_out[14]
port 89 nsew default tristate
rlabel metal3 s 19520 8576 20000 8696 6 chanx_right_out[15]
port 90 nsew default tristate
rlabel metal3 s 19520 8848 20000 8968 6 chanx_right_out[16]
port 91 nsew default tristate
rlabel metal3 s 19520 9256 20000 9376 6 chanx_right_out[17]
port 92 nsew default tristate
rlabel metal3 s 19520 9528 20000 9648 6 chanx_right_out[18]
port 93 nsew default tristate
rlabel metal3 s 19520 9936 20000 10056 6 chanx_right_out[19]
port 94 nsew default tristate
rlabel metal3 s 19520 3952 20000 4072 6 chanx_right_out[1]
port 95 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 chanx_right_out[2]
port 96 nsew default tristate
rlabel metal3 s 19520 4632 20000 4752 6 chanx_right_out[3]
port 97 nsew default tristate
rlabel metal3 s 19520 5040 20000 5160 6 chanx_right_out[4]
port 98 nsew default tristate
rlabel metal3 s 19520 5312 20000 5432 6 chanx_right_out[5]
port 99 nsew default tristate
rlabel metal3 s 19520 5584 20000 5704 6 chanx_right_out[6]
port 100 nsew default tristate
rlabel metal3 s 19520 5992 20000 6112 6 chanx_right_out[7]
port 101 nsew default tristate
rlabel metal3 s 19520 6264 20000 6384 6 chanx_right_out[8]
port 102 nsew default tristate
rlabel metal3 s 19520 6672 20000 6792 6 chanx_right_out[9]
port 103 nsew default tristate
rlabel metal3 s 19520 3408 20000 3528 6 clk_1_E_in
port 104 nsew default input
rlabel metal2 s 8298 16520 8354 17000 6 clk_1_N_out
port 105 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 clk_1_S_out
port 106 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 clk_1_W_in
port 107 nsew default input
rlabel metal3 s 19520 3000 20000 3120 6 clk_2_E_in
port 108 nsew default input
rlabel metal3 s 19520 1368 20000 1488 6 clk_2_E_out
port 109 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 clk_2_W_in
port 110 nsew default input
rlabel metal3 s 0 14696 480 14816 6 clk_2_W_out
port 111 nsew default tristate
rlabel metal3 s 19520 2728 20000 2848 6 clk_3_E_in
port 112 nsew default input
rlabel metal3 s 19520 1096 20000 1216 6 clk_3_E_out
port 113 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 clk_3_W_in
port 114 nsew default input
rlabel metal3 s 0 14424 480 14544 6 clk_3_W_out
port 115 nsew default tristate
rlabel metal2 s 11610 16520 11666 17000 6 prog_clk_0_N_in
port 116 nsew default input
rlabel metal2 s 14922 16520 14978 17000 6 prog_clk_0_W_out
port 117 nsew default tristate
rlabel metal3 s 19520 2320 20000 2440 6 prog_clk_1_E_in
port 118 nsew default input
rlabel metal3 s 19520 688 20000 808 6 prog_clk_1_N_out
port 119 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 prog_clk_1_S_out
port 120 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 prog_clk_1_W_in
port 121 nsew default input
rlabel metal3 s 19520 2048 20000 2168 6 prog_clk_2_E_in
port 122 nsew default input
rlabel metal3 s 19520 416 20000 536 6 prog_clk_2_E_out
port 123 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 prog_clk_2_W_in
port 124 nsew default input
rlabel metal3 s 0 14016 480 14136 6 prog_clk_2_W_out
port 125 nsew default tristate
rlabel metal3 s 19520 1776 20000 1896 6 prog_clk_3_E_in
port 126 nsew default input
rlabel metal3 s 19520 144 20000 264 6 prog_clk_3_E_out
port 127 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 prog_clk_3_W_in
port 128 nsew default input
rlabel metal3 s 0 13744 480 13864 6 prog_clk_3_W_out
port 129 nsew default tristate
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 130 nsew default input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 131 nsew default input
<< properties >>
string FIXED_BBOX 0 0 20000 17000
<< end >>
