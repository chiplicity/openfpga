magic
tech EFS8A
magscale 1 2
timestamp 1603801549
<< locali >>
rect 10885 13787 10919 13889
rect 17601 6103 17635 6409
rect 8953 5015 8987 5321
<< viali >>
rect 1476 24225 1510 24259
rect 1547 24021 1581 24055
rect 2237 23817 2271 23851
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 1547 23477 1581 23511
rect 1476 22525 1510 22559
rect 1869 22525 1903 22559
rect 1547 22389 1581 22423
rect 1476 21437 1510 21471
rect 1869 21437 1903 21471
rect 1547 21301 1581 21335
rect 1444 20961 1478 20995
rect 1547 20757 1581 20791
rect 1593 20553 1627 20587
rect 1476 19873 1510 19907
rect 1547 19669 1581 19703
rect 1593 19465 1627 19499
rect 5952 18785 5986 18819
rect 6055 18581 6089 18615
rect 5917 18377 5951 18411
rect 1476 18173 1510 18207
rect 1869 18173 1903 18207
rect 1547 18037 1581 18071
rect 1444 17697 1478 17731
rect 2488 17697 2522 17731
rect 11196 17697 11230 17731
rect 1547 17561 1581 17595
rect 2145 17493 2179 17527
rect 2559 17493 2593 17527
rect 11299 17493 11333 17527
rect 11161 17289 11195 17323
rect 2145 17085 2179 17119
rect 3652 17085 3686 17119
rect 4077 17085 4111 17119
rect 2053 17017 2087 17051
rect 1593 16949 1627 16983
rect 3065 16949 3099 16983
rect 3755 16949 3789 16983
rect 1961 16609 1995 16643
rect 2053 16609 2087 16643
rect 4128 16609 4162 16643
rect 4215 16609 4249 16643
rect 4905 16065 4939 16099
rect 2421 15997 2455 16031
rect 3985 15997 4019 16031
rect 1777 15861 1811 15895
rect 2237 15861 2271 15895
rect 2605 15861 2639 15895
rect 3709 15861 3743 15895
rect 4169 15861 4203 15895
rect 5457 15861 5491 15895
rect 1961 15521 1995 15555
rect 4629 15521 4663 15555
rect 10368 15521 10402 15555
rect 15612 15521 15646 15555
rect 4537 15453 4571 15487
rect 6101 15453 6135 15487
rect 2145 15317 2179 15351
rect 10471 15317 10505 15351
rect 15715 15317 15749 15351
rect 10609 15113 10643 15147
rect 15577 15113 15611 15147
rect 1869 14909 1903 14943
rect 3249 14909 3283 14943
rect 3985 14909 4019 14943
rect 5089 14909 5123 14943
rect 5549 14909 5583 14943
rect 8192 14909 8226 14943
rect 9848 14909 9882 14943
rect 10241 14909 10275 14943
rect 11228 14909 11262 14943
rect 5825 14841 5859 14875
rect 1685 14773 1719 14807
rect 2237 14773 2271 14807
rect 3617 14773 3651 14807
rect 4629 14773 4663 14807
rect 4997 14773 5031 14807
rect 8263 14773 8297 14807
rect 8677 14773 8711 14807
rect 9919 14773 9953 14807
rect 11299 14773 11333 14807
rect 11713 14773 11747 14807
rect 1476 14433 1510 14467
rect 2237 14433 2271 14467
rect 3065 14433 3099 14467
rect 5457 14433 5491 14467
rect 8652 14433 8686 14467
rect 10517 14433 10551 14467
rect 12081 14433 12115 14467
rect 15612 14433 15646 14467
rect 4353 14365 4387 14399
rect 6929 14365 6963 14399
rect 1869 14297 1903 14331
rect 1547 14229 1581 14263
rect 2881 14229 2915 14263
rect 5181 14229 5215 14263
rect 5641 14229 5675 14263
rect 8723 14229 8757 14263
rect 10701 14229 10735 14263
rect 12265 14229 12299 14263
rect 15715 14229 15749 14263
rect 2605 14025 2639 14059
rect 3801 14025 3835 14059
rect 4261 14025 4295 14059
rect 5457 14025 5491 14059
rect 11069 14025 11103 14059
rect 15577 14025 15611 14059
rect 3249 13957 3283 13991
rect 6285 13957 6319 13991
rect 9229 13957 9263 13991
rect 9735 13957 9769 13991
rect 10793 13957 10827 13991
rect 12633 13957 12667 13991
rect 1501 13889 1535 13923
rect 4445 13889 4479 13923
rect 8539 13889 8573 13923
rect 10885 13889 10919 13923
rect 11437 13889 11471 13923
rect 1593 13821 1627 13855
rect 2973 13821 3007 13855
rect 3065 13821 3099 13855
rect 6653 13821 6687 13855
rect 7113 13821 7147 13855
rect 7389 13821 7423 13855
rect 8436 13821 8470 13855
rect 8953 13821 8987 13855
rect 9664 13821 9698 13855
rect 10057 13821 10091 13855
rect 10609 13821 10643 13855
rect 12081 13821 12115 13855
rect 12449 13821 12483 13855
rect 12909 13821 12943 13855
rect 13496 13821 13530 13855
rect 13599 13821 13633 13855
rect 13921 13821 13955 13855
rect 4537 13753 4571 13787
rect 5089 13753 5123 13787
rect 10885 13753 10919 13787
rect 7113 13685 7147 13719
rect 1593 13481 1627 13515
rect 4215 13481 4249 13515
rect 8769 13481 8803 13515
rect 10793 13481 10827 13515
rect 2145 13413 2179 13447
rect 5549 13413 5583 13447
rect 7113 13413 7147 13447
rect 4144 13345 4178 13379
rect 8585 13345 8619 13379
rect 9689 13345 9723 13379
rect 11805 13345 11839 13379
rect 13001 13345 13035 13379
rect 14013 13345 14047 13379
rect 15428 13345 15462 13379
rect 2053 13277 2087 13311
rect 5457 13277 5491 13311
rect 7021 13277 7055 13311
rect 7297 13277 7331 13311
rect 2605 13209 2639 13243
rect 6009 13209 6043 13243
rect 3065 13141 3099 13175
rect 4905 13141 4939 13175
rect 9873 13141 9907 13175
rect 10425 13141 10459 13175
rect 11713 13141 11747 13175
rect 13185 13141 13219 13175
rect 14197 13141 14231 13175
rect 15531 13141 15565 13175
rect 1685 12937 1719 12971
rect 2053 12937 2087 12971
rect 3341 12937 3375 12971
rect 4169 12937 4203 12971
rect 5825 12937 5859 12971
rect 7113 12937 7147 12971
rect 10498 12937 10532 12971
rect 11805 12937 11839 12971
rect 13461 12937 13495 12971
rect 14473 12937 14507 12971
rect 15853 12937 15887 12971
rect 2973 12869 3007 12903
rect 5457 12869 5491 12903
rect 6561 12869 6595 12903
rect 8677 12869 8711 12903
rect 10609 12869 10643 12903
rect 2421 12801 2455 12835
rect 4905 12801 4939 12835
rect 7481 12801 7515 12835
rect 7941 12801 7975 12835
rect 10701 12801 10735 12835
rect 9137 12733 9171 12767
rect 9689 12733 9723 12767
rect 10057 12733 10091 12767
rect 12265 12733 12299 12767
rect 12541 12733 12575 12767
rect 14013 12733 14047 12767
rect 14841 12733 14875 12767
rect 15060 12733 15094 12767
rect 15485 12733 15519 12767
rect 16072 12733 16106 12767
rect 16497 12733 16531 12767
rect 2513 12665 2547 12699
rect 4721 12665 4755 12699
rect 4997 12665 5031 12699
rect 6193 12665 6227 12699
rect 7665 12665 7699 12699
rect 7757 12665 7791 12699
rect 10333 12665 10367 12699
rect 13185 12665 13219 12699
rect 15163 12665 15197 12699
rect 9321 12597 9355 12631
rect 10977 12597 11011 12631
rect 11437 12597 11471 12631
rect 14197 12597 14231 12631
rect 16175 12597 16209 12631
rect 5917 12393 5951 12427
rect 7665 12393 7699 12427
rect 12633 12393 12667 12427
rect 2145 12325 2179 12359
rect 2697 12325 2731 12359
rect 4905 12325 4939 12359
rect 5359 12325 5393 12359
rect 7066 12325 7100 12359
rect 11621 12325 11655 12359
rect 13185 12325 13219 12359
rect 9781 12257 9815 12291
rect 15393 12257 15427 12291
rect 2053 12189 2087 12223
rect 4997 12189 5031 12223
rect 6745 12189 6779 12223
rect 8493 12189 8527 12223
rect 9689 12189 9723 12223
rect 11529 12189 11563 12223
rect 13093 12189 13127 12223
rect 12081 12121 12115 12155
rect 13645 12121 13679 12155
rect 1685 12053 1719 12087
rect 2973 12053 3007 12087
rect 7941 12053 7975 12087
rect 10793 12053 10827 12087
rect 15761 12053 15795 12087
rect 2053 11849 2087 11883
rect 2329 11849 2363 11883
rect 6101 11849 6135 11883
rect 9781 11849 9815 11883
rect 11529 11849 11563 11883
rect 12679 11849 12713 11883
rect 13553 11849 13587 11883
rect 13921 11849 13955 11883
rect 14473 11849 14507 11883
rect 11805 11781 11839 11815
rect 12817 11781 12851 11815
rect 3065 11713 3099 11747
rect 6653 11713 6687 11747
rect 7849 11713 7883 11747
rect 10333 11713 10367 11747
rect 10793 11713 10827 11747
rect 12909 11713 12943 11747
rect 1409 11645 1443 11679
rect 4813 11645 4847 11679
rect 5733 11645 5767 11679
rect 8585 11645 8619 11679
rect 9321 11645 9355 11679
rect 12541 11645 12575 11679
rect 2789 11577 2823 11611
rect 2881 11577 2915 11611
rect 4721 11577 4755 11611
rect 5175 11577 5209 11611
rect 7205 11577 7239 11611
rect 7297 11577 7331 11611
rect 9413 11577 9447 11611
rect 10425 11577 10459 11611
rect 13277 11577 13311 11611
rect 14565 11577 14599 11611
rect 15117 11577 15151 11611
rect 15669 11577 15703 11611
rect 15761 11577 15795 11611
rect 16313 11577 16347 11611
rect 1593 11509 1627 11543
rect 3709 11509 3743 11543
rect 4261 11509 4295 11543
rect 8125 11509 8159 11543
rect 10149 11509 10183 11543
rect 12265 11509 12299 11543
rect 15485 11509 15519 11543
rect 1547 11305 1581 11339
rect 3433 11305 3467 11339
rect 5733 11305 5767 11339
rect 6377 11305 6411 11339
rect 7481 11305 7515 11339
rect 10701 11305 10735 11339
rect 11345 11305 11379 11339
rect 12817 11305 12851 11339
rect 13093 11305 13127 11339
rect 13553 11305 13587 11339
rect 3157 11237 3191 11271
rect 5175 11237 5209 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 12218 11237 12252 11271
rect 13737 11237 13771 11271
rect 13829 11237 13863 11271
rect 15485 11237 15519 11271
rect 16037 11237 16071 11271
rect 1476 11169 1510 11203
rect 1961 11169 1995 11203
rect 2697 11169 2731 11203
rect 2973 11169 3007 11203
rect 6561 11169 6595 11203
rect 7205 11169 7239 11203
rect 7665 11169 7699 11203
rect 7757 11169 7791 11203
rect 16865 11169 16899 11203
rect 16957 11169 16991 11203
rect 18496 11169 18530 11203
rect 4813 11101 4847 11135
rect 9781 11101 9815 11135
rect 11897 11101 11931 11135
rect 14013 11101 14047 11135
rect 15393 11101 15427 11135
rect 2237 11033 2271 11067
rect 6745 11033 6779 11067
rect 11713 11033 11747 11067
rect 18567 11033 18601 11067
rect 8769 10965 8803 10999
rect 1685 10761 1719 10795
rect 4813 10761 4847 10795
rect 6285 10761 6319 10795
rect 7481 10761 7515 10795
rect 8861 10761 8895 10795
rect 9229 10761 9263 10795
rect 10609 10761 10643 10795
rect 10885 10761 10919 10795
rect 11621 10761 11655 10795
rect 13553 10761 13587 10795
rect 15025 10761 15059 10795
rect 15761 10761 15795 10795
rect 16957 10761 16991 10795
rect 17233 10761 17267 10795
rect 9597 10693 9631 10727
rect 11989 10693 12023 10727
rect 16497 10693 16531 10727
rect 1869 10625 1903 10659
rect 4077 10625 4111 10659
rect 12541 10625 12575 10659
rect 3433 10557 3467 10591
rect 3801 10557 3835 10591
rect 4445 10557 4479 10591
rect 5181 10557 5215 10591
rect 5457 10557 5491 10591
rect 7941 10557 7975 10591
rect 9689 10557 9723 10591
rect 14105 10557 14139 10591
rect 17877 10557 17911 10591
rect 18153 10557 18187 10591
rect 1961 10489 1995 10523
rect 2513 10489 2547 10523
rect 3249 10489 3283 10523
rect 7849 10489 7883 10523
rect 8303 10489 8337 10523
rect 10051 10489 10085 10523
rect 12633 10489 12667 10523
rect 13185 10489 13219 10523
rect 14426 10489 14460 10523
rect 15945 10489 15979 10523
rect 16037 10489 16071 10523
rect 19073 10489 19107 10523
rect 2881 10421 2915 10455
rect 4997 10421 5031 10455
rect 6009 10421 6043 10455
rect 6837 10421 6871 10455
rect 14013 10421 14047 10455
rect 15301 10421 15335 10455
rect 18337 10421 18371 10455
rect 1961 10217 1995 10251
rect 2329 10217 2363 10251
rect 4813 10217 4847 10251
rect 4997 10217 5031 10251
rect 6607 10217 6641 10251
rect 8769 10217 8803 10251
rect 12357 10217 12391 10251
rect 12725 10217 12759 10251
rect 13185 10217 13219 10251
rect 14381 10217 14415 10251
rect 15025 10217 15059 10251
rect 16405 10217 16439 10251
rect 2605 10149 2639 10183
rect 7573 10149 7607 10183
rect 10609 10149 10643 10183
rect 11799 10149 11833 10183
rect 13823 10149 13857 10183
rect 15485 10149 15519 10183
rect 16037 10149 16071 10183
rect 1476 10081 1510 10115
rect 5181 10081 5215 10115
rect 5365 10081 5399 10115
rect 6504 10081 6538 10115
rect 7941 10081 7975 10115
rect 8125 10081 8159 10115
rect 8493 10081 8527 10115
rect 10517 10081 10551 10115
rect 17141 10081 17175 10115
rect 17325 10081 17359 10115
rect 19073 10081 19107 10115
rect 23616 10081 23650 10115
rect 2513 10013 2547 10047
rect 3157 10013 3191 10047
rect 3525 10013 3559 10047
rect 7205 10013 7239 10047
rect 11437 10013 11471 10047
rect 13461 10013 13495 10047
rect 15393 10013 15427 10047
rect 17417 10013 17451 10047
rect 18429 10013 18463 10047
rect 14657 9945 14691 9979
rect 1547 9877 1581 9911
rect 9413 9877 9447 9911
rect 11345 9877 11379 9911
rect 18153 9877 18187 9911
rect 23719 9877 23753 9911
rect 2697 9673 2731 9707
rect 9229 9673 9263 9707
rect 9965 9673 9999 9707
rect 11897 9673 11931 9707
rect 13829 9673 13863 9707
rect 15853 9673 15887 9707
rect 17785 9673 17819 9707
rect 19073 9673 19107 9707
rect 23489 9673 23523 9707
rect 6009 9605 6043 9639
rect 6975 9605 7009 9639
rect 10701 9605 10735 9639
rect 14749 9605 14783 9639
rect 4721 9537 4755 9571
rect 7297 9537 7331 9571
rect 11529 9537 11563 9571
rect 13461 9537 13495 9571
rect 16497 9537 16531 9571
rect 3065 9469 3099 9503
rect 3433 9469 3467 9503
rect 3709 9469 3743 9503
rect 6904 9469 6938 9503
rect 7757 9469 7791 9503
rect 8401 9469 8435 9503
rect 8585 9469 8619 9503
rect 8953 9469 8987 9503
rect 10793 9469 10827 9503
rect 11253 9469 11287 9503
rect 13001 9469 13035 9503
rect 13277 9469 13311 9503
rect 14841 9469 14875 9503
rect 15301 9469 15335 9503
rect 17141 9469 17175 9503
rect 18153 9469 18187 9503
rect 19533 9469 19567 9503
rect 19717 9469 19751 9503
rect 21256 9469 21290 9503
rect 21649 9469 21683 9503
rect 23708 9469 23742 9503
rect 24133 9469 24167 9503
rect 1685 9401 1719 9435
rect 1777 9401 1811 9435
rect 2329 9401 2363 9435
rect 3893 9401 3927 9435
rect 4629 9401 4663 9435
rect 5083 9401 5117 9435
rect 9505 9401 9539 9435
rect 10333 9401 10367 9435
rect 12173 9401 12207 9435
rect 15577 9401 15611 9435
rect 16313 9401 16347 9435
rect 16589 9401 16623 9435
rect 20361 9401 20395 9435
rect 4169 9333 4203 9367
rect 5641 9333 5675 9367
rect 6469 9333 6503 9367
rect 14105 9333 14139 9367
rect 17509 9333 17543 9367
rect 18337 9333 18371 9367
rect 21327 9333 21361 9367
rect 23811 9333 23845 9367
rect 2145 9129 2179 9163
rect 3525 9129 3559 9163
rect 4629 9129 4663 9163
rect 8217 9129 8251 9163
rect 10425 9129 10459 9163
rect 10793 9129 10827 9163
rect 11437 9129 11471 9163
rect 14933 9129 14967 9163
rect 15301 9129 15335 9163
rect 15761 9129 15795 9163
rect 19165 9129 19199 9163
rect 2605 9061 2639 9095
rect 5134 9061 5168 9095
rect 9781 9061 9815 9095
rect 13645 9061 13679 9095
rect 16589 9061 16623 9095
rect 16681 9061 16715 9095
rect 17233 9061 17267 9095
rect 18245 9061 18279 9095
rect 1476 8993 1510 9027
rect 4813 8993 4847 9027
rect 7113 8993 7147 9027
rect 11345 8993 11379 9027
rect 11759 8993 11793 9027
rect 13093 8993 13127 9027
rect 13369 8993 13403 9027
rect 21960 8993 21994 9027
rect 2513 8925 2547 8959
rect 2789 8925 2823 8959
rect 3801 8925 3835 8959
rect 7021 8925 7055 8959
rect 8585 8925 8619 8959
rect 10149 8925 10183 8959
rect 11253 8925 11287 8959
rect 18153 8925 18187 8959
rect 18429 8925 18463 8959
rect 19625 8925 19659 8959
rect 20913 8925 20947 8959
rect 6561 8857 6595 8891
rect 9946 8857 9980 8891
rect 1547 8789 1581 8823
rect 5733 8789 5767 8823
rect 6929 8789 6963 8823
rect 9413 8789 9447 8823
rect 10057 8789 10091 8823
rect 12633 8789 12667 8823
rect 14289 8789 14323 8823
rect 22063 8789 22097 8823
rect 1961 8585 1995 8619
rect 3065 8585 3099 8619
rect 6285 8585 6319 8619
rect 9321 8585 9355 8619
rect 9873 8585 9907 8619
rect 10517 8585 10551 8619
rect 11069 8585 11103 8619
rect 12909 8585 12943 8619
rect 13277 8585 13311 8619
rect 13737 8585 13771 8619
rect 15669 8585 15703 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 18521 8585 18555 8619
rect 20453 8585 20487 8619
rect 10747 8517 10781 8551
rect 10885 8517 10919 8551
rect 12265 8517 12299 8551
rect 12798 8517 12832 8551
rect 16773 8517 16807 8551
rect 17049 8517 17083 8551
rect 18245 8517 18279 8551
rect 19717 8517 19751 8551
rect 21281 8517 21315 8551
rect 2145 8449 2179 8483
rect 3525 8449 3559 8483
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 7389 8449 7423 8483
rect 9045 8449 9079 8483
rect 10977 8449 11011 8483
rect 13001 8449 13035 8483
rect 15853 8449 15887 8483
rect 19165 8449 19199 8483
rect 20729 8449 20763 8483
rect 3893 8381 3927 8415
rect 4169 8381 4203 8415
rect 8309 8381 8343 8415
rect 8677 8381 8711 8415
rect 9137 8381 9171 8415
rect 10609 8381 10643 8415
rect 14105 8381 14139 8415
rect 14197 8381 14231 8415
rect 14657 8381 14691 8415
rect 18061 8381 18095 8415
rect 18889 8381 18923 8415
rect 22236 8381 22270 8415
rect 22661 8381 22695 8415
rect 2237 8313 2271 8347
rect 2789 8313 2823 8347
rect 4353 8313 4387 8347
rect 5365 8313 5399 8347
rect 6653 8313 6687 8347
rect 7297 8313 7331 8347
rect 7710 8313 7744 8347
rect 11805 8313 11839 8347
rect 12633 8313 12667 8347
rect 16174 8313 16208 8347
rect 19257 8313 19291 8347
rect 20821 8313 20855 8347
rect 21925 8313 21959 8347
rect 22339 8313 22373 8347
rect 4905 8245 4939 8279
rect 14289 8245 14323 8279
rect 1685 8041 1719 8075
rect 3157 8041 3191 8075
rect 3709 8041 3743 8075
rect 6009 8041 6043 8075
rect 7757 8041 7791 8075
rect 9505 8041 9539 8075
rect 11989 8041 12023 8075
rect 13553 8041 13587 8075
rect 15853 8041 15887 8075
rect 17601 8041 17635 8075
rect 19073 8041 19107 8075
rect 19349 8041 19383 8075
rect 19717 8041 19751 8075
rect 20729 8041 20763 8075
rect 1869 7973 1903 8007
rect 1961 7973 1995 8007
rect 2789 7973 2823 8007
rect 5083 7973 5117 8007
rect 7205 7973 7239 8007
rect 7573 7973 7607 8007
rect 9965 7973 9999 8007
rect 12173 7973 12207 8007
rect 16681 7973 16715 8007
rect 16773 7973 16807 8007
rect 17325 7973 17359 8007
rect 18474 7973 18508 8007
rect 4721 7905 4755 7939
rect 6469 7905 6503 7939
rect 7941 7905 7975 7939
rect 8217 7905 8251 7939
rect 8493 7905 8527 7939
rect 10609 7905 10643 7939
rect 12817 7905 12851 7939
rect 21005 7905 21039 7939
rect 22477 7905 22511 7939
rect 23556 7905 23590 7939
rect 2513 7837 2547 7871
rect 10517 7837 10551 7871
rect 10977 7837 11011 7871
rect 11713 7837 11747 7871
rect 13737 7837 13771 7871
rect 15301 7837 15335 7871
rect 16497 7837 16531 7871
rect 18153 7837 18187 7871
rect 20913 7837 20947 7871
rect 6653 7769 6687 7803
rect 10747 7769 10781 7803
rect 10885 7769 10919 7803
rect 11069 7769 11103 7803
rect 5641 7701 5675 7735
rect 13185 7701 13219 7735
rect 14289 7701 14323 7735
rect 21925 7701 21959 7735
rect 22661 7701 22695 7735
rect 23627 7701 23661 7735
rect 1869 7497 1903 7531
rect 3525 7497 3559 7531
rect 5917 7497 5951 7531
rect 9045 7497 9079 7531
rect 10701 7497 10735 7531
rect 12265 7497 12299 7531
rect 12725 7497 12759 7531
rect 13369 7497 13403 7531
rect 16865 7497 16899 7531
rect 17417 7497 17451 7531
rect 21446 7497 21480 7531
rect 22293 7497 22327 7531
rect 22661 7497 22695 7531
rect 2789 7429 2823 7463
rect 4629 7429 4663 7463
rect 10333 7429 10367 7463
rect 21557 7429 21591 7463
rect 2237 7361 2271 7395
rect 4721 7361 4755 7395
rect 6285 7361 6319 7395
rect 11161 7361 11195 7395
rect 13737 7361 13771 7395
rect 15485 7361 15519 7395
rect 15945 7361 15979 7395
rect 18797 7361 18831 7395
rect 19073 7361 19107 7395
rect 19809 7361 19843 7395
rect 21097 7361 21131 7395
rect 21741 7361 21775 7395
rect 23489 7361 23523 7395
rect 3760 7293 3794 7327
rect 5641 7293 5675 7327
rect 7113 7293 7147 7327
rect 7481 7293 7515 7327
rect 7849 7293 7883 7327
rect 8217 7293 8251 7327
rect 8401 7293 8435 7327
rect 9540 7293 9574 7327
rect 10793 7293 10827 7327
rect 11529 7293 11563 7327
rect 12633 7293 12667 7327
rect 14105 7293 14139 7327
rect 14289 7293 14323 7327
rect 18061 7293 18095 7327
rect 18521 7293 18555 7327
rect 20453 7293 20487 7327
rect 21281 7293 21315 7327
rect 21620 7293 21654 7327
rect 23673 7293 23707 7327
rect 24133 7293 24167 7327
rect 24720 7293 24754 7327
rect 25145 7293 25179 7327
rect 2329 7225 2363 7259
rect 3249 7225 3283 7259
rect 3847 7225 3881 7259
rect 5083 7225 5117 7259
rect 9413 7225 9447 7259
rect 11897 7225 11931 7259
rect 12449 7225 12483 7259
rect 15853 7225 15887 7259
rect 16307 7225 16341 7259
rect 19901 7225 19935 7259
rect 20821 7225 20855 7259
rect 4169 7157 4203 7191
rect 7665 7157 7699 7191
rect 9643 7157 9677 7191
rect 13921 7157 13955 7191
rect 17877 7157 17911 7191
rect 19625 7157 19659 7191
rect 23857 7157 23891 7191
rect 24823 7157 24857 7191
rect 2605 6953 2639 6987
rect 4813 6953 4847 6987
rect 6469 6953 6503 6987
rect 9413 6953 9447 6987
rect 17509 6953 17543 6987
rect 18153 6953 18187 6987
rect 19533 6953 19567 6987
rect 20729 6953 20763 6987
rect 1777 6885 1811 6919
rect 7113 6885 7147 6919
rect 18934 6885 18968 6919
rect 21097 6885 21131 6919
rect 4077 6817 4111 6851
rect 5181 6817 5215 6851
rect 5641 6817 5675 6851
rect 8033 6817 8067 6851
rect 8544 6817 8578 6851
rect 9689 6817 9723 6851
rect 10333 6817 10367 6851
rect 10885 6817 10919 6851
rect 11621 6817 11655 6851
rect 11897 6817 11931 6851
rect 13093 6817 13127 6851
rect 13645 6817 13679 6851
rect 15301 6817 15335 6851
rect 16313 6817 16347 6851
rect 16865 6817 16899 6851
rect 22477 6817 22511 6851
rect 22569 6817 22603 6851
rect 24041 6817 24075 6851
rect 25212 6817 25246 6851
rect 1685 6749 1719 6783
rect 5733 6749 5767 6783
rect 7021 6749 7055 6783
rect 7389 6749 7423 6783
rect 8631 6749 8665 6783
rect 12817 6749 12851 6783
rect 14013 6749 14047 6783
rect 15669 6749 15703 6783
rect 15761 6749 15795 6783
rect 17233 6749 17267 6783
rect 18613 6749 18647 6783
rect 21005 6749 21039 6783
rect 21281 6749 21315 6783
rect 2237 6681 2271 6715
rect 4261 6681 4295 6715
rect 6837 6681 6871 6715
rect 15577 6681 15611 6715
rect 16681 6681 16715 6715
rect 17141 6681 17175 6715
rect 8401 6613 8435 6647
rect 11529 6613 11563 6647
rect 13553 6613 13587 6647
rect 13783 6613 13817 6647
rect 13921 6613 13955 6647
rect 14289 6613 14323 6647
rect 14749 6613 14783 6647
rect 15466 6613 15500 6647
rect 17030 6613 17064 6647
rect 18429 6613 18463 6647
rect 19901 6613 19935 6647
rect 21925 6613 21959 6647
rect 24225 6613 24259 6647
rect 25283 6613 25317 6647
rect 4905 6409 4939 6443
rect 7205 6409 7239 6443
rect 9781 6409 9815 6443
rect 11713 6409 11747 6443
rect 12725 6409 12759 6443
rect 17601 6409 17635 6443
rect 18521 6409 18555 6443
rect 19073 6409 19107 6443
rect 19441 6409 19475 6443
rect 21005 6409 21039 6443
rect 21354 6409 21388 6443
rect 22937 6409 22971 6443
rect 24133 6409 24167 6443
rect 2605 6341 2639 6375
rect 5917 6341 5951 6375
rect 10333 6341 10367 6375
rect 12265 6341 12299 6375
rect 14289 6341 14323 6375
rect 17417 6341 17451 6375
rect 1593 6273 1627 6307
rect 6653 6273 6687 6307
rect 7297 6273 7331 6307
rect 12596 6273 12630 6307
rect 12817 6273 12851 6307
rect 12909 6273 12943 6307
rect 14381 6273 14415 6307
rect 15301 6273 15335 6307
rect 16497 6273 16531 6307
rect 3341 6205 3375 6239
rect 3709 6205 3743 6239
rect 3985 6205 4019 6239
rect 4169 6205 4203 6239
rect 4997 6205 5031 6239
rect 8493 6205 8527 6239
rect 9080 6205 9114 6239
rect 10425 6205 10459 6239
rect 10977 6205 11011 6239
rect 14160 6205 14194 6239
rect 1685 6137 1719 6171
rect 2237 6137 2271 6171
rect 5318 6137 5352 6171
rect 6285 6137 6319 6171
rect 7618 6137 7652 6171
rect 12449 6137 12483 6171
rect 14013 6137 14047 6171
rect 14749 6137 14783 6171
rect 16313 6137 16347 6171
rect 16589 6137 16623 6171
rect 17141 6137 17175 6171
rect 17877 6341 17911 6375
rect 18337 6341 18371 6375
rect 21465 6341 21499 6375
rect 22293 6341 22327 6375
rect 24869 6341 24903 6375
rect 18429 6273 18463 6307
rect 20177 6273 20211 6307
rect 21557 6273 21591 6307
rect 22569 6273 22603 6307
rect 18208 6205 18242 6239
rect 19625 6205 19659 6239
rect 20085 6205 20119 6239
rect 21189 6205 21223 6239
rect 24685 6205 24719 6239
rect 25145 6205 25179 6239
rect 18061 6137 18095 6171
rect 2973 6069 3007 6103
rect 4445 6069 4479 6103
rect 8217 6069 8251 6103
rect 8861 6069 8895 6103
rect 9183 6069 9217 6103
rect 10701 6069 10735 6103
rect 13737 6069 13771 6103
rect 15761 6069 15795 6103
rect 17601 6069 17635 6103
rect 21833 6069 21867 6103
rect 23673 6069 23707 6103
rect 25513 6069 25547 6103
rect 1593 5865 1627 5899
rect 2973 5865 3007 5899
rect 3525 5865 3559 5899
rect 4261 5865 4295 5899
rect 4721 5865 4755 5899
rect 5825 5865 5859 5899
rect 7113 5865 7147 5899
rect 7757 5865 7791 5899
rect 12541 5865 12575 5899
rect 14473 5865 14507 5899
rect 14841 5865 14875 5899
rect 15485 5865 15519 5899
rect 15853 5865 15887 5899
rect 17049 5865 17083 5899
rect 18153 5865 18187 5899
rect 19625 5865 19659 5899
rect 20729 5865 20763 5899
rect 22017 5865 22051 5899
rect 22569 5865 22603 5899
rect 2145 5797 2179 5831
rect 5226 5797 5260 5831
rect 9873 5797 9907 5831
rect 11253 5797 11287 5831
rect 16491 5797 16525 5831
rect 17417 5797 17451 5831
rect 18678 5797 18712 5831
rect 4905 5729 4939 5763
rect 6720 5729 6754 5763
rect 7665 5729 7699 5763
rect 8125 5729 8159 5763
rect 12817 5729 12851 5763
rect 16129 5729 16163 5763
rect 20913 5729 20947 5763
rect 21465 5729 21499 5763
rect 22477 5729 22511 5763
rect 22937 5729 22971 5763
rect 24041 5729 24075 5763
rect 25145 5729 25179 5763
rect 2053 5661 2087 5695
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 11161 5661 11195 5695
rect 11400 5661 11434 5695
rect 11621 5661 11655 5695
rect 13185 5661 13219 5695
rect 14013 5661 14047 5695
rect 17785 5661 17819 5695
rect 18337 5661 18371 5695
rect 21373 5661 21407 5695
rect 2605 5593 2639 5627
rect 10793 5593 10827 5627
rect 13277 5593 13311 5627
rect 25329 5593 25363 5627
rect 6791 5525 6825 5559
rect 7481 5525 7515 5559
rect 11529 5525 11563 5559
rect 11713 5525 11747 5559
rect 12955 5525 12989 5559
rect 13093 5525 13127 5559
rect 19257 5525 19291 5559
rect 19993 5525 20027 5559
rect 24225 5525 24259 5559
rect 2789 5321 2823 5355
rect 4997 5321 5031 5355
rect 6561 5321 6595 5355
rect 7389 5321 7423 5355
rect 8769 5321 8803 5355
rect 8953 5321 8987 5355
rect 11023 5321 11057 5355
rect 11437 5321 11471 5355
rect 12081 5321 12115 5355
rect 15025 5321 15059 5355
rect 15485 5321 15519 5355
rect 16221 5321 16255 5355
rect 18613 5321 18647 5355
rect 20453 5321 20487 5355
rect 22109 5321 22143 5355
rect 22477 5321 22511 5355
rect 24685 5321 24719 5355
rect 25145 5321 25179 5355
rect 1869 5185 1903 5219
rect 2329 5185 2363 5219
rect 3525 5185 3559 5219
rect 5917 5185 5951 5219
rect 7573 5185 7607 5219
rect 3893 5117 3927 5151
rect 4169 5117 4203 5151
rect 5457 5117 5491 5151
rect 5733 5117 5767 5151
rect 1961 5049 1995 5083
rect 6285 5049 6319 5083
rect 7894 5049 7928 5083
rect 18889 5253 18923 5287
rect 20085 5253 20119 5287
rect 23029 5253 23063 5287
rect 25421 5253 25455 5287
rect 9137 5185 9171 5219
rect 9689 5185 9723 5219
rect 10793 5185 10827 5219
rect 16497 5185 16531 5219
rect 17141 5185 17175 5219
rect 19533 5185 19567 5219
rect 21097 5185 21131 5219
rect 21741 5185 21775 5219
rect 10952 5117 10986 5151
rect 11713 5117 11747 5151
rect 12449 5117 12483 5151
rect 12909 5117 12943 5151
rect 14197 5117 14231 5151
rect 14565 5117 14599 5151
rect 23765 5117 23799 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 9413 5049 9447 5083
rect 9505 5049 9539 5083
rect 10425 5049 10459 5083
rect 13185 5049 13219 5083
rect 13921 5049 13955 5083
rect 14749 5049 14783 5083
rect 15853 5049 15887 5083
rect 16589 5049 16623 5083
rect 19349 5049 19383 5083
rect 19625 5049 19659 5083
rect 21189 5049 21223 5083
rect 23673 5049 23707 5083
rect 1685 4981 1719 5015
rect 3893 4981 3927 5015
rect 7021 4981 7055 5015
rect 8493 4981 8527 5015
rect 8953 4981 8987 5015
rect 13461 4981 13495 5015
rect 18061 4981 18095 5015
rect 20913 4981 20947 5015
rect 22569 4981 22603 5015
rect 23489 4981 23523 5015
rect 1869 4777 1903 4811
rect 3249 4777 3283 4811
rect 3709 4777 3743 4811
rect 4721 4777 4755 4811
rect 5641 4777 5675 4811
rect 9321 4777 9355 4811
rect 9965 4777 9999 4811
rect 11345 4777 11379 4811
rect 12909 4777 12943 4811
rect 14381 4777 14415 4811
rect 16405 4777 16439 4811
rect 16773 4777 16807 4811
rect 18429 4777 18463 4811
rect 19809 4777 19843 4811
rect 20729 4777 20763 4811
rect 2421 4709 2455 4743
rect 6377 4709 6411 4743
rect 7941 4709 7975 4743
rect 10419 4709 10453 4743
rect 11621 4709 11655 4743
rect 17141 4709 17175 4743
rect 19210 4709 19244 4743
rect 21097 4709 21131 4743
rect 4629 4641 4663 4675
rect 5181 4641 5215 4675
rect 10057 4641 10091 4675
rect 11805 4641 11839 4675
rect 14013 4641 14047 4675
rect 15301 4641 15335 4675
rect 15853 4641 15887 4675
rect 18889 4641 18923 4675
rect 22661 4641 22695 4675
rect 24685 4641 24719 4675
rect 2329 4573 2363 4607
rect 2973 4573 3007 4607
rect 6285 4573 6319 4607
rect 6929 4573 6963 4607
rect 7297 4573 7331 4607
rect 7849 4573 7883 4607
rect 8493 4573 8527 4607
rect 12173 4573 12207 4607
rect 13369 4573 13403 4607
rect 17049 4573 17083 4607
rect 17325 4573 17359 4607
rect 21005 4573 21039 4607
rect 21649 4573 21683 4607
rect 22477 4573 22511 4607
rect 10977 4505 11011 4539
rect 15393 4505 15427 4539
rect 7665 4437 7699 4471
rect 11943 4437 11977 4471
rect 12081 4437 12115 4471
rect 12449 4437 12483 4471
rect 13185 4437 13219 4471
rect 14841 4437 14875 4471
rect 24317 4437 24351 4471
rect 2237 4233 2271 4267
rect 3893 4233 3927 4267
rect 4353 4233 4387 4267
rect 4721 4233 4755 4267
rect 6285 4233 6319 4267
rect 6561 4233 6595 4267
rect 7573 4233 7607 4267
rect 10977 4233 11011 4267
rect 19073 4233 19107 4267
rect 21649 4233 21683 4267
rect 22753 4233 22787 4267
rect 2421 4097 2455 4131
rect 3065 4097 3099 4131
rect 4813 4097 4847 4131
rect 7297 4097 7331 4131
rect 7757 4097 7791 4131
rect 9045 4097 9079 4131
rect 9597 4097 9631 4131
rect 9873 4097 9907 4131
rect 12725 4097 12759 4131
rect 14013 4097 14047 4131
rect 19441 4097 19475 4131
rect 20085 4097 20119 4131
rect 21373 4097 21407 4131
rect 22109 4097 22143 4131
rect 10609 4029 10643 4063
rect 11136 4029 11170 4063
rect 11529 4029 11563 4063
rect 15117 4029 15151 4063
rect 15301 4029 15335 4063
rect 16221 4029 16255 4063
rect 16405 4029 16439 4063
rect 16865 4029 16899 4063
rect 17785 4029 17819 4063
rect 18061 4029 18095 4063
rect 18521 4029 18555 4063
rect 22201 4029 22235 4063
rect 23765 4029 23799 4063
rect 25237 4029 25271 4063
rect 25789 4029 25823 4063
rect 2513 3961 2547 3995
rect 3341 3961 3375 3995
rect 5134 3961 5168 3995
rect 8078 3961 8112 3995
rect 9413 3961 9447 3995
rect 9689 3961 9723 3995
rect 12265 3961 12299 3995
rect 12817 3961 12851 3995
rect 13369 3961 13403 3995
rect 15577 3961 15611 3995
rect 17141 3961 17175 3995
rect 20729 3961 20763 3995
rect 20821 3961 20855 3995
rect 1869 3893 1903 3927
rect 5733 3893 5767 3927
rect 8677 3893 8711 3927
rect 11207 3893 11241 3927
rect 13737 3893 13771 3927
rect 14749 3893 14783 3927
rect 15853 3893 15887 3927
rect 17509 3893 17543 3927
rect 18153 3893 18187 3927
rect 19625 3893 19659 3927
rect 20545 3893 20579 3927
rect 22385 3893 22419 3927
rect 23489 3893 23523 3927
rect 23949 3893 23983 3927
rect 24685 3893 24719 3927
rect 25421 3893 25455 3927
rect 2329 3689 2363 3723
rect 4721 3689 4755 3723
rect 6101 3689 6135 3723
rect 10149 3689 10183 3723
rect 11989 3689 12023 3723
rect 12449 3689 12483 3723
rect 12817 3689 12851 3723
rect 13277 3689 13311 3723
rect 14289 3689 14323 3723
rect 15669 3689 15703 3723
rect 17049 3689 17083 3723
rect 17693 3689 17727 3723
rect 19349 3689 19383 3723
rect 20729 3689 20763 3723
rect 24317 3689 24351 3723
rect 1961 3621 1995 3655
rect 2513 3621 2547 3655
rect 2605 3621 2639 3655
rect 5134 3621 5168 3655
rect 6469 3621 6503 3655
rect 6653 3621 6687 3655
rect 6745 3621 6779 3655
rect 9827 3621 9861 3655
rect 10517 3621 10551 3655
rect 11134 3621 11168 3655
rect 13731 3621 13765 3655
rect 14933 3621 14967 3655
rect 16102 3621 16136 3655
rect 18153 3621 18187 3655
rect 18791 3621 18825 3655
rect 20913 3621 20947 3655
rect 1476 3553 1510 3587
rect 4813 3553 4847 3587
rect 8125 3553 8159 3587
rect 9724 3553 9758 3587
rect 10793 3553 10827 3587
rect 13369 3553 13403 3587
rect 18429 3553 18463 3587
rect 21005 3553 21039 3587
rect 22569 3553 22603 3587
rect 24133 3553 24167 3587
rect 3433 3485 3467 3519
rect 7297 3485 7331 3519
rect 7849 3485 7883 3519
rect 15761 3485 15795 3519
rect 22477 3485 22511 3519
rect 3065 3417 3099 3451
rect 5733 3417 5767 3451
rect 11713 3417 11747 3451
rect 1547 3349 1581 3383
rect 3893 3349 3927 3383
rect 4261 3349 4295 3383
rect 8309 3349 8343 3383
rect 16681 3349 16715 3383
rect 17325 3349 17359 3383
rect 19625 3349 19659 3383
rect 3249 3145 3283 3179
rect 5181 3145 5215 3179
rect 5549 3145 5583 3179
rect 9965 3145 9999 3179
rect 11897 3145 11931 3179
rect 12265 3145 12299 3179
rect 15025 3145 15059 3179
rect 15669 3145 15703 3179
rect 17417 3145 17451 3179
rect 19073 3145 19107 3179
rect 19533 3145 19567 3179
rect 20637 3145 20671 3179
rect 22569 3145 22603 3179
rect 23489 3145 23523 3179
rect 24685 3145 24719 3179
rect 4905 3077 4939 3111
rect 11069 3077 11103 3111
rect 16129 3077 16163 3111
rect 25421 3077 25455 3111
rect 2973 3009 3007 3043
rect 3893 3009 3927 3043
rect 7941 3009 7975 3043
rect 8493 3009 8527 3043
rect 8769 3009 8803 3043
rect 9505 3009 9539 3043
rect 10517 3009 10551 3043
rect 13001 3009 13035 3043
rect 13829 3009 13863 3043
rect 16221 3009 16255 3043
rect 18153 3009 18187 3043
rect 18797 3009 18831 3043
rect 19717 3009 19751 3043
rect 21281 3009 21315 3043
rect 5365 2941 5399 2975
rect 6285 2941 6319 2975
rect 6653 2941 6687 2975
rect 7481 2941 7515 2975
rect 12449 2941 12483 2975
rect 12633 2941 12667 2975
rect 13277 2941 13311 2975
rect 14749 2941 14783 2975
rect 17141 2941 17175 2975
rect 23765 2941 23799 2975
rect 25237 2941 25271 2975
rect 25789 2941 25823 2975
rect 1777 2873 1811 2907
rect 2329 2873 2363 2907
rect 2421 2873 2455 2907
rect 3709 2873 3743 2907
rect 3985 2873 4019 2907
rect 4537 2873 4571 2907
rect 8309 2873 8343 2907
rect 8585 2873 8619 2907
rect 10609 2873 10643 2907
rect 13737 2873 13771 2907
rect 14191 2873 14225 2907
rect 16542 2873 16576 2907
rect 18245 2873 18279 2907
rect 19809 2873 19843 2907
rect 20361 2873 20395 2907
rect 21097 2873 21131 2907
rect 21373 2873 21407 2907
rect 21925 2873 21959 2907
rect 23673 2873 23707 2907
rect 2145 2805 2179 2839
rect 7113 2805 7147 2839
rect 10333 2805 10367 2839
rect 11529 2805 11563 2839
rect 17877 2805 17911 2839
rect 2329 2601 2363 2635
rect 5365 2601 5399 2635
rect 5825 2601 5859 2635
rect 8125 2601 8159 2635
rect 9137 2601 9171 2635
rect 9505 2601 9539 2635
rect 13829 2601 13863 2635
rect 18153 2601 18187 2635
rect 19809 2601 19843 2635
rect 21005 2601 21039 2635
rect 23397 2601 23431 2635
rect 2605 2533 2639 2567
rect 3157 2533 3191 2567
rect 3893 2533 3927 2567
rect 4261 2533 4295 2567
rect 6745 2533 6779 2567
rect 7113 2533 7147 2567
rect 10425 2533 10459 2567
rect 10517 2533 10551 2567
rect 12449 2533 12483 2567
rect 12909 2533 12943 2567
rect 13461 2533 13495 2567
rect 15623 2533 15657 2567
rect 16405 2533 16439 2567
rect 16681 2533 16715 2567
rect 17233 2533 17267 2567
rect 17785 2533 17819 2567
rect 18429 2533 18463 2567
rect 18521 2533 18555 2567
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 5641 2465 5675 2499
rect 8493 2465 8527 2499
rect 14324 2465 14358 2499
rect 14749 2465 14783 2499
rect 15520 2465 15554 2499
rect 15945 2465 15979 2499
rect 19901 2465 19935 2499
rect 21281 2465 21315 2499
rect 22753 2465 22787 2499
rect 23857 2465 23891 2499
rect 24133 2465 24167 2499
rect 2513 2397 2547 2431
rect 3525 2397 3559 2431
rect 4169 2397 4203 2431
rect 4537 2397 4571 2431
rect 7021 2397 7055 2431
rect 7297 2397 7331 2431
rect 11989 2397 12023 2431
rect 12817 2397 12851 2431
rect 16589 2397 16623 2431
rect 18797 2397 18831 2431
rect 21189 2397 21223 2431
rect 24041 2397 24075 2431
rect 25605 2397 25639 2431
rect 1547 2329 1581 2363
rect 6285 2329 6319 2363
rect 10977 2329 11011 2363
rect 20085 2329 20119 2363
rect 8677 2261 8711 2295
rect 10241 2261 10275 2295
rect 14427 2261 14461 2295
rect 15301 2261 15335 2295
rect 20545 2261 20579 2295
rect 22937 2261 22971 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1486 24265 1492 24268
rect 1464 24259 1492 24265
rect 1464 24225 1476 24259
rect 1464 24219 1492 24225
rect 1486 24216 1492 24219
rect 1544 24216 1550 24268
rect 1535 24055 1593 24061
rect 1535 24021 1547 24055
rect 1581 24052 1593 24055
rect 1762 24052 1768 24064
rect 1581 24024 1768 24052
rect 1581 24021 1593 24024
rect 1535 24015 1593 24021
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1486 23808 1492 23860
rect 1544 23848 1550 23860
rect 2225 23851 2283 23857
rect 2225 23848 2237 23851
rect 1544 23820 2237 23848
rect 1544 23808 1550 23820
rect 2225 23817 2237 23820
rect 2271 23817 2283 23851
rect 2225 23811 2283 23817
rect 1394 23604 1400 23656
rect 1452 23653 1458 23656
rect 1452 23647 1490 23653
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1452 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 1452 23604 1458 23607
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1854 23508 1860 23520
rect 1581 23480 1860 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1854 23468 1860 23480
rect 1912 23468 1918 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1464 22559 1522 22565
rect 1464 22525 1476 22559
rect 1510 22556 1522 22559
rect 1578 22556 1584 22568
rect 1510 22528 1584 22556
rect 1510 22525 1522 22528
rect 1464 22519 1522 22525
rect 1578 22516 1584 22528
rect 1636 22556 1642 22568
rect 1857 22559 1915 22565
rect 1857 22556 1869 22559
rect 1636 22528 1869 22556
rect 1636 22516 1642 22528
rect 1857 22525 1869 22528
rect 1903 22525 1915 22559
rect 1857 22519 1915 22525
rect 1535 22423 1593 22429
rect 1535 22389 1547 22423
rect 1581 22420 1593 22423
rect 2498 22420 2504 22432
rect 1581 22392 2504 22420
rect 1581 22389 1593 22392
rect 1535 22383 1593 22389
rect 2498 22380 2504 22392
rect 2556 22380 2562 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21477 1492 21480
rect 1464 21471 1492 21477
rect 1464 21437 1476 21471
rect 1544 21468 1550 21480
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1544 21440 1869 21468
rect 1464 21431 1492 21437
rect 1486 21428 1492 21431
rect 1544 21428 1550 21440
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 1578 21341 1584 21344
rect 1535 21335 1584 21341
rect 1535 21301 1547 21335
rect 1581 21301 1584 21335
rect 1535 21295 1584 21301
rect 1578 21292 1584 21295
rect 1636 21292 1642 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1394 20952 1400 21004
rect 1452 21001 1458 21004
rect 1452 20995 1490 21001
rect 1478 20961 1490 20995
rect 1452 20955 1490 20961
rect 1452 20952 1458 20955
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 1670 20788 1676 20800
rect 1581 20760 1676 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 1670 20748 1676 20760
rect 1728 20748 1734 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1394 20544 1400 20596
rect 1452 20584 1458 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1452 20556 1593 20584
rect 1452 20544 1458 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1486 19913 1492 19916
rect 1464 19907 1492 19913
rect 1464 19873 1476 19907
rect 1464 19867 1492 19873
rect 1486 19864 1492 19867
rect 1544 19864 1550 19916
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 2590 19700 2596 19712
rect 1581 19672 2596 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 1581 19499 1639 19505
rect 1581 19496 1593 19499
rect 1544 19468 1593 19496
rect 1544 19456 1550 19468
rect 1581 19465 1593 19468
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 3326 19360 3332 19372
rect 2004 19332 3332 19360
rect 2004 19320 2010 19332
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 5534 18776 5540 18828
rect 5592 18816 5598 18828
rect 5940 18819 5998 18825
rect 5940 18816 5952 18819
rect 5592 18788 5952 18816
rect 5592 18776 5598 18788
rect 5940 18785 5952 18788
rect 5986 18785 5998 18819
rect 5940 18779 5998 18785
rect 6043 18615 6101 18621
rect 6043 18581 6055 18615
rect 6089 18612 6101 18615
rect 6270 18612 6276 18624
rect 6089 18584 6276 18612
rect 6089 18581 6101 18584
rect 6043 18575 6101 18581
rect 6270 18572 6276 18584
rect 6328 18572 6334 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 5534 18368 5540 18420
rect 5592 18408 5598 18420
rect 5905 18411 5963 18417
rect 5905 18408 5917 18411
rect 5592 18380 5917 18408
rect 5592 18368 5598 18380
rect 5905 18377 5917 18380
rect 5951 18377 5963 18411
rect 5905 18371 5963 18377
rect 1464 18207 1522 18213
rect 1464 18173 1476 18207
rect 1510 18204 1522 18207
rect 1578 18204 1584 18216
rect 1510 18176 1584 18204
rect 1510 18173 1522 18176
rect 1464 18167 1522 18173
rect 1578 18164 1584 18176
rect 1636 18204 1642 18216
rect 1857 18207 1915 18213
rect 1857 18204 1869 18207
rect 1636 18176 1869 18204
rect 1636 18164 1642 18176
rect 1857 18173 1869 18176
rect 1903 18173 1915 18207
rect 1857 18167 1915 18173
rect 1486 18028 1492 18080
rect 1544 18077 1550 18080
rect 1544 18071 1593 18077
rect 1544 18037 1547 18071
rect 1581 18037 1593 18071
rect 1544 18031 1593 18037
rect 1544 18028 1550 18031
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1394 17688 1400 17740
rect 1452 17737 1458 17740
rect 1452 17731 1490 17737
rect 1478 17697 1490 17731
rect 1452 17691 1490 17697
rect 2476 17731 2534 17737
rect 2476 17697 2488 17731
rect 2522 17728 2534 17731
rect 2958 17728 2964 17740
rect 2522 17700 2964 17728
rect 2522 17697 2534 17700
rect 2476 17691 2534 17697
rect 1452 17688 1458 17691
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 11146 17688 11152 17740
rect 11204 17737 11210 17740
rect 11204 17731 11242 17737
rect 11230 17697 11242 17731
rect 11204 17691 11242 17697
rect 11204 17688 11210 17691
rect 1535 17595 1593 17601
rect 1535 17561 1547 17595
rect 1581 17592 1593 17595
rect 2406 17592 2412 17604
rect 1581 17564 2412 17592
rect 1581 17561 1593 17564
rect 1535 17555 1593 17561
rect 2406 17552 2412 17564
rect 2464 17552 2470 17604
rect 2130 17524 2136 17536
rect 2091 17496 2136 17524
rect 2130 17484 2136 17496
rect 2188 17484 2194 17536
rect 2590 17533 2596 17536
rect 2547 17527 2596 17533
rect 2547 17493 2559 17527
rect 2593 17493 2596 17527
rect 2547 17487 2596 17493
rect 2590 17484 2596 17487
rect 2648 17484 2654 17536
rect 11287 17527 11345 17533
rect 11287 17493 11299 17527
rect 11333 17524 11345 17527
rect 12158 17524 12164 17536
rect 11333 17496 12164 17524
rect 11333 17493 11345 17496
rect 11287 17487 11345 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 11146 17320 11152 17332
rect 11107 17292 11152 17320
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 2130 17116 2136 17128
rect 2091 17088 2136 17116
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 3510 17076 3516 17128
rect 3568 17116 3574 17128
rect 3640 17119 3698 17125
rect 3640 17116 3652 17119
rect 3568 17088 3652 17116
rect 3568 17076 3574 17088
rect 3640 17085 3652 17088
rect 3686 17116 3698 17119
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 3686 17088 4077 17116
rect 3686 17085 3698 17088
rect 3640 17079 3698 17085
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 2038 17048 2044 17060
rect 1999 17020 2044 17048
rect 2038 17008 2044 17020
rect 2096 17008 2102 17060
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1452 16952 1593 16980
rect 1452 16940 1458 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3053 16983 3111 16989
rect 3053 16980 3065 16983
rect 3016 16952 3065 16980
rect 3016 16940 3022 16952
rect 3053 16949 3065 16952
rect 3099 16949 3111 16983
rect 3053 16943 3111 16949
rect 3234 16940 3240 16992
rect 3292 16980 3298 16992
rect 3743 16983 3801 16989
rect 3743 16980 3755 16983
rect 3292 16952 3755 16980
rect 3292 16940 3298 16952
rect 3743 16949 3755 16952
rect 3789 16949 3801 16983
rect 3743 16943 3801 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3878 16668 3884 16720
rect 3936 16708 3942 16720
rect 3936 16680 4154 16708
rect 3936 16668 3942 16680
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 4126 16649 4154 16680
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16609 2099 16643
rect 2041 16603 2099 16609
rect 4116 16643 4174 16649
rect 4116 16609 4128 16643
rect 4162 16609 4174 16643
rect 4116 16603 4174 16609
rect 4203 16643 4261 16649
rect 4203 16609 4215 16643
rect 4249 16640 4261 16643
rect 4338 16640 4344 16652
rect 4249 16612 4344 16640
rect 4249 16609 4261 16612
rect 4203 16603 4261 16609
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 2056 16572 2084 16603
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 1728 16544 2084 16572
rect 1728 16532 1734 16544
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 4893 16099 4951 16105
rect 4893 16096 4905 16099
rect 3936 16068 4905 16096
rect 3936 16056 3942 16068
rect 4893 16065 4905 16068
rect 4939 16065 4951 16099
rect 4893 16059 4951 16065
rect 2409 16031 2467 16037
rect 2409 16028 2421 16031
rect 2240 16000 2421 16028
rect 2240 15904 2268 16000
rect 2409 15997 2421 16000
rect 2455 15997 2467 16031
rect 2409 15991 2467 15997
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 1765 15895 1823 15901
rect 1765 15892 1777 15895
rect 1728 15864 1777 15892
rect 1728 15852 1734 15864
rect 1765 15861 1777 15864
rect 1811 15861 1823 15895
rect 2222 15892 2228 15904
rect 2183 15864 2228 15892
rect 1765 15855 1823 15861
rect 2222 15852 2228 15864
rect 2280 15852 2286 15904
rect 2590 15892 2596 15904
rect 2551 15864 2596 15892
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 3697 15895 3755 15901
rect 3697 15892 3709 15895
rect 3476 15864 3709 15892
rect 3476 15852 3482 15864
rect 3697 15861 3709 15864
rect 3743 15892 3755 15895
rect 3988 15892 4016 15991
rect 3743 15864 4016 15892
rect 4157 15895 4215 15901
rect 3743 15861 3755 15864
rect 3697 15855 3755 15861
rect 4157 15861 4169 15895
rect 4203 15892 4215 15895
rect 4246 15892 4252 15904
rect 4203 15864 4252 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5445 15895 5503 15901
rect 5445 15892 5457 15895
rect 5040 15864 5457 15892
rect 5040 15852 5046 15864
rect 5445 15861 5457 15864
rect 5491 15861 5503 15895
rect 5445 15855 5503 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1210 15648 1216 15700
rect 1268 15688 1274 15700
rect 1854 15688 1860 15700
rect 1268 15660 1860 15688
rect 1268 15648 1274 15660
rect 1854 15648 1860 15660
rect 1912 15648 1918 15700
rect 1854 15512 1860 15564
rect 1912 15552 1918 15564
rect 1949 15555 2007 15561
rect 1949 15552 1961 15555
rect 1912 15524 1961 15552
rect 1912 15512 1918 15524
rect 1949 15521 1961 15524
rect 1995 15521 2007 15555
rect 4614 15552 4620 15564
rect 4575 15524 4620 15552
rect 1949 15515 2007 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 10356 15555 10414 15561
rect 10356 15552 10368 15555
rect 10192 15524 10368 15552
rect 10192 15512 10198 15524
rect 10356 15521 10368 15524
rect 10402 15521 10414 15555
rect 10356 15515 10414 15521
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 15600 15555 15658 15561
rect 15600 15552 15612 15555
rect 15528 15524 15612 15552
rect 15528 15512 15534 15524
rect 15600 15521 15612 15524
rect 15646 15521 15658 15555
rect 15600 15515 15658 15521
rect 4522 15484 4528 15496
rect 4483 15456 4528 15484
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15484 6147 15487
rect 6178 15484 6184 15496
rect 6135 15456 6184 15484
rect 6135 15453 6147 15456
rect 6089 15447 6147 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 2130 15348 2136 15360
rect 2091 15320 2136 15348
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 10459 15351 10517 15357
rect 10459 15317 10471 15351
rect 10505 15348 10517 15351
rect 10686 15348 10692 15360
rect 10505 15320 10692 15348
rect 10505 15317 10517 15320
rect 10459 15311 10517 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 15703 15351 15761 15357
rect 15703 15317 15715 15351
rect 15749 15348 15761 15351
rect 16298 15348 16304 15360
rect 15749 15320 16304 15348
rect 15749 15317 15761 15320
rect 15703 15311 15761 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 10192 15116 10609 15144
rect 10192 15104 10198 15116
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 10597 15107 10655 15113
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15528 15116 15577 15144
rect 15528 15104 15534 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 1857 14943 1915 14949
rect 1857 14940 1869 14943
rect 1452 14912 1869 14940
rect 1452 14900 1458 14912
rect 1857 14909 1869 14912
rect 1903 14909 1915 14943
rect 1857 14903 1915 14909
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14940 3295 14943
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3283 14912 3985 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 3973 14909 3985 14912
rect 4019 14940 4031 14943
rect 4062 14940 4068 14952
rect 4019 14912 4068 14940
rect 4019 14909 4031 14912
rect 3973 14903 4031 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14909 5135 14943
rect 5077 14903 5135 14909
rect 5092 14816 5120 14903
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 5537 14943 5595 14949
rect 5537 14940 5549 14943
rect 5316 14912 5549 14940
rect 5316 14900 5322 14912
rect 5537 14909 5549 14912
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 8180 14943 8238 14949
rect 8180 14909 8192 14943
rect 8226 14940 8238 14943
rect 9836 14943 9894 14949
rect 8226 14912 8708 14940
rect 8226 14909 8238 14912
rect 8180 14903 8238 14909
rect 5813 14875 5871 14881
rect 5813 14841 5825 14875
rect 5859 14872 5871 14875
rect 6086 14872 6092 14884
rect 5859 14844 6092 14872
rect 5859 14841 5871 14844
rect 5813 14835 5871 14841
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 1854 14804 1860 14816
rect 1719 14776 1860 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 2222 14804 2228 14816
rect 2183 14776 2228 14804
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5074 14804 5080 14816
rect 5031 14776 5080 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 8018 14764 8024 14816
rect 8076 14804 8082 14816
rect 8680 14813 8708 14912
rect 9836 14909 9848 14943
rect 9882 14940 9894 14943
rect 9950 14940 9956 14952
rect 9882 14912 9956 14940
rect 9882 14909 9894 14912
rect 9836 14903 9894 14909
rect 9950 14900 9956 14912
rect 10008 14940 10014 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10008 14912 10241 14940
rect 10008 14900 10014 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 11216 14943 11274 14949
rect 11216 14909 11228 14943
rect 11262 14940 11274 14943
rect 11262 14912 11744 14940
rect 11262 14909 11274 14912
rect 11216 14903 11274 14909
rect 8251 14807 8309 14813
rect 8251 14804 8263 14807
rect 8076 14776 8263 14804
rect 8076 14764 8082 14776
rect 8251 14773 8263 14776
rect 8297 14773 8309 14807
rect 8251 14767 8309 14773
rect 8665 14807 8723 14813
rect 8665 14773 8677 14807
rect 8711 14804 8723 14807
rect 9122 14804 9128 14816
rect 8711 14776 9128 14804
rect 8711 14773 8723 14776
rect 8665 14767 8723 14773
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9907 14807 9965 14813
rect 9907 14773 9919 14807
rect 9953 14804 9965 14807
rect 10134 14804 10140 14816
rect 9953 14776 10140 14804
rect 9953 14773 9965 14776
rect 9907 14767 9965 14773
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 11287 14807 11345 14813
rect 11287 14773 11299 14807
rect 11333 14804 11345 14807
rect 11514 14804 11520 14816
rect 11333 14776 11520 14804
rect 11333 14773 11345 14776
rect 11287 14767 11345 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 11716 14813 11744 14912
rect 11701 14807 11759 14813
rect 11701 14773 11713 14807
rect 11747 14804 11759 14807
rect 12342 14804 12348 14816
rect 11747 14776 12348 14804
rect 11747 14773 11759 14776
rect 11701 14767 11759 14773
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1464 14467 1522 14473
rect 1464 14433 1476 14467
rect 1510 14464 1522 14467
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 1510 14436 2237 14464
rect 1510 14433 1522 14436
rect 1464 14427 1522 14433
rect 2225 14433 2237 14436
rect 2271 14464 2283 14467
rect 2682 14464 2688 14476
rect 2271 14436 2688 14464
rect 2271 14433 2283 14436
rect 2225 14427 2283 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 5442 14464 5448 14476
rect 5403 14436 5448 14464
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 8640 14467 8698 14473
rect 8640 14433 8652 14467
rect 8686 14464 8698 14467
rect 8938 14464 8944 14476
rect 8686 14436 8944 14464
rect 8686 14433 8698 14436
rect 8640 14427 8698 14433
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 10502 14464 10508 14476
rect 10463 14436 10508 14464
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11940 14436 12081 14464
rect 11940 14424 11946 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 15562 14424 15568 14476
rect 15620 14473 15626 14476
rect 15620 14467 15658 14473
rect 15646 14433 15658 14467
rect 15620 14427 15658 14433
rect 15620 14424 15626 14427
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 5166 14396 5172 14408
rect 4387 14368 5172 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 7374 14396 7380 14408
rect 6963 14368 7380 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 1857 14331 1915 14337
rect 1857 14328 1869 14331
rect 1452 14300 1869 14328
rect 1452 14288 1458 14300
rect 1857 14297 1869 14300
rect 1903 14297 1915 14331
rect 1857 14291 1915 14297
rect 1535 14263 1593 14269
rect 1535 14229 1547 14263
rect 1581 14260 1593 14263
rect 1762 14260 1768 14272
rect 1581 14232 1768 14260
rect 1581 14229 1593 14232
rect 1535 14223 1593 14229
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 2832 14232 2881 14260
rect 2832 14220 2838 14232
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 2869 14223 2927 14229
rect 5169 14263 5227 14269
rect 5169 14229 5181 14263
rect 5215 14260 5227 14263
rect 5258 14260 5264 14272
rect 5215 14232 5264 14260
rect 5215 14229 5227 14232
rect 5169 14223 5227 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5629 14263 5687 14269
rect 5629 14260 5641 14263
rect 5592 14232 5641 14260
rect 5592 14220 5598 14232
rect 5629 14229 5641 14232
rect 5675 14229 5687 14263
rect 5629 14223 5687 14229
rect 8711 14263 8769 14269
rect 8711 14229 8723 14263
rect 8757 14260 8769 14263
rect 8846 14260 8852 14272
rect 8757 14232 8852 14260
rect 8757 14229 8769 14232
rect 8711 14223 8769 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 10689 14263 10747 14269
rect 10689 14229 10701 14263
rect 10735 14260 10747 14263
rect 11422 14260 11428 14272
rect 10735 14232 11428 14260
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 12253 14263 12311 14269
rect 12253 14260 12265 14263
rect 12032 14232 12265 14260
rect 12032 14220 12038 14232
rect 12253 14229 12265 14232
rect 12299 14229 12311 14263
rect 12253 14223 12311 14229
rect 15703 14263 15761 14269
rect 15703 14229 15715 14263
rect 15749 14260 15761 14263
rect 15930 14260 15936 14272
rect 15749 14232 15936 14260
rect 15749 14229 15761 14232
rect 15703 14223 15761 14229
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1118 14016 1124 14068
rect 1176 14056 1182 14068
rect 1486 14056 1492 14068
rect 1176 14028 1492 14056
rect 1176 14016 1182 14028
rect 1486 14016 1492 14028
rect 1544 14016 1550 14068
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 3050 14056 3056 14068
rect 2639 14028 3056 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3786 14056 3792 14068
rect 3747 14028 3792 14056
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14056 4307 14059
rect 4522 14056 4528 14068
rect 4295 14028 4528 14056
rect 4295 14025 4307 14028
rect 4249 14019 4307 14025
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 5442 14056 5448 14068
rect 5403 14028 5448 14056
rect 5442 14016 5448 14028
rect 5500 14056 5506 14068
rect 7006 14056 7012 14068
rect 5500 14028 7012 14056
rect 5500 14016 5506 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7466 14056 7472 14068
rect 7116 14028 7472 14056
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 3200 13960 3249 13988
rect 3200 13948 3206 13960
rect 3237 13957 3249 13960
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 1486 13920 1492 13932
rect 1447 13892 1492 13920
rect 1486 13880 1492 13892
rect 1544 13880 1550 13932
rect 3804 13920 3832 14016
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 6273 13991 6331 13997
rect 6273 13988 6285 13991
rect 5316 13960 6285 13988
rect 5316 13948 5322 13960
rect 6273 13957 6285 13960
rect 6319 13988 6331 13991
rect 7116 13988 7144 14028
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 10870 14056 10876 14068
rect 10560 14028 10876 14056
rect 10560 14016 10566 14028
rect 10870 14016 10876 14028
rect 10928 14056 10934 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10928 14028 11069 14056
rect 10928 14016 10934 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 12894 14056 12900 14068
rect 11057 14019 11115 14025
rect 12544 14028 12900 14056
rect 6319 13960 7144 13988
rect 6319 13957 6331 13960
rect 6273 13951 6331 13957
rect 7282 13948 7288 14000
rect 7340 13948 7346 14000
rect 9217 13991 9275 13997
rect 9217 13988 9229 13991
rect 8404 13960 9229 13988
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 3804 13892 4445 13920
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 7300 13920 7328 13948
rect 4433 13883 4491 13889
rect 7116 13892 8248 13920
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 7116 13861 7144 13892
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3053 13855 3111 13861
rect 3053 13852 3065 13855
rect 3007 13824 3065 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3053 13821 3065 13824
rect 3099 13852 3111 13855
rect 6641 13855 6699 13861
rect 3099 13824 4108 13852
rect 3099 13821 3111 13824
rect 3053 13815 3111 13821
rect 4080 13784 4108 13824
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 6687 13824 7113 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13852 7435 13855
rect 7466 13852 7472 13864
rect 7423 13824 7472 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 4154 13784 4160 13796
rect 4080 13756 4160 13784
rect 4154 13744 4160 13756
rect 4212 13744 4218 13796
rect 4522 13744 4528 13796
rect 4580 13784 4586 13796
rect 5077 13787 5135 13793
rect 4580 13756 4625 13784
rect 4580 13744 4586 13756
rect 5077 13753 5089 13787
rect 5123 13784 5135 13787
rect 5442 13784 5448 13796
rect 5123 13756 5448 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 8220 13784 8248 13892
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8404 13861 8432 13960
rect 9217 13957 9229 13960
rect 9263 13957 9275 13991
rect 9217 13951 9275 13957
rect 9723 13991 9781 13997
rect 9723 13957 9735 13991
rect 9769 13988 9781 13991
rect 10686 13988 10692 14000
rect 9769 13960 10692 13988
rect 9769 13957 9781 13960
rect 9723 13951 9781 13957
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 12544 13988 12572 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 10827 13960 12572 13988
rect 12621 13991 12679 13997
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 12621 13957 12633 13991
rect 12667 13988 12679 13991
rect 12710 13988 12716 14000
rect 12667 13960 12716 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 8527 13923 8585 13929
rect 8527 13889 8539 13923
rect 8573 13920 8585 13923
rect 9030 13920 9036 13932
rect 8573 13892 9036 13920
rect 8573 13889 8585 13892
rect 8527 13883 8585 13889
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 10919 13892 11437 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 11425 13889 11437 13892
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 13464 13892 13952 13920
rect 8404 13855 8482 13861
rect 8404 13852 8436 13855
rect 8352 13824 8436 13852
rect 8352 13812 8358 13824
rect 8424 13821 8436 13824
rect 8470 13821 8482 13855
rect 8938 13852 8944 13864
rect 8899 13824 8944 13852
rect 8424 13815 8482 13821
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 9652 13855 9710 13861
rect 9652 13821 9664 13855
rect 9698 13852 9710 13855
rect 9858 13852 9864 13864
rect 9698 13824 9864 13852
rect 9698 13821 9710 13824
rect 9652 13815 9710 13821
rect 9858 13812 9864 13824
rect 9916 13852 9922 13864
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 9916 13824 10057 13852
rect 9916 13812 9922 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 8754 13784 8760 13796
rect 8220 13756 8760 13784
rect 8754 13744 8760 13756
rect 8812 13744 8818 13796
rect 10612 13784 10640 13815
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 11940 13824 12081 13852
rect 11940 13812 11946 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 12069 13815 12127 13821
rect 12434 13812 12440 13824
rect 12492 13852 12498 13864
rect 13464 13861 13492 13892
rect 13924 13864 13952 13892
rect 13630 13861 13636 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12492 13824 12909 13852
rect 12492 13812 12498 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 13464 13855 13542 13861
rect 13464 13824 13496 13855
rect 12897 13815 12955 13821
rect 13484 13821 13496 13824
rect 13530 13821 13542 13855
rect 13484 13815 13542 13821
rect 13587 13855 13636 13861
rect 13587 13821 13599 13855
rect 13633 13821 13636 13855
rect 13587 13815 13636 13821
rect 13630 13812 13636 13815
rect 13688 13812 13694 13864
rect 13906 13852 13912 13864
rect 13867 13824 13912 13852
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 10778 13784 10784 13796
rect 10612 13756 10784 13784
rect 10778 13744 10784 13756
rect 10836 13784 10842 13796
rect 10873 13787 10931 13793
rect 10873 13784 10885 13787
rect 10836 13756 10885 13784
rect 10836 13744 10842 13756
rect 10873 13753 10885 13756
rect 10919 13753 10931 13787
rect 10873 13747 10931 13753
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2130 13716 2136 13728
rect 1820 13688 2136 13716
rect 1820 13676 1826 13688
rect 2130 13676 2136 13688
rect 2188 13676 2194 13728
rect 7098 13716 7104 13728
rect 7059 13688 7104 13716
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 4154 13472 4160 13524
rect 4212 13521 4218 13524
rect 4212 13515 4261 13521
rect 4212 13481 4215 13515
rect 4249 13481 4261 13515
rect 8754 13512 8760 13524
rect 8715 13484 8760 13512
rect 4212 13475 4261 13481
rect 4212 13472 4218 13475
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 10778 13512 10784 13524
rect 10739 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 2130 13444 2136 13456
rect 2091 13416 2136 13444
rect 2130 13404 2136 13416
rect 2188 13404 2194 13456
rect 5534 13444 5540 13456
rect 5495 13416 5540 13444
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 7101 13447 7159 13453
rect 7101 13444 7113 13447
rect 7064 13416 7113 13444
rect 7064 13404 7070 13416
rect 7101 13413 7113 13416
rect 7147 13413 7159 13447
rect 7101 13407 7159 13413
rect 4154 13385 4160 13388
rect 4132 13379 4160 13385
rect 4132 13376 4144 13379
rect 4067 13348 4144 13376
rect 4132 13345 4144 13348
rect 4212 13376 4218 13388
rect 8573 13379 8631 13385
rect 4212 13348 5120 13376
rect 4132 13339 4160 13345
rect 4154 13336 4160 13339
rect 4212 13336 4218 13348
rect 1210 13268 1216 13320
rect 1268 13308 1274 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1268 13280 2053 13308
rect 1268 13268 1274 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 1118 13200 1124 13252
rect 1176 13240 1182 13252
rect 2314 13240 2320 13252
rect 1176 13212 2320 13240
rect 1176 13200 1182 13212
rect 2314 13200 2320 13212
rect 2372 13200 2378 13252
rect 2593 13243 2651 13249
rect 2593 13209 2605 13243
rect 2639 13209 2651 13243
rect 5092 13240 5120 13348
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 8662 13376 8668 13388
rect 8619 13348 8668 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 11790 13376 11796 13388
rect 9732 13348 9777 13376
rect 11751 13348 11796 13376
rect 9732 13336 9738 13348
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13345 13047 13379
rect 13998 13376 14004 13388
rect 13959 13348 14004 13376
rect 12989 13339 13047 13345
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5445 13311 5503 13317
rect 5445 13308 5457 13311
rect 5224 13280 5457 13308
rect 5224 13268 5230 13280
rect 5445 13277 5457 13280
rect 5491 13277 5503 13311
rect 7006 13308 7012 13320
rect 6967 13280 7012 13308
rect 5445 13271 5503 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 5997 13243 6055 13249
rect 5997 13240 6009 13243
rect 5092 13212 6009 13240
rect 2593 13203 2651 13209
rect 5997 13209 6009 13212
rect 6043 13240 6055 13243
rect 7300 13240 7328 13271
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 13004 13308 13032 13339
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 15378 13336 15384 13388
rect 15436 13385 15442 13388
rect 15436 13379 15474 13385
rect 15462 13345 15474 13379
rect 15436 13339 15474 13345
rect 15436 13336 15442 13339
rect 13446 13308 13452 13320
rect 11204 13280 13452 13308
rect 11204 13268 11210 13280
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 6043 13212 7328 13240
rect 6043 13209 6055 13212
rect 5997 13203 6055 13209
rect 2608 13172 2636 13203
rect 3050 13172 3056 13184
rect 2608 13144 3056 13172
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 4890 13172 4896 13184
rect 4851 13144 4896 13172
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 9861 13175 9919 13181
rect 9861 13172 9873 13175
rect 9824 13144 9873 13172
rect 9824 13132 9830 13144
rect 9861 13141 9873 13144
rect 9907 13141 9919 13175
rect 10410 13172 10416 13184
rect 10371 13144 10416 13172
rect 9861 13135 9919 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 11698 13172 11704 13184
rect 11659 13144 11704 13172
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 13354 13172 13360 13184
rect 13219 13144 13360 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 14185 13175 14243 13181
rect 14185 13141 14197 13175
rect 14231 13172 14243 13175
rect 14642 13172 14648 13184
rect 14231 13144 14648 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 15519 13175 15577 13181
rect 15519 13141 15531 13175
rect 15565 13172 15577 13175
rect 16390 13172 16396 13184
rect 15565 13144 16396 13172
rect 15565 13141 15577 13144
rect 15519 13135 15577 13141
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 1762 12968 1768 12980
rect 1719 12940 1768 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 2041 12971 2099 12977
rect 2041 12937 2053 12971
rect 2087 12968 2099 12971
rect 2130 12968 2136 12980
rect 2087 12940 2136 12968
rect 2087 12937 2099 12940
rect 2041 12931 2099 12937
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 2424 12940 3341 12968
rect 1210 12860 1216 12912
rect 1268 12900 1274 12912
rect 2424 12900 2452 12940
rect 3329 12937 3341 12940
rect 3375 12937 3387 12971
rect 4154 12968 4160 12980
rect 4115 12940 4160 12968
rect 3329 12931 3387 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5592 12940 5825 12968
rect 5592 12928 5598 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7101 12971 7159 12977
rect 7101 12968 7113 12971
rect 6972 12940 7113 12968
rect 6972 12928 6978 12940
rect 7101 12937 7113 12940
rect 7147 12968 7159 12971
rect 7190 12968 7196 12980
rect 7147 12940 7196 12968
rect 7147 12937 7159 12940
rect 7101 12931 7159 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 10486 12971 10544 12977
rect 10486 12937 10498 12971
rect 10532 12968 10544 12971
rect 11514 12968 11520 12980
rect 10532 12940 11520 12968
rect 10532 12937 10544 12940
rect 10486 12931 10544 12937
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13446 12968 13452 12980
rect 13407 12940 13452 12968
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 14461 12971 14519 12977
rect 14461 12968 14473 12971
rect 14056 12940 14473 12968
rect 14056 12928 14062 12940
rect 14461 12937 14473 12940
rect 14507 12937 14519 12971
rect 14461 12931 14519 12937
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15436 12940 15853 12968
rect 15436 12928 15442 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 15841 12931 15899 12937
rect 1268 12872 2452 12900
rect 1268 12860 1274 12872
rect 2682 12860 2688 12912
rect 2740 12900 2746 12912
rect 2961 12903 3019 12909
rect 2961 12900 2973 12903
rect 2740 12872 2973 12900
rect 2740 12860 2746 12872
rect 2961 12869 2973 12872
rect 3007 12869 3019 12903
rect 5442 12900 5448 12912
rect 5403 12872 5448 12900
rect 2961 12863 3019 12869
rect 5442 12860 5448 12872
rect 5500 12900 5506 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 5500 12872 6561 12900
rect 5500 12860 5506 12872
rect 6549 12869 6561 12872
rect 6595 12900 6607 12903
rect 7006 12900 7012 12912
rect 6595 12872 7012 12900
rect 6595 12869 6607 12872
rect 6549 12863 6607 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 8662 12900 8668 12912
rect 8623 12872 8668 12900
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 10597 12903 10655 12909
rect 10597 12869 10609 12903
rect 10643 12900 10655 12903
rect 10870 12900 10876 12912
rect 10643 12872 10876 12900
rect 10643 12869 10655 12872
rect 10597 12863 10655 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 3050 12832 3056 12844
rect 2455 12804 3056 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 4890 12832 4896 12844
rect 4851 12804 4896 12832
rect 4890 12792 4896 12804
rect 4948 12832 4954 12844
rect 5350 12832 5356 12844
rect 4948 12804 5356 12832
rect 4948 12792 4954 12804
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 7466 12832 7472 12844
rect 7379 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12832 7530 12844
rect 7742 12832 7748 12844
rect 7524 12804 7748 12832
rect 7524 12792 7530 12804
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 10686 12832 10692 12844
rect 10647 12804 10692 12832
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 14608 12804 15091 12832
rect 14608 12792 14614 12804
rect 9125 12767 9183 12773
rect 9125 12733 9137 12767
rect 9171 12764 9183 12767
rect 9674 12764 9680 12776
rect 9171 12736 9680 12764
rect 9171 12733 9183 12736
rect 9125 12727 9183 12733
rect 9674 12724 9680 12736
rect 9732 12764 9738 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9732 12736 10057 12764
rect 9732 12724 9738 12736
rect 10045 12733 10057 12736
rect 10091 12764 10103 12767
rect 10226 12764 10232 12776
rect 10091 12736 10232 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10704 12764 10732 12792
rect 10870 12764 10876 12776
rect 10704 12736 10876 12764
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 12299 12736 12541 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12529 12733 12541 12736
rect 12575 12764 12587 12767
rect 12802 12764 12808 12776
rect 12575 12736 12808 12764
rect 12575 12733 12587 12736
rect 12529 12727 12587 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 14001 12767 14059 12773
rect 14001 12733 14013 12767
rect 14047 12764 14059 12767
rect 14090 12764 14096 12776
rect 14047 12736 14096 12764
rect 14047 12733 14059 12736
rect 14001 12727 14059 12733
rect 14090 12724 14096 12736
rect 14148 12764 14154 12776
rect 15063 12773 15091 12804
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 14148 12736 14841 12764
rect 14148 12724 14154 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 15048 12767 15106 12773
rect 15048 12733 15060 12767
rect 15094 12764 15106 12767
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 15094 12736 15485 12764
rect 15094 12733 15106 12736
rect 15048 12727 15106 12733
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 16022 12724 16028 12776
rect 16080 12773 16086 12776
rect 16080 12767 16118 12773
rect 16106 12764 16118 12767
rect 16485 12767 16543 12773
rect 16485 12764 16497 12767
rect 16106 12736 16497 12764
rect 16106 12733 16118 12736
rect 16080 12727 16118 12733
rect 16485 12733 16497 12736
rect 16531 12733 16543 12767
rect 16485 12727 16543 12733
rect 16080 12724 16086 12727
rect 1118 12656 1124 12708
rect 1176 12696 1182 12708
rect 1670 12696 1676 12708
rect 1176 12668 1676 12696
rect 1176 12656 1182 12668
rect 1670 12656 1676 12668
rect 1728 12656 1734 12708
rect 1762 12656 1768 12708
rect 1820 12696 1826 12708
rect 2501 12699 2559 12705
rect 2501 12696 2513 12699
rect 1820 12668 2513 12696
rect 1820 12656 1826 12668
rect 2501 12665 2513 12668
rect 2547 12665 2559 12699
rect 2501 12659 2559 12665
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 4709 12699 4767 12705
rect 4709 12696 4721 12699
rect 4672 12668 4721 12696
rect 4672 12656 4678 12668
rect 4709 12665 4721 12668
rect 4755 12696 4767 12699
rect 4985 12699 5043 12705
rect 4985 12696 4997 12699
rect 4755 12668 4997 12696
rect 4755 12665 4767 12668
rect 4709 12659 4767 12665
rect 4985 12665 4997 12668
rect 5031 12665 5043 12699
rect 4985 12659 5043 12665
rect 1210 12588 1216 12640
rect 1268 12628 1274 12640
rect 1394 12628 1400 12640
rect 1268 12600 1400 12628
rect 1268 12588 1274 12600
rect 1394 12588 1400 12600
rect 1452 12588 1458 12640
rect 5000 12628 5028 12659
rect 5166 12656 5172 12708
rect 5224 12696 5230 12708
rect 6181 12699 6239 12705
rect 6181 12696 6193 12699
rect 5224 12668 6193 12696
rect 5224 12656 5230 12668
rect 6181 12665 6193 12668
rect 6227 12665 6239 12699
rect 7650 12696 7656 12708
rect 7611 12668 7656 12696
rect 6181 12659 6239 12665
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 10321 12699 10379 12705
rect 7800 12668 7845 12696
rect 7800 12656 7806 12668
rect 10321 12665 10333 12699
rect 10367 12696 10379 12699
rect 10410 12696 10416 12708
rect 10367 12668 10416 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 10410 12656 10416 12668
rect 10468 12696 10474 12708
rect 11146 12696 11152 12708
rect 10468 12668 11152 12696
rect 10468 12656 10474 12668
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 13170 12696 13176 12708
rect 13131 12668 13176 12696
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 15151 12699 15209 12705
rect 15151 12696 15163 12699
rect 13596 12668 15163 12696
rect 13596 12656 13602 12668
rect 15151 12665 15163 12668
rect 15197 12665 15209 12699
rect 15151 12659 15209 12665
rect 5902 12628 5908 12640
rect 5000 12600 5908 12628
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 9306 12628 9312 12640
rect 9267 12600 9312 12628
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10100 12600 10977 12628
rect 10100 12588 10106 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11425 12631 11483 12637
rect 11425 12597 11437 12631
rect 11471 12628 11483 12631
rect 11514 12628 11520 12640
rect 11471 12600 11520 12628
rect 11471 12597 11483 12600
rect 11425 12591 11483 12597
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 16206 12637 16212 12640
rect 16163 12631 16212 12637
rect 16163 12597 16175 12631
rect 16209 12597 16212 12631
rect 16163 12591 16212 12597
rect 16206 12588 16212 12591
rect 16264 12588 16270 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 5902 12424 5908 12436
rect 5863 12396 5908 12424
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7248 12396 7665 12424
rect 7248 12384 7254 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 9674 12424 9680 12436
rect 8720 12396 9680 12424
rect 8720 12384 8726 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 9824 12396 11100 12424
rect 9824 12384 9830 12396
rect 11072 12368 11100 12396
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12584 12396 12633 12424
rect 12584 12384 12590 12396
rect 12621 12393 12633 12396
rect 12667 12424 12679 12427
rect 14182 12424 14188 12436
rect 12667 12396 14188 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 2133 12359 2191 12365
rect 2133 12356 2145 12359
rect 2096 12328 2145 12356
rect 2096 12316 2102 12328
rect 2133 12325 2145 12328
rect 2179 12325 2191 12359
rect 2682 12356 2688 12368
rect 2643 12328 2688 12356
rect 2133 12319 2191 12325
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 4893 12359 4951 12365
rect 4893 12325 4905 12359
rect 4939 12356 4951 12359
rect 5166 12356 5172 12368
rect 4939 12328 5172 12356
rect 4939 12325 4951 12328
rect 4893 12319 4951 12325
rect 5166 12316 5172 12328
rect 5224 12356 5230 12368
rect 5347 12359 5405 12365
rect 5347 12356 5359 12359
rect 5224 12328 5359 12356
rect 5224 12316 5230 12328
rect 5347 12325 5359 12328
rect 5393 12356 5405 12359
rect 7006 12356 7012 12368
rect 5393 12328 7012 12356
rect 5393 12325 5405 12328
rect 5347 12319 5405 12325
rect 7006 12316 7012 12328
rect 7064 12365 7070 12368
rect 7064 12359 7112 12365
rect 7064 12325 7066 12359
rect 7100 12325 7112 12359
rect 7064 12319 7112 12325
rect 7064 12316 7070 12319
rect 11054 12316 11060 12368
rect 11112 12316 11118 12368
rect 11606 12356 11612 12368
rect 11567 12328 11612 12356
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 13170 12356 13176 12368
rect 13131 12328 13176 12356
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 9766 12288 9772 12300
rect 9727 12260 9772 12288
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 15378 12288 15384 12300
rect 15339 12260 15384 12288
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2130 12220 2136 12232
rect 2087 12192 2136 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 6086 12220 6092 12232
rect 5031 12192 6092 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 7098 12220 7104 12232
rect 6779 12192 7104 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 7098 12180 7104 12192
rect 7156 12220 7162 12232
rect 7466 12220 7472 12232
rect 7156 12192 7472 12220
rect 7156 12180 7162 12192
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9640 12192 9689 12220
rect 9640 12180 9646 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 11330 12220 11336 12232
rect 10928 12192 11336 12220
rect 10928 12180 10934 12192
rect 11330 12180 11336 12192
rect 11388 12220 11394 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11388 12192 11529 12220
rect 11388 12180 11394 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 12158 12180 12164 12232
rect 12216 12220 12222 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12216 12192 13093 12220
rect 12216 12180 12222 12192
rect 13081 12189 13093 12192
rect 13127 12220 13139 12223
rect 13722 12220 13728 12232
rect 13127 12192 13728 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 12069 12155 12127 12161
rect 12069 12121 12081 12155
rect 12115 12152 12127 12155
rect 12342 12152 12348 12164
rect 12115 12124 12348 12152
rect 12115 12121 12127 12124
rect 12069 12115 12127 12121
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 13633 12155 13691 12161
rect 13633 12121 13645 12155
rect 13679 12152 13691 12155
rect 13998 12152 14004 12164
rect 13679 12124 14004 12152
rect 13679 12121 13691 12124
rect 13633 12115 13691 12121
rect 13998 12112 14004 12124
rect 14056 12112 14062 12164
rect 1670 12084 1676 12096
rect 1631 12056 1676 12084
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 2961 12087 3019 12093
rect 2961 12084 2973 12087
rect 2924 12056 2973 12084
rect 2924 12044 2930 12056
rect 2961 12053 2973 12056
rect 3007 12084 3019 12087
rect 3418 12084 3424 12096
rect 3007 12056 3424 12084
rect 3007 12053 3019 12056
rect 2961 12047 3019 12053
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7892 12056 7941 12084
rect 7892 12044 7898 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 10781 12087 10839 12093
rect 10781 12053 10793 12087
rect 10827 12084 10839 12087
rect 10870 12084 10876 12096
rect 10827 12056 10876 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 15746 12084 15752 12096
rect 15707 12056 15752 12084
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 2188 11852 2329 11880
rect 2188 11840 2194 11852
rect 2317 11849 2329 11852
rect 2363 11849 2375 11883
rect 6086 11880 6092 11892
rect 6047 11852 6092 11880
rect 2317 11843 2375 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 9766 11880 9772 11892
rect 9727 11852 9772 11880
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11606 11880 11612 11892
rect 11563 11852 11612 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 12618 11840 12624 11892
rect 12676 11889 12682 11892
rect 12676 11883 12725 11889
rect 12676 11849 12679 11883
rect 12713 11849 12725 11883
rect 12676 11843 12725 11849
rect 12676 11840 12682 11843
rect 13170 11840 13176 11892
rect 13228 11880 13234 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13228 11852 13553 11880
rect 13228 11840 13234 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13780 11852 13921 11880
rect 13780 11840 13786 11852
rect 13909 11849 13921 11852
rect 13955 11849 13967 11883
rect 13909 11843 13967 11849
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 15378 11880 15384 11892
rect 14507 11852 15384 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 11793 11815 11851 11821
rect 11793 11812 11805 11815
rect 11480 11784 11805 11812
rect 11480 11772 11486 11784
rect 11793 11781 11805 11784
rect 11839 11781 11851 11815
rect 12805 11815 12863 11821
rect 12805 11812 12817 11815
rect 11793 11775 11851 11781
rect 12452 11784 12817 11812
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7006 11744 7012 11756
rect 6687 11716 7012 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7006 11704 7012 11716
rect 7064 11744 7070 11756
rect 7650 11744 7656 11756
rect 7064 11716 7656 11744
rect 7064 11704 7070 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 7926 11744 7932 11756
rect 7883 11716 7932 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 7926 11704 7932 11716
rect 7984 11744 7990 11756
rect 10042 11744 10048 11756
rect 7984 11716 10048 11744
rect 7984 11704 7990 11716
rect 10042 11704 10048 11716
rect 10100 11744 10106 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 10100 11716 10333 11744
rect 10100 11704 10106 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10321 11707 10379 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11808 11744 11836 11775
rect 12452 11744 12480 11784
rect 12805 11781 12817 11784
rect 12851 11812 12863 11815
rect 12851 11784 13032 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 12894 11744 12900 11756
rect 11808 11716 12480 11744
rect 12855 11716 12900 11744
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1670 11676 1676 11688
rect 1443 11648 1676 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 4801 11679 4859 11685
rect 4801 11676 4813 11679
rect 4264 11648 4813 11676
rect 2777 11611 2835 11617
rect 2777 11577 2789 11611
rect 2823 11577 2835 11611
rect 2777 11571 2835 11577
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2792 11540 2820 11571
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 2924 11580 2969 11608
rect 2924 11568 2930 11580
rect 4264 11552 4292 11648
rect 4801 11645 4813 11648
rect 4847 11645 4859 11679
rect 5718 11676 5724 11688
rect 5679 11648 5724 11676
rect 4801 11639 4859 11645
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 8619 11648 9321 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9309 11645 9321 11648
rect 9355 11676 9367 11679
rect 12526 11676 12532 11688
rect 9355 11648 10180 11676
rect 12487 11648 12532 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 5166 11617 5172 11620
rect 4709 11611 4767 11617
rect 4709 11577 4721 11611
rect 4755 11608 4767 11611
rect 5163 11608 5172 11617
rect 4755 11580 5172 11608
rect 4755 11577 4767 11580
rect 4709 11571 4767 11577
rect 5163 11571 5172 11580
rect 5166 11568 5172 11571
rect 5224 11568 5230 11620
rect 7190 11608 7196 11620
rect 7151 11580 7196 11608
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 7282 11568 7288 11620
rect 7340 11608 7346 11620
rect 9398 11608 9404 11620
rect 7340 11580 7385 11608
rect 9359 11580 9404 11608
rect 7340 11568 7346 11580
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 3694 11540 3700 11552
rect 2792 11512 3700 11540
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 4246 11540 4252 11552
rect 4207 11512 4252 11540
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 7208 11540 7236 11568
rect 10152 11549 10180 11648
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 10413 11611 10471 11617
rect 10413 11577 10425 11611
rect 10459 11608 10471 11611
rect 10686 11608 10692 11620
rect 10459 11580 10692 11608
rect 10459 11577 10471 11580
rect 10413 11571 10471 11577
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 7208 11512 8125 11540
rect 8113 11509 8125 11512
rect 8159 11509 8171 11543
rect 8113 11503 8171 11509
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10428 11540 10456 11571
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 12894 11568 12900 11620
rect 12952 11608 12958 11620
rect 13004 11608 13032 11784
rect 12952 11580 13032 11608
rect 13265 11611 13323 11617
rect 12952 11568 12958 11580
rect 13265 11577 13277 11611
rect 13311 11608 13323 11611
rect 13354 11608 13360 11620
rect 13311 11580 13360 11608
rect 13311 11577 13323 11580
rect 13265 11571 13323 11577
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 14553 11611 14611 11617
rect 14553 11577 14565 11611
rect 14599 11608 14611 11611
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 14599 11580 15117 11608
rect 14599 11577 14611 11580
rect 14553 11571 14611 11577
rect 15105 11577 15117 11580
rect 15151 11608 15163 11611
rect 15657 11611 15715 11617
rect 15657 11608 15669 11611
rect 15151 11580 15669 11608
rect 15151 11577 15163 11580
rect 15105 11571 15163 11577
rect 15657 11577 15669 11580
rect 15703 11577 15715 11611
rect 15657 11571 15715 11577
rect 15749 11611 15807 11617
rect 15749 11577 15761 11611
rect 15795 11608 15807 11611
rect 16114 11608 16120 11620
rect 15795 11580 16120 11608
rect 15795 11577 15807 11580
rect 15749 11571 15807 11577
rect 10183 11512 10456 11540
rect 12253 11543 12311 11549
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12618 11540 12624 11552
rect 12299 11512 12624 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 15473 11543 15531 11549
rect 15473 11509 15485 11543
rect 15519 11540 15531 11543
rect 15764 11540 15792 11571
rect 16114 11568 16120 11580
rect 16172 11568 16178 11620
rect 16298 11608 16304 11620
rect 16259 11580 16304 11608
rect 16298 11568 16304 11580
rect 16356 11568 16362 11620
rect 15519 11512 15792 11540
rect 15519 11509 15531 11512
rect 15473 11503 15531 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1535 11339 1593 11345
rect 1535 11305 1547 11339
rect 1581 11336 1593 11339
rect 1670 11336 1676 11348
rect 1581 11308 1676 11336
rect 1581 11305 1593 11308
rect 1535 11299 1593 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2556 11308 3433 11336
rect 2556 11296 2562 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5592 11308 5733 11336
rect 5592 11296 5598 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 6362 11336 6368 11348
rect 6323 11308 6368 11336
rect 5721 11299 5779 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 7466 11336 7472 11348
rect 7427 11308 7472 11336
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 10100 11308 10701 11336
rect 10100 11296 10106 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 10689 11299 10747 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 12802 11336 12808 11348
rect 12763 11308 12808 11336
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 13044 11308 13093 11336
rect 13044 11296 13050 11308
rect 13081 11305 13093 11308
rect 13127 11336 13139 11339
rect 13446 11336 13452 11348
rect 13127 11308 13452 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13630 11336 13636 11348
rect 13587 11308 13636 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13630 11296 13636 11308
rect 13688 11336 13694 11348
rect 13688 11308 13768 11336
rect 13688 11296 13694 11308
rect 3145 11271 3203 11277
rect 3145 11237 3157 11271
rect 3191 11268 3203 11271
rect 4246 11268 4252 11280
rect 3191 11240 4252 11268
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 5166 11277 5172 11280
rect 5163 11268 5172 11277
rect 5127 11240 5172 11268
rect 5163 11231 5172 11240
rect 5166 11228 5172 11231
rect 5224 11228 5230 11280
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 1670 11200 1676 11212
rect 1510 11172 1676 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 1670 11160 1676 11172
rect 1728 11200 1734 11212
rect 1949 11203 2007 11209
rect 1728 11172 1900 11200
rect 1728 11160 1734 11172
rect 1872 11132 1900 11172
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 2038 11200 2044 11212
rect 1995 11172 2044 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2866 11200 2872 11212
rect 2731 11172 2872 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 3510 11200 3516 11212
rect 3007 11172 3516 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 6380 11200 6408 11296
rect 7558 11228 7564 11280
rect 7616 11268 7622 11280
rect 7616 11240 7788 11268
rect 7616 11228 7622 11240
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 6380 11172 6561 11200
rect 6549 11169 6561 11172
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11200 7251 11203
rect 7282 11200 7288 11212
rect 7239 11172 7288 11200
rect 7239 11169 7251 11172
rect 7193 11163 7251 11169
rect 7282 11160 7288 11172
rect 7340 11200 7346 11212
rect 7760 11209 7788 11240
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9456 11240 9873 11268
rect 9456 11228 9462 11240
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 9861 11231 9919 11237
rect 10410 11228 10416 11240
rect 10468 11268 10474 11280
rect 10778 11268 10784 11280
rect 10468 11240 10784 11268
rect 10468 11228 10474 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 10928 11240 11008 11268
rect 10928 11228 10934 11240
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7340 11172 7665 11200
rect 7340 11160 7346 11172
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 3326 11132 3332 11144
rect 1872 11104 3332 11132
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 4212 11104 4813 11132
rect 4212 11092 4218 11104
rect 4801 11101 4813 11104
rect 4847 11132 4859 11135
rect 5442 11132 5448 11144
rect 4847 11104 5448 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 8536 11104 9781 11132
rect 8536 11092 8542 11104
rect 9769 11101 9781 11104
rect 9815 11132 9827 11135
rect 10870 11132 10876 11144
rect 9815 11104 10876 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2225 11067 2283 11073
rect 2225 11064 2237 11067
rect 2188 11036 2237 11064
rect 2188 11024 2194 11036
rect 2225 11033 2237 11036
rect 2271 11033 2283 11067
rect 6730 11064 6736 11076
rect 6691 11036 6736 11064
rect 2225 11027 2283 11033
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 10980 11064 11008 11240
rect 12158 11228 12164 11280
rect 12216 11277 12222 11280
rect 13740 11277 13768 11308
rect 15488 11308 16988 11336
rect 12216 11271 12264 11277
rect 12216 11237 12218 11271
rect 12252 11237 12264 11271
rect 12216 11231 12264 11237
rect 13725 11271 13783 11277
rect 13725 11237 13737 11271
rect 13771 11237 13783 11271
rect 13725 11231 13783 11237
rect 12216 11228 12222 11231
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 13872 11240 13917 11268
rect 13872 11228 13878 11240
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 15488 11277 15516 11308
rect 15473 11271 15531 11277
rect 15473 11268 15485 11271
rect 14884 11240 15485 11268
rect 14884 11228 14890 11240
rect 15473 11237 15485 11240
rect 15519 11237 15531 11271
rect 15473 11231 15531 11237
rect 16025 11271 16083 11277
rect 16025 11237 16037 11271
rect 16071 11268 16083 11271
rect 16298 11268 16304 11280
rect 16071 11240 16304 11268
rect 16071 11237 16083 11240
rect 16025 11231 16083 11237
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 16960 11212 16988 11308
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 16172 11172 16865 11200
rect 16172 11160 16178 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 16853 11163 16911 11169
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 18506 11209 18512 11212
rect 18484 11203 18512 11209
rect 17000 11172 17045 11200
rect 17000 11160 17006 11172
rect 18484 11169 18496 11203
rect 18484 11163 18512 11169
rect 18506 11160 18512 11163
rect 18564 11160 18570 11212
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11101 11943 11135
rect 13998 11132 14004 11144
rect 13959 11104 14004 11132
rect 11885 11095 11943 11101
rect 11698 11064 11704 11076
rect 10100 11036 11008 11064
rect 11659 11036 11704 11064
rect 10100 11024 10106 11036
rect 11698 11024 11704 11036
rect 11756 11064 11762 11076
rect 11900 11064 11928 11095
rect 13998 11092 14004 11104
rect 14056 11132 14062 11144
rect 14734 11132 14740 11144
rect 14056 11104 14740 11132
rect 14056 11092 14062 11104
rect 14734 11092 14740 11104
rect 14792 11132 14798 11144
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 14792 11104 15393 11132
rect 14792 11092 14798 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 11756 11036 11928 11064
rect 11756 11024 11762 11036
rect 12986 11024 12992 11076
rect 13044 11064 13050 11076
rect 14550 11064 14556 11076
rect 13044 11036 14556 11064
rect 13044 11024 13050 11036
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 18555 11067 18613 11073
rect 18555 11033 18567 11067
rect 18601 11064 18613 11067
rect 20162 11064 20168 11076
rect 18601 11036 20168 11064
rect 18601 11033 18613 11036
rect 18555 11027 18613 11033
rect 20162 11024 20168 11036
rect 20220 11024 20226 11076
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11146 10996 11152 11008
rect 10836 10968 11152 10996
rect 10836 10956 10842 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 3694 10752 3700 10804
rect 3752 10792 3758 10804
rect 4062 10792 4068 10804
rect 3752 10764 4068 10792
rect 3752 10752 3758 10764
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4801 10795 4859 10801
rect 4801 10761 4813 10795
rect 4847 10792 4859 10795
rect 5166 10792 5172 10804
rect 4847 10764 5172 10792
rect 4847 10761 4859 10764
rect 4801 10755 4859 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6273 10795 6331 10801
rect 6273 10792 6285 10795
rect 5500 10764 6285 10792
rect 5500 10752 5506 10764
rect 6273 10761 6285 10764
rect 6319 10761 6331 10795
rect 6273 10755 6331 10761
rect 7469 10795 7527 10801
rect 7469 10761 7481 10795
rect 7515 10792 7527 10795
rect 7558 10792 7564 10804
rect 7515 10764 7564 10792
rect 7515 10761 7527 10764
rect 7469 10755 7527 10761
rect 7558 10752 7564 10764
rect 7616 10792 7622 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 7616 10764 8861 10792
rect 7616 10752 7622 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 9398 10792 9404 10804
rect 9263 10764 9404 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 10686 10792 10692 10804
rect 10643 10764 10692 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 10870 10792 10876 10804
rect 10831 10764 10876 10792
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11609 10795 11667 10801
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 11790 10792 11796 10804
rect 11655 10764 11796 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 11790 10752 11796 10764
rect 11848 10792 11854 10804
rect 12434 10792 12440 10804
rect 11848 10764 12440 10792
rect 11848 10752 11854 10764
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13541 10795 13599 10801
rect 13541 10792 13553 10795
rect 12860 10764 13553 10792
rect 12860 10752 12866 10764
rect 13541 10761 13553 10764
rect 13587 10792 13599 10795
rect 13722 10792 13728 10804
rect 13587 10764 13728 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14826 10752 14832 10804
rect 14884 10792 14890 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 14884 10764 15025 10792
rect 14884 10752 14890 10764
rect 15013 10761 15025 10764
rect 15059 10761 15071 10795
rect 15746 10792 15752 10804
rect 15707 10764 15752 10792
rect 15013 10755 15071 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16942 10792 16948 10804
rect 16903 10764 16948 10792
rect 16942 10752 16948 10764
rect 17000 10792 17006 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 17000 10764 17233 10792
rect 17000 10752 17006 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 17221 10755 17279 10761
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 9631 10696 11989 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 1210 10616 1216 10668
rect 1268 10656 1274 10668
rect 1394 10656 1400 10668
rect 1268 10628 1400 10656
rect 1268 10616 1274 10628
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 2498 10656 2504 10668
rect 1903 10628 2504 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 4062 10656 4068 10668
rect 4023 10628 4068 10656
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 1946 10520 1952 10532
rect 1907 10492 1952 10520
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 2498 10520 2504 10532
rect 2459 10492 2504 10520
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3436 10520 3464 10551
rect 3510 10548 3516 10600
rect 3568 10588 3574 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3568 10560 3801 10588
rect 3568 10548 3574 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 5166 10588 5172 10600
rect 4479 10560 5172 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 4062 10520 4068 10532
rect 3283 10492 4068 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 4062 10480 4068 10492
rect 4120 10520 4126 10532
rect 4448 10520 4476 10551
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 7929 10591 7987 10597
rect 5491 10560 6040 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 4120 10492 4476 10520
rect 4120 10480 4126 10492
rect 2866 10452 2872 10464
rect 2779 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10452 2930 10464
rect 3418 10452 3424 10464
rect 2924 10424 3424 10452
rect 2924 10412 2930 10424
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 6012 10461 6040 10560
rect 7929 10557 7941 10591
rect 7975 10588 7987 10591
rect 8754 10588 8760 10600
rect 7975 10560 8760 10588
rect 7975 10557 7987 10560
rect 7929 10551 7987 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9272 10560 9689 10588
rect 9272 10548 9278 10560
rect 9677 10557 9689 10560
rect 9723 10557 9735 10591
rect 9677 10551 9735 10557
rect 7650 10480 7656 10532
rect 7708 10520 7714 10532
rect 10060 10529 10088 10696
rect 11977 10693 11989 10696
rect 12023 10724 12035 10727
rect 12158 10724 12164 10736
rect 12023 10696 12164 10724
rect 12023 10693 12035 10696
rect 11977 10687 12035 10693
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 12342 10684 12348 10736
rect 12400 10724 12406 10736
rect 13170 10724 13176 10736
rect 12400 10696 13176 10724
rect 12400 10684 12406 10696
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 16482 10724 16488 10736
rect 16443 10696 16488 10724
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 13538 10656 13544 10668
rect 12575 10628 13544 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 13872 10560 14105 10588
rect 13872 10548 13878 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 16908 10560 17877 10588
rect 16908 10548 16914 10560
rect 17865 10557 17877 10560
rect 17911 10588 17923 10591
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 17911 10560 18153 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 7837 10523 7895 10529
rect 7837 10520 7849 10523
rect 7708 10492 7849 10520
rect 7708 10480 7714 10492
rect 7837 10489 7849 10492
rect 7883 10520 7895 10523
rect 8291 10523 8349 10529
rect 8291 10520 8303 10523
rect 7883 10492 8303 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8291 10489 8303 10492
rect 8337 10520 8349 10523
rect 10039 10523 10097 10529
rect 10039 10520 10051 10523
rect 8337 10492 10051 10520
rect 8337 10489 8349 10492
rect 8291 10483 8349 10489
rect 10039 10489 10051 10492
rect 10085 10489 10097 10523
rect 10039 10483 10097 10489
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10489 12679 10523
rect 13170 10520 13176 10532
rect 13131 10492 13176 10520
rect 12621 10483 12679 10489
rect 4985 10455 5043 10461
rect 4985 10452 4997 10455
rect 4856 10424 4997 10452
rect 4856 10412 4862 10424
rect 4985 10421 4997 10424
rect 5031 10421 5043 10455
rect 4985 10415 5043 10421
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6454 10452 6460 10464
rect 6043 10424 6460 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12636 10452 12664 10483
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 14414 10523 14472 10529
rect 14414 10520 14426 10523
rect 14016 10492 14426 10520
rect 14016 10464 14044 10492
rect 14414 10489 14426 10492
rect 14460 10489 14472 10523
rect 15933 10523 15991 10529
rect 15933 10520 15945 10523
rect 14414 10483 14472 10489
rect 15304 10492 15945 10520
rect 15304 10464 15332 10492
rect 15933 10489 15945 10492
rect 15979 10489 15991 10523
rect 15933 10483 15991 10489
rect 16025 10523 16083 10529
rect 16025 10489 16037 10523
rect 16071 10489 16083 10523
rect 16025 10483 16083 10489
rect 13998 10452 14004 10464
rect 12492 10424 12664 10452
rect 13959 10424 14004 10452
rect 12492 10412 12498 10424
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 15286 10452 15292 10464
rect 15247 10424 15292 10452
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 16040 10452 16068 10483
rect 17678 10480 17684 10532
rect 17736 10520 17742 10532
rect 18506 10520 18512 10532
rect 17736 10492 18512 10520
rect 17736 10480 17742 10492
rect 18506 10480 18512 10492
rect 18564 10520 18570 10532
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 18564 10492 19073 10520
rect 18564 10480 18570 10492
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19061 10483 19119 10489
rect 18322 10452 18328 10464
rect 15804 10424 16068 10452
rect 18283 10424 18328 10452
rect 15804 10412 15810 10424
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2038 10208 2044 10260
rect 2096 10208 2102 10260
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 3510 10248 3516 10260
rect 2363 10220 3516 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 4798 10248 4804 10260
rect 4759 10220 4804 10248
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 4948 10220 4997 10248
rect 4948 10208 4954 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 4985 10211 5043 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6595 10251 6653 10257
rect 6595 10248 6607 10251
rect 5592 10220 6607 10248
rect 5592 10208 5598 10220
rect 6595 10217 6607 10220
rect 6641 10217 6653 10251
rect 8754 10248 8760 10260
rect 8715 10220 8760 10248
rect 6595 10211 6653 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 12434 10248 12440 10260
rect 12391 10220 12440 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13173 10251 13231 10257
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 13538 10248 13544 10260
rect 13219 10220 13544 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 14369 10251 14427 10257
rect 14369 10217 14381 10251
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 2056 10112 2084 10208
rect 2593 10183 2651 10189
rect 2593 10149 2605 10183
rect 2639 10180 2651 10183
rect 2682 10180 2688 10192
rect 2639 10152 2688 10180
rect 2639 10149 2651 10152
rect 2593 10143 2651 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 7561 10183 7619 10189
rect 7561 10180 7573 10183
rect 7156 10152 7573 10180
rect 7156 10140 7162 10152
rect 7561 10149 7573 10152
rect 7607 10180 7619 10183
rect 10597 10183 10655 10189
rect 7607 10152 8524 10180
rect 7607 10149 7619 10152
rect 7561 10143 7619 10149
rect 1510 10084 2084 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 5074 10112 5080 10124
rect 3476 10084 5080 10112
rect 3476 10072 3482 10084
rect 5074 10072 5080 10084
rect 5132 10112 5138 10124
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 5132 10084 5181 10112
rect 5132 10072 5138 10084
rect 5169 10081 5181 10084
rect 5215 10112 5227 10115
rect 5258 10112 5264 10124
rect 5215 10084 5264 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10013 2559 10047
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 2501 10007 2559 10013
rect 2516 9976 2544 10007
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3510 10044 3516 10056
rect 3471 10016 3516 10044
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 5368 10044 5396 10075
rect 6178 10072 6184 10124
rect 6236 10112 6242 10124
rect 6492 10115 6550 10121
rect 6492 10112 6504 10115
rect 6236 10084 6504 10112
rect 6236 10072 6242 10084
rect 6492 10081 6504 10084
rect 6538 10081 6550 10115
rect 7926 10112 7932 10124
rect 7887 10084 7932 10112
rect 6492 10075 6550 10081
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8496 10121 8524 10152
rect 10597 10149 10609 10183
rect 10643 10180 10655 10183
rect 10686 10180 10692 10192
rect 10643 10152 10692 10180
rect 10643 10149 10655 10152
rect 10597 10143 10655 10149
rect 10686 10140 10692 10152
rect 10744 10180 10750 10192
rect 10962 10180 10968 10192
rect 10744 10152 10968 10180
rect 10744 10140 10750 10152
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 11787 10183 11845 10189
rect 11787 10149 11799 10183
rect 11833 10180 11845 10183
rect 12158 10180 12164 10192
rect 11833 10152 12164 10180
rect 11833 10149 11845 10152
rect 11787 10143 11845 10149
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 13811 10183 13869 10189
rect 13811 10149 13823 10183
rect 13857 10180 13869 10183
rect 13998 10180 14004 10192
rect 13857 10152 14004 10180
rect 13857 10149 13869 10152
rect 13811 10143 13869 10149
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 14384 10180 14412 10211
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14792 10220 15025 10248
rect 14792 10208 14798 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 16390 10248 16396 10260
rect 16351 10220 16396 10248
rect 15013 10211 15071 10217
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 15378 10180 15384 10192
rect 14384 10152 15384 10180
rect 15378 10140 15384 10152
rect 15436 10180 15442 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15436 10152 15485 10180
rect 15436 10140 15442 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 15473 10143 15531 10149
rect 16025 10183 16083 10189
rect 16025 10149 16037 10183
rect 16071 10180 16083 10183
rect 16482 10180 16488 10192
rect 16071 10152 16488 10180
rect 16071 10149 16083 10152
rect 16025 10143 16083 10149
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 17494 10180 17500 10192
rect 17144 10152 17500 10180
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8754 10112 8760 10124
rect 8527 10084 8760 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 4212 10016 5396 10044
rect 7193 10047 7251 10053
rect 4212 10004 4218 10016
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 8128 10044 8156 10075
rect 8754 10072 8760 10084
rect 8812 10112 8818 10124
rect 9306 10112 9312 10124
rect 8812 10084 9312 10112
rect 8812 10072 8818 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10870 10112 10876 10124
rect 10551 10084 10876 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 17144 10121 17172 10152
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 17770 10112 17776 10124
rect 17359 10084 17776 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 19058 10112 19064 10124
rect 19019 10084 19064 10112
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 23474 10072 23480 10124
rect 23532 10112 23538 10124
rect 23604 10115 23662 10121
rect 23604 10112 23616 10115
rect 23532 10084 23616 10112
rect 23532 10072 23538 10084
rect 23604 10081 23616 10084
rect 23650 10081 23662 10115
rect 23604 10075 23662 10081
rect 8570 10044 8576 10056
rect 7239 10016 8576 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 13446 10044 13452 10056
rect 13407 10016 13452 10044
rect 11425 10007 11483 10013
rect 2774 9976 2780 9988
rect 2516 9948 2780 9976
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 11440 9920 11468 10007
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 15746 10044 15752 10056
rect 15427 10016 15752 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 16540 10016 17417 10044
rect 16540 10004 16546 10016
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17405 10007 17463 10013
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 18417 10047 18475 10053
rect 18417 10044 18429 10047
rect 18012 10016 18429 10044
rect 18012 10004 18018 10016
rect 18417 10013 18429 10016
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 14645 9979 14703 9985
rect 14645 9976 14657 9979
rect 13872 9948 14657 9976
rect 13872 9936 13878 9948
rect 14645 9945 14657 9948
rect 14691 9945 14703 9979
rect 14645 9939 14703 9945
rect 1535 9911 1593 9917
rect 1535 9877 1547 9911
rect 1581 9908 1593 9911
rect 1762 9908 1768 9920
rect 1581 9880 1768 9908
rect 1581 9877 1593 9880
rect 1535 9871 1593 9877
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 3234 9908 3240 9920
rect 2924 9880 3240 9908
rect 2924 9868 2930 9880
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 9272 9880 9413 9908
rect 9272 9868 9278 9880
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 11333 9911 11391 9917
rect 11333 9877 11345 9911
rect 11379 9908 11391 9911
rect 11422 9908 11428 9920
rect 11379 9880 11428 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 23707 9911 23765 9917
rect 23707 9877 23719 9911
rect 23753 9908 23765 9911
rect 24118 9908 24124 9920
rect 23753 9880 24124 9908
rect 23753 9877 23765 9880
rect 23707 9871 23765 9877
rect 24118 9868 24124 9880
rect 24176 9868 24182 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2314 9704 2320 9716
rect 1596 9676 2320 9704
rect 1596 9648 1624 9676
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2682 9704 2688 9716
rect 2643 9676 2688 9704
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 6454 9704 6460 9716
rect 2924 9676 3004 9704
rect 2924 9664 2930 9676
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 2038 9636 2044 9648
rect 1688 9608 2044 9636
rect 1210 9528 1216 9580
rect 1268 9568 1274 9580
rect 1688 9568 1716 9608
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 2976 9636 3004 9676
rect 4080 9676 6460 9704
rect 3234 9636 3240 9648
rect 2976 9608 3240 9636
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 1268 9540 1716 9568
rect 1268 9528 1274 9540
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3418 9500 3424 9512
rect 3099 9472 3424 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3697 9503 3755 9509
rect 3697 9500 3709 9503
rect 3568 9472 3709 9500
rect 3568 9460 3574 9472
rect 3697 9469 3709 9472
rect 3743 9500 3755 9503
rect 4080 9500 4108 9676
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 7098 9704 7104 9716
rect 6840 9676 7104 9704
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 5592 9608 6009 9636
rect 5592 9596 5598 9608
rect 5997 9605 6009 9608
rect 6043 9636 6055 9639
rect 6840 9636 6868 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 9953 9707 10011 9713
rect 9272 9676 9317 9704
rect 9272 9664 9278 9676
rect 9953 9673 9965 9707
rect 9999 9704 10011 9707
rect 10870 9704 10876 9716
rect 9999 9676 10876 9704
rect 9999 9673 10011 9676
rect 9953 9667 10011 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 12158 9704 12164 9716
rect 11931 9676 12164 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 12158 9664 12164 9676
rect 12216 9704 12222 9716
rect 13817 9707 13875 9713
rect 13817 9704 13829 9707
rect 12216 9676 13829 9704
rect 12216 9664 12222 9676
rect 13817 9673 13829 9676
rect 13863 9704 13875 9707
rect 13998 9704 14004 9716
rect 13863 9676 14004 9704
rect 13863 9673 13875 9676
rect 13817 9667 13875 9673
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15436 9676 15853 9704
rect 15436 9664 15442 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 17494 9704 17500 9716
rect 15841 9667 15899 9673
rect 15948 9676 17500 9704
rect 6043 9608 6868 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 6914 9596 6920 9648
rect 6972 9645 6978 9648
rect 6972 9639 7021 9645
rect 6972 9605 6975 9639
rect 7009 9605 7021 9639
rect 6972 9599 7021 9605
rect 6972 9596 6978 9599
rect 7374 9596 7380 9648
rect 7432 9596 7438 9648
rect 10689 9639 10747 9645
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 10962 9636 10968 9648
rect 10735 9608 10968 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4798 9568 4804 9580
rect 4755 9540 4804 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7392 9568 7420 9596
rect 7331 9540 8708 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 8680 9512 8708 9540
rect 3743 9472 4108 9500
rect 6892 9503 6950 9509
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 6892 9469 6904 9503
rect 6938 9500 6950 9503
rect 7374 9500 7380 9512
rect 6938 9472 7380 9500
rect 6938 9469 6950 9472
rect 6892 9463 6950 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 7926 9500 7932 9512
rect 7791 9472 7932 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 7926 9460 7932 9472
rect 7984 9500 7990 9512
rect 8386 9500 8392 9512
rect 7984 9472 8392 9500
rect 7984 9460 7990 9472
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 10796 9509 10824 9608
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 14737 9639 14795 9645
rect 14737 9605 14749 9639
rect 14783 9636 14795 9639
rect 15948 9636 15976 9676
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 17770 9704 17776 9716
rect 17731 9676 17776 9704
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 19058 9704 19064 9716
rect 19019 9676 19064 9704
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 23474 9704 23480 9716
rect 23435 9676 23480 9704
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 14783 9608 15976 9636
rect 14783 9605 14795 9608
rect 14737 9599 14795 9605
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11698 9568 11704 9580
rect 11563 9540 11704 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13814 9568 13820 9580
rect 13495 9540 13820 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8720 9472 8953 9500
rect 8720 9460 8726 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9469 11299 9503
rect 11241 9463 11299 9469
rect 1673 9435 1731 9441
rect 1673 9401 1685 9435
rect 1719 9401 1731 9435
rect 1673 9395 1731 9401
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 2038 9432 2044 9444
rect 1811 9404 2044 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 1688 9364 1716 9395
rect 2038 9392 2044 9404
rect 2096 9392 2102 9444
rect 2130 9392 2136 9444
rect 2188 9392 2194 9444
rect 2317 9435 2375 9441
rect 2317 9401 2329 9435
rect 2363 9432 2375 9435
rect 2498 9432 2504 9444
rect 2363 9404 2504 9432
rect 2363 9401 2375 9404
rect 2317 9395 2375 9401
rect 2498 9392 2504 9404
rect 2556 9432 2562 9444
rect 2682 9432 2688 9444
rect 2556 9404 2688 9432
rect 2556 9392 2562 9404
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 3878 9432 3884 9444
rect 3839 9404 3884 9432
rect 3878 9392 3884 9404
rect 3936 9392 3942 9444
rect 5074 9441 5080 9444
rect 4617 9435 4675 9441
rect 4617 9401 4629 9435
rect 4663 9432 4675 9435
rect 5071 9432 5080 9441
rect 4663 9404 5080 9432
rect 4663 9401 4675 9404
rect 4617 9395 4675 9401
rect 5071 9395 5080 9404
rect 5074 9392 5080 9395
rect 5132 9392 5138 9444
rect 8588 9432 8616 9460
rect 9306 9432 9312 9444
rect 8588 9404 9312 9432
rect 9306 9392 9312 9404
rect 9364 9432 9370 9444
rect 9493 9435 9551 9441
rect 9493 9432 9505 9435
rect 9364 9404 9505 9432
rect 9364 9392 9370 9404
rect 9493 9401 9505 9404
rect 9539 9401 9551 9435
rect 9493 9395 9551 9401
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9432 10379 9435
rect 11256 9432 11284 9463
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12768 9472 13001 9500
rect 12768 9460 12774 9472
rect 12989 9469 13001 9472
rect 13035 9500 13047 9503
rect 13078 9500 13084 9512
rect 13035 9472 13084 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14844 9509 14872 9608
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 16448 9608 16528 9636
rect 16448 9596 16454 9608
rect 16500 9577 16528 9608
rect 20162 9596 20168 9648
rect 20220 9636 20226 9648
rect 20438 9636 20444 9648
rect 20220 9608 20444 9636
rect 20220 9596 20226 9608
rect 20438 9596 20444 9608
rect 20496 9596 20502 9648
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14240 9472 14841 9500
rect 14240 9460 14246 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 14918 9460 14924 9512
rect 14976 9500 14982 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 14976 9472 15301 9500
rect 14976 9460 14982 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 17218 9500 17224 9512
rect 17175 9472 17224 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 18138 9500 18144 9512
rect 18099 9472 18144 9500
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 19150 9460 19156 9512
rect 19208 9500 19214 9512
rect 21266 9509 21272 9512
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19208 9472 19533 9500
rect 19208 9460 19214 9472
rect 19521 9469 19533 9472
rect 19567 9500 19579 9503
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 19567 9472 19717 9500
rect 19567 9469 19579 9472
rect 19521 9463 19579 9469
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 21244 9503 21272 9509
rect 21244 9469 21256 9503
rect 21324 9500 21330 9512
rect 21637 9503 21695 9509
rect 21637 9500 21649 9503
rect 21324 9472 21649 9500
rect 21244 9463 21272 9469
rect 21266 9460 21272 9463
rect 21324 9460 21330 9472
rect 21637 9469 21649 9472
rect 21683 9469 21695 9503
rect 21637 9463 21695 9469
rect 23658 9460 23664 9512
rect 23716 9509 23722 9512
rect 23716 9503 23754 9509
rect 23742 9500 23754 9503
rect 24121 9503 24179 9509
rect 24121 9500 24133 9503
rect 23742 9472 24133 9500
rect 23742 9469 23754 9472
rect 23716 9463 23754 9469
rect 24121 9469 24133 9472
rect 24167 9469 24179 9503
rect 24121 9463 24179 9469
rect 23716 9460 23722 9463
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 10367 9404 12173 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 12161 9401 12173 9404
rect 12207 9432 12219 9435
rect 13280 9432 13308 9460
rect 15562 9432 15568 9444
rect 12207 9404 13308 9432
rect 15523 9404 15568 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 15562 9392 15568 9404
rect 15620 9392 15626 9444
rect 16301 9435 16359 9441
rect 16301 9401 16313 9435
rect 16347 9432 16359 9435
rect 16577 9435 16635 9441
rect 16577 9432 16589 9435
rect 16347 9404 16589 9432
rect 16347 9401 16359 9404
rect 16301 9395 16359 9401
rect 16577 9401 16589 9404
rect 16623 9401 16635 9435
rect 17862 9432 17868 9444
rect 16577 9395 16635 9401
rect 17236 9404 17868 9432
rect 2148 9364 2176 9392
rect 2958 9364 2964 9376
rect 1688 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 4154 9364 4160 9376
rect 4115 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 5626 9364 5632 9376
rect 5587 9336 5632 9364
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6236 9336 6469 9364
rect 6236 9324 6242 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 6457 9327 6515 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 16592 9364 16620 9395
rect 17236 9364 17264 9404
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 20346 9432 20352 9444
rect 20307 9404 20352 9432
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 17494 9364 17500 9376
rect 16592 9336 17264 9364
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 18288 9336 18337 9364
rect 18288 9324 18294 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 21315 9367 21373 9373
rect 21315 9333 21327 9367
rect 21361 9364 21373 9367
rect 21542 9364 21548 9376
rect 21361 9336 21548 9364
rect 21361 9333 21373 9336
rect 21315 9327 21373 9333
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 23799 9367 23857 9373
rect 23799 9333 23811 9367
rect 23845 9364 23857 9367
rect 24026 9364 24032 9376
rect 23845 9336 24032 9364
rect 23845 9333 23857 9336
rect 23799 9327 23857 9333
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2130 9160 2136 9172
rect 2091 9132 2136 9160
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 3510 9160 3516 9172
rect 3471 9132 3516 9160
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 3936 9132 4629 9160
rect 3936 9120 3942 9132
rect 4617 9129 4629 9132
rect 4663 9160 4675 9163
rect 8205 9163 8263 9169
rect 4663 9132 4844 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 1118 9052 1124 9104
rect 1176 9092 1182 9104
rect 2038 9092 2044 9104
rect 1176 9064 2044 9092
rect 1176 9052 1182 9064
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2593 9095 2651 9101
rect 2593 9092 2605 9095
rect 2556 9064 2605 9092
rect 2556 9052 2562 9064
rect 2593 9061 2605 9064
rect 2639 9092 2651 9095
rect 2774 9092 2780 9104
rect 2639 9064 2780 9092
rect 2639 9061 2651 9064
rect 2593 9055 2651 9061
rect 2774 9052 2780 9064
rect 2832 9052 2838 9104
rect 4816 9033 4844 9132
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8386 9160 8392 9172
rect 8251 9132 8392 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 9640 9132 10425 9160
rect 9640 9120 9646 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10778 9160 10784 9172
rect 10739 9132 10784 9160
rect 10413 9123 10471 9129
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 11422 9160 11428 9172
rect 11383 9132 11428 9160
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 14918 9160 14924 9172
rect 14879 9132 14924 9160
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15746 9160 15752 9172
rect 15707 9132 15752 9160
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 16758 9160 16764 9172
rect 16671 9132 16764 9160
rect 5074 9052 5080 9104
rect 5132 9101 5138 9104
rect 5132 9095 5180 9101
rect 5132 9061 5134 9095
rect 5168 9061 5180 9095
rect 5132 9055 5180 9061
rect 9769 9095 9827 9101
rect 9769 9061 9781 9095
rect 9815 9092 9827 9095
rect 10226 9092 10232 9104
rect 9815 9064 10232 9092
rect 9815 9061 9827 9064
rect 9769 9055 9827 9061
rect 5132 9052 5138 9055
rect 10226 9052 10232 9064
rect 10284 9092 10290 9104
rect 10870 9092 10876 9104
rect 10284 9064 10876 9092
rect 10284 9052 10290 9064
rect 10870 9052 10876 9064
rect 10928 9052 10934 9104
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 11146 9092 11152 9104
rect 11020 9064 11152 9092
rect 11020 9052 11026 9064
rect 11146 9052 11152 9064
rect 11204 9092 11210 9104
rect 11882 9092 11888 9104
rect 11204 9064 11888 9092
rect 11204 9052 11210 9064
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 8993 1522 9027
rect 1464 8987 1522 8993
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 8993 4859 9027
rect 7098 9024 7104 9036
rect 7059 8996 7104 9024
rect 4801 8987 4859 8993
rect 1479 8888 1507 8987
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 11348 9033 11376 9064
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 13446 9052 13452 9104
rect 13504 9092 13510 9104
rect 13633 9095 13691 9101
rect 13633 9092 13645 9095
rect 13504 9064 13645 9092
rect 13504 9052 13510 9064
rect 13633 9061 13645 9064
rect 13679 9092 13691 9095
rect 14090 9092 14096 9104
rect 13679 9064 14096 9092
rect 13679 9061 13691 9064
rect 13633 9055 13691 9061
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 16574 9092 16580 9104
rect 16535 9064 16580 9092
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 16684 9101 16712 9132
rect 16758 9120 16764 9132
rect 16816 9160 16822 9172
rect 18966 9160 18972 9172
rect 16816 9132 18972 9160
rect 16816 9120 16822 9132
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 19150 9160 19156 9172
rect 19111 9132 19156 9160
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 16669 9095 16727 9101
rect 16669 9061 16681 9095
rect 16715 9061 16727 9095
rect 17218 9092 17224 9104
rect 17179 9064 17224 9092
rect 16669 9055 16727 9061
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 18233 9095 18291 9101
rect 18233 9061 18245 9095
rect 18279 9092 18291 9095
rect 18322 9092 18328 9104
rect 18279 9064 18328 9092
rect 18279 9061 18291 9064
rect 18233 9055 18291 9061
rect 18322 9052 18328 9064
rect 18380 9052 18386 9104
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11698 8984 11704 9036
rect 11756 9033 11762 9036
rect 11756 9027 11805 9033
rect 11756 8993 11759 9027
rect 11793 8993 11805 9027
rect 13078 9024 13084 9036
rect 13039 8996 13084 9024
rect 11756 8987 11805 8993
rect 11756 8984 11762 8987
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13354 9024 13360 9036
rect 13315 8996 13360 9024
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 21910 8984 21916 9036
rect 21968 9033 21974 9036
rect 21968 9027 22006 9033
rect 21994 8993 22006 9027
rect 21968 8987 22006 8993
rect 21968 8984 21974 8987
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2682 8956 2688 8968
rect 2547 8928 2688 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 3142 8956 3148 8968
rect 2823 8928 3148 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 2792 8888 2820 8919
rect 3142 8916 3148 8928
rect 3200 8956 3206 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3200 8928 3801 8956
rect 3200 8916 3206 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6328 8928 7021 8956
rect 6328 8916 6334 8928
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8536 8928 8585 8956
rect 8536 8916 8542 8928
rect 8573 8925 8585 8928
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9272 8928 10149 8956
rect 9272 8916 9278 8928
rect 10137 8925 10149 8928
rect 10183 8956 10195 8959
rect 10686 8956 10692 8968
rect 10183 8928 10692 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11020 8928 11253 8956
rect 11020 8916 11026 8928
rect 11241 8925 11253 8928
rect 11287 8956 11299 8959
rect 13722 8956 13728 8968
rect 11287 8928 13728 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 17862 8956 17868 8968
rect 15988 8928 17868 8956
rect 15988 8916 15994 8928
rect 17862 8916 17868 8928
rect 17920 8956 17926 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 17920 8928 18153 8956
rect 17920 8916 17926 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 19610 8956 19616 8968
rect 19571 8928 19616 8956
rect 18417 8919 18475 8925
rect 1479 8860 2820 8888
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 6052 8860 6561 8888
rect 6052 8848 6058 8860
rect 6549 8857 6561 8860
rect 6595 8888 6607 8891
rect 7374 8888 7380 8900
rect 6595 8860 7380 8888
rect 6595 8857 6607 8860
rect 6549 8851 6607 8857
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 9934 8891 9992 8897
rect 9934 8888 9946 8891
rect 9640 8860 9946 8888
rect 9640 8848 9646 8860
rect 9934 8857 9946 8860
rect 9980 8888 9992 8891
rect 11514 8888 11520 8900
rect 9980 8860 11520 8888
rect 9980 8857 9992 8860
rect 9934 8851 9992 8857
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 18432 8888 18460 8919
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 20898 8956 20904 8968
rect 20859 8928 20904 8956
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 18012 8860 18460 8888
rect 18012 8848 18018 8860
rect 1535 8823 1593 8829
rect 1535 8789 1547 8823
rect 1581 8820 1593 8823
rect 1854 8820 1860 8832
rect 1581 8792 1860 8820
rect 1581 8789 1593 8792
rect 1535 8783 1593 8789
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 5721 8823 5779 8829
rect 5721 8820 5733 8823
rect 2096 8792 5733 8820
rect 2096 8780 2102 8792
rect 5721 8789 5733 8792
rect 5767 8789 5779 8823
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 5721 8783 5779 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 9398 8820 9404 8832
rect 9359 8792 9404 8820
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12492 8792 12633 8820
rect 12492 8780 12498 8792
rect 12621 8789 12633 8792
rect 12667 8820 12679 8823
rect 13170 8820 13176 8832
rect 12667 8792 13176 8820
rect 12667 8789 12679 8792
rect 12621 8783 12679 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 14274 8820 14280 8832
rect 14235 8792 14280 8820
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 22002 8780 22008 8832
rect 22060 8829 22066 8832
rect 22060 8823 22109 8829
rect 22060 8789 22063 8823
rect 22097 8820 22109 8823
rect 22097 8792 22153 8820
rect 22097 8789 22109 8792
rect 22060 8783 22109 8789
rect 22060 8780 22066 8783
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2314 8616 2320 8628
rect 1995 8588 2320 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2924 8588 3065 8616
rect 2924 8576 2930 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 6270 8616 6276 8628
rect 5408 8588 6276 8616
rect 5408 8576 5414 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 9306 8616 9312 8628
rect 9267 8588 9312 8616
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9861 8619 9919 8625
rect 9861 8585 9873 8619
rect 9907 8616 9919 8619
rect 10226 8616 10232 8628
rect 9907 8588 10232 8616
rect 9907 8585 9919 8588
rect 9861 8579 9919 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 11054 8616 11060 8628
rect 10551 8588 10916 8616
rect 11015 8588 11060 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10888 8560 10916 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 12894 8616 12900 8628
rect 11808 8588 12900 8616
rect 8386 8508 8392 8560
rect 8444 8548 8450 8560
rect 9122 8548 9128 8560
rect 8444 8520 9128 8548
rect 8444 8508 8450 8520
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 10686 8548 10692 8560
rect 9456 8520 10692 8548
rect 9456 8508 9462 8520
rect 10686 8508 10692 8520
rect 10744 8557 10750 8560
rect 10744 8551 10793 8557
rect 10744 8517 10747 8551
rect 10781 8517 10793 8551
rect 10870 8548 10876 8560
rect 10831 8520 10876 8548
rect 10744 8511 10793 8517
rect 10744 8508 10750 8511
rect 10870 8508 10876 8520
rect 10928 8508 10934 8560
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 4062 8480 4068 8492
rect 3559 8452 4068 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3896 8421 3924 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5442 8480 5448 8492
rect 5307 8452 5448 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5994 8480 6000 8492
rect 5951 8452 6000 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6972 8452 7389 8480
rect 6972 8440 6978 8452
rect 7377 8449 7389 8452
rect 7423 8480 7435 8483
rect 7742 8480 7748 8492
rect 7423 8452 7748 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9214 8480 9220 8492
rect 9079 8452 9220 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 10962 8480 10968 8492
rect 10923 8452 10968 8480
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 4154 8412 4160 8424
rect 4115 8384 4160 8412
rect 3881 8375 3939 8381
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 7116 8384 8309 8412
rect 7116 8356 7144 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 9122 8412 9128 8424
rect 8711 8384 9128 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10778 8412 10784 8424
rect 10643 8384 10784 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8344 2283 8347
rect 2314 8344 2320 8356
rect 2271 8316 2320 8344
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3326 8344 3332 8356
rect 2823 8316 3332 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 3326 8304 3332 8316
rect 3384 8304 3390 8356
rect 4338 8344 4344 8356
rect 4299 8316 4344 8344
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 6641 8347 6699 8353
rect 5408 8316 5453 8344
rect 5408 8304 5414 8316
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 7098 8344 7104 8356
rect 6687 8316 7104 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 7208 8316 7297 8344
rect 7208 8288 7236 8316
rect 7285 8313 7297 8316
rect 7331 8344 7343 8347
rect 7650 8344 7656 8356
rect 7331 8316 7656 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7650 8304 7656 8316
rect 7708 8353 7714 8356
rect 7708 8347 7756 8353
rect 7708 8313 7710 8347
rect 7744 8313 7756 8347
rect 7708 8307 7756 8313
rect 7708 8304 7714 8307
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 11514 8304 11520 8356
rect 11572 8344 11578 8356
rect 11808 8353 11836 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13262 8616 13268 8628
rect 13223 8588 13268 8616
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13722 8616 13728 8628
rect 13683 8588 13728 8616
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 14056 8588 15669 8616
rect 14056 8576 14062 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 12802 8557 12808 8560
rect 12253 8551 12311 8557
rect 12253 8517 12265 8551
rect 12299 8548 12311 8551
rect 12786 8551 12808 8557
rect 12786 8548 12798 8551
rect 12299 8520 12798 8548
rect 12299 8517 12311 8520
rect 12253 8511 12311 8517
rect 12786 8517 12798 8520
rect 12786 8511 12808 8517
rect 12802 8508 12808 8511
rect 12860 8508 12866 8560
rect 12434 8440 12440 8492
rect 12492 8440 12498 8492
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8480 13047 8483
rect 13740 8480 13768 8576
rect 15672 8548 15700 8579
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 16632 8588 17417 8616
rect 16632 8576 16638 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17405 8579 17463 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18322 8576 18328 8628
rect 18380 8616 18386 8628
rect 18509 8619 18567 8625
rect 18509 8616 18521 8619
rect 18380 8588 18521 8616
rect 18380 8576 18386 8588
rect 18509 8585 18521 8588
rect 18555 8585 18567 8619
rect 18509 8579 18567 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20404 8588 20453 8616
rect 20404 8576 20410 8588
rect 20441 8585 20453 8588
rect 20487 8616 20499 8619
rect 20806 8616 20812 8628
rect 20487 8588 20812 8616
rect 20487 8585 20499 8588
rect 20441 8579 20499 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 15746 8548 15752 8560
rect 15659 8520 15752 8548
rect 15746 8508 15752 8520
rect 15804 8548 15810 8560
rect 16758 8548 16764 8560
rect 15804 8520 16205 8548
rect 16719 8520 16764 8548
rect 15804 8508 15810 8520
rect 13035 8452 13768 8480
rect 13035 8449 13047 8452
rect 12989 8443 13047 8449
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15620 8452 15853 8480
rect 15620 8440 15626 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 15841 8443 15899 8449
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 11572 8316 11805 8344
rect 11572 8304 11578 8316
rect 11793 8313 11805 8316
rect 11839 8313 11851 8347
rect 11793 8307 11851 8313
rect 12452 8344 12480 8440
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8412 14151 8415
rect 14182 8412 14188 8424
rect 14139 8384 14188 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14332 8384 14657 8412
rect 14332 8372 14338 8384
rect 14645 8381 14657 8384
rect 14691 8412 14703 8415
rect 14826 8412 14832 8424
rect 14691 8384 14832 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 12452 8316 12633 8344
rect 4893 8279 4951 8285
rect 4893 8245 4905 8279
rect 4939 8276 4951 8279
rect 5074 8276 5080 8288
rect 4939 8248 5080 8276
rect 4939 8245 4951 8248
rect 4893 8239 4951 8245
rect 5074 8236 5080 8248
rect 5132 8276 5138 8288
rect 7190 8276 7196 8288
rect 5132 8248 7196 8276
rect 5132 8236 5138 8248
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 10244 8276 10272 8304
rect 12452 8288 12480 8316
rect 12621 8313 12633 8316
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 16177 8353 16205 8520
rect 16758 8508 16764 8520
rect 16816 8548 16822 8560
rect 17037 8551 17095 8557
rect 17037 8548 17049 8551
rect 16816 8520 17049 8548
rect 16816 8508 16822 8520
rect 17037 8517 17049 8520
rect 17083 8517 17095 8551
rect 17037 8511 17095 8517
rect 18233 8551 18291 8557
rect 18233 8517 18245 8551
rect 18279 8548 18291 8551
rect 18414 8548 18420 8560
rect 18279 8520 18420 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 19705 8551 19763 8557
rect 19705 8517 19717 8551
rect 19751 8548 19763 8551
rect 21266 8548 21272 8560
rect 19751 8520 21272 8548
rect 19751 8517 19763 8520
rect 19705 8511 19763 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 17218 8440 17224 8492
rect 17276 8480 17282 8492
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 17276 8452 19165 8480
rect 17276 8440 17282 8452
rect 19153 8449 19165 8452
rect 19199 8480 19211 8483
rect 19334 8480 19340 8492
rect 19199 8452 19340 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 20714 8480 20720 8492
rect 19668 8452 20720 8480
rect 19668 8440 19674 8452
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 16298 8372 16304 8424
rect 16356 8412 16362 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 16356 8384 18061 8412
rect 16356 8372 16362 8384
rect 18049 8381 18061 8384
rect 18095 8412 18107 8415
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 18095 8384 18889 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18877 8381 18889 8384
rect 18923 8381 18935 8415
rect 18877 8375 18935 8381
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22224 8415 22282 8421
rect 22224 8412 22236 8415
rect 22152 8384 22236 8412
rect 22152 8372 22158 8384
rect 22224 8381 22236 8384
rect 22270 8412 22282 8415
rect 22649 8415 22707 8421
rect 22649 8412 22661 8415
rect 22270 8384 22661 8412
rect 22270 8381 22282 8384
rect 22224 8375 22282 8381
rect 22649 8381 22661 8384
rect 22695 8381 22707 8415
rect 22649 8375 22707 8381
rect 16162 8347 16220 8353
rect 13596 8316 14320 8344
rect 13596 8304 13602 8316
rect 10778 8276 10784 8288
rect 10244 8248 10784 8276
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 12434 8236 12440 8288
rect 12492 8236 12498 8288
rect 14292 8285 14320 8316
rect 16162 8313 16174 8347
rect 16208 8313 16220 8347
rect 16162 8307 16220 8313
rect 19150 8304 19156 8356
rect 19208 8344 19214 8356
rect 19245 8347 19303 8353
rect 19245 8344 19257 8347
rect 19208 8316 19257 8344
rect 19208 8304 19214 8316
rect 19245 8313 19257 8316
rect 19291 8313 19303 8347
rect 19245 8307 19303 8313
rect 20806 8304 20812 8356
rect 20864 8344 20870 8356
rect 20864 8316 20909 8344
rect 20864 8304 20870 8316
rect 21450 8304 21456 8356
rect 21508 8344 21514 8356
rect 21910 8344 21916 8356
rect 21508 8316 21916 8344
rect 21508 8304 21514 8316
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 22327 8347 22385 8353
rect 22327 8313 22339 8347
rect 22373 8344 22385 8347
rect 23290 8344 23296 8356
rect 22373 8316 23296 8344
rect 22373 8313 22385 8316
rect 22327 8307 22385 8313
rect 23290 8304 23296 8316
rect 23348 8304 23354 8356
rect 14277 8279 14335 8285
rect 14277 8245 14289 8279
rect 14323 8245 14335 8279
rect 14277 8239 14335 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 2038 8072 2044 8084
rect 1719 8044 2044 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2740 8044 3157 8072
rect 2740 8032 2746 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3145 8035 3203 8041
rect 3697 8075 3755 8081
rect 3697 8041 3709 8075
rect 3743 8072 3755 8075
rect 4062 8072 4068 8084
rect 3743 8044 4068 8072
rect 3743 8041 3755 8044
rect 3697 8035 3755 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5592 8044 6009 8072
rect 5592 8032 5598 8044
rect 5997 8041 6009 8044
rect 6043 8072 6055 8075
rect 6822 8072 6828 8084
rect 6043 8044 6828 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7742 8072 7748 8084
rect 7703 8044 7748 8072
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9582 8072 9588 8084
rect 9539 8044 9588 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11940 8044 11989 8072
rect 11940 8032 11946 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13412 8044 13553 8072
rect 13412 8032 13418 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 15562 8032 15568 8084
rect 15620 8072 15626 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 15620 8044 15853 8072
rect 15620 8032 15626 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 15841 8035 15899 8041
rect 16684 8044 17601 8072
rect 1578 7964 1584 8016
rect 1636 8004 1642 8016
rect 1857 8007 1915 8013
rect 1857 8004 1869 8007
rect 1636 7976 1869 8004
rect 1636 7964 1642 7976
rect 1857 7973 1869 7976
rect 1903 7973 1915 8007
rect 1857 7967 1915 7973
rect 1949 8007 2007 8013
rect 1949 7973 1961 8007
rect 1995 8004 2007 8007
rect 2222 8004 2228 8016
rect 1995 7976 2228 8004
rect 1995 7973 2007 7976
rect 1949 7967 2007 7973
rect 2222 7964 2228 7976
rect 2280 7964 2286 8016
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 5074 8013 5080 8016
rect 5071 8004 5080 8013
rect 2832 7976 2877 8004
rect 5035 7976 5080 8004
rect 2832 7964 2838 7976
rect 5071 7967 5080 7976
rect 5074 7964 5080 7967
rect 5132 7964 5138 8016
rect 7193 8007 7251 8013
rect 7193 7973 7205 8007
rect 7239 8004 7251 8007
rect 7561 8007 7619 8013
rect 7561 8004 7573 8007
rect 7239 7976 7573 8004
rect 7239 7973 7251 7976
rect 7193 7967 7251 7973
rect 7561 7973 7573 7976
rect 7607 8004 7619 8007
rect 9306 8004 9312 8016
rect 7607 7976 9312 8004
rect 7607 7973 7619 7976
rect 7561 7967 7619 7973
rect 8220 7948 8248 7976
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 8004 10011 8007
rect 10042 8004 10048 8016
rect 9999 7976 10048 8004
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 10042 7964 10048 7976
rect 10100 8004 10106 8016
rect 12161 8007 12219 8013
rect 12161 8004 12173 8007
rect 10100 7976 12173 8004
rect 10100 7964 10106 7976
rect 12161 7973 12173 7976
rect 12207 7973 12219 8007
rect 13372 8004 13400 8032
rect 16684 8016 16712 8044
rect 17589 8041 17601 8044
rect 17635 8041 17647 8075
rect 17589 8035 17647 8041
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19150 8072 19156 8084
rect 19107 8044 19156 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 19334 8072 19340 8084
rect 19295 8044 19340 8072
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19705 8075 19763 8081
rect 19705 8072 19717 8075
rect 19484 8044 19717 8072
rect 19484 8032 19490 8044
rect 19705 8041 19717 8044
rect 19751 8041 19763 8075
rect 20714 8072 20720 8084
rect 20675 8044 20720 8072
rect 19705 8035 19763 8041
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 16666 8004 16672 8016
rect 12161 7967 12219 7973
rect 12268 7976 13400 8004
rect 16627 7976 16672 8004
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 4890 7936 4896 7948
rect 4755 7908 4896 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 6454 7936 6460 7948
rect 6415 7908 6460 7936
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 7926 7936 7932 7948
rect 7887 7908 7932 7936
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8202 7936 8208 7948
rect 8115 7908 8208 7936
rect 8202 7896 8208 7908
rect 8260 7936 8266 7948
rect 8481 7939 8539 7945
rect 8260 7908 8285 7936
rect 8260 7896 8266 7908
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8570 7936 8576 7948
rect 8527 7908 8576 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 10778 7936 10784 7948
rect 10643 7908 10784 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 2498 7868 2504 7880
rect 2459 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 8294 7868 8300 7880
rect 3292 7840 8300 7868
rect 3292 7828 3298 7840
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7868 10563 7871
rect 10962 7868 10968 7880
rect 10551 7840 10968 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11698 7868 11704 7880
rect 11611 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7868 11762 7880
rect 12268 7868 12296 7976
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 16761 8007 16819 8013
rect 16761 7973 16773 8007
rect 16807 8004 16819 8007
rect 16850 8004 16856 8016
rect 16807 7976 16856 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 16850 7964 16856 7976
rect 16908 7964 16914 8016
rect 17313 8007 17371 8013
rect 17313 7973 17325 8007
rect 17359 8004 17371 8007
rect 17954 8004 17960 8016
rect 17359 7976 17960 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 18414 7964 18420 8016
rect 18472 8013 18478 8016
rect 18472 8007 18520 8013
rect 18472 7973 18474 8007
rect 18508 7973 18520 8007
rect 18472 7967 18520 7973
rect 18472 7964 18478 7967
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 11756 7840 12296 7868
rect 11756 7828 11762 7840
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 2682 7800 2688 7812
rect 2464 7772 2688 7800
rect 2464 7760 2470 7772
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 6641 7803 6699 7809
rect 6641 7800 6653 7803
rect 2792 7772 6653 7800
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 2792 7732 2820 7772
rect 6641 7769 6653 7772
rect 6687 7769 6699 7803
rect 6641 7763 6699 7769
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 10042 7800 10048 7812
rect 9916 7772 10048 7800
rect 9916 7760 9922 7772
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 10686 7760 10692 7812
rect 10744 7809 10750 7812
rect 10744 7803 10793 7809
rect 10744 7769 10747 7803
rect 10781 7769 10793 7803
rect 10870 7800 10876 7812
rect 10831 7772 10876 7800
rect 10744 7763 10793 7769
rect 10744 7760 10750 7763
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 11054 7800 11060 7812
rect 11015 7772 11060 7800
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12820 7800 12848 7899
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 16298 7936 16304 7948
rect 12952 7908 16304 7936
rect 12952 7896 12958 7908
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 20990 7936 20996 7948
rect 20951 7908 20996 7936
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 22462 7936 22468 7948
rect 22423 7908 22468 7936
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 23566 7945 23572 7948
rect 23544 7939 23572 7945
rect 23544 7905 23556 7939
rect 23544 7899 23572 7905
rect 23566 7896 23572 7899
rect 23624 7896 23630 7948
rect 13354 7828 13360 7880
rect 13412 7868 13418 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13412 7840 13737 7868
rect 13412 7828 13418 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 13725 7831 13783 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16850 7868 16856 7880
rect 16531 7840 16856 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 18138 7868 18144 7880
rect 18099 7840 18144 7868
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 17034 7800 17040 7812
rect 12400 7772 17040 7800
rect 12400 7760 12406 7772
rect 17034 7760 17040 7772
rect 17092 7760 17098 7812
rect 1912 7704 2820 7732
rect 1912 7692 1918 7704
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5629 7735 5687 7741
rect 5629 7732 5641 7735
rect 5592 7704 5641 7732
rect 5592 7692 5598 7704
rect 5629 7701 5641 7704
rect 5675 7701 5687 7735
rect 10704 7732 10732 7760
rect 11238 7732 11244 7744
rect 10704 7704 11244 7732
rect 5629 7695 5687 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 13170 7732 13176 7744
rect 13131 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 14274 7732 14280 7744
rect 14235 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 21266 7692 21272 7744
rect 21324 7732 21330 7744
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 21324 7704 21925 7732
rect 21324 7692 21330 7704
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 21913 7695 21971 7701
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22649 7735 22707 7741
rect 22649 7732 22661 7735
rect 22244 7704 22661 7732
rect 22244 7692 22250 7704
rect 22649 7701 22661 7704
rect 22695 7701 22707 7735
rect 22649 7695 22707 7701
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 23615 7735 23673 7741
rect 23615 7732 23627 7735
rect 23440 7704 23627 7732
rect 23440 7692 23446 7704
rect 23615 7701 23627 7704
rect 23661 7701 23673 7735
rect 23615 7695 23673 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 2222 7528 2228 7540
rect 1903 7500 2228 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 3513 7531 3571 7537
rect 3513 7528 3525 7531
rect 2424 7500 3525 7528
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 2424 7460 2452 7500
rect 3513 7497 3525 7500
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5905 7531 5963 7537
rect 5905 7528 5917 7531
rect 4948 7500 5917 7528
rect 4948 7488 4954 7500
rect 5905 7497 5917 7500
rect 5951 7497 5963 7531
rect 5905 7491 5963 7497
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9398 7528 9404 7540
rect 9079 7500 9404 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 10870 7528 10876 7540
rect 10735 7500 10876 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 10870 7488 10876 7500
rect 10928 7528 10934 7540
rect 12253 7531 12311 7537
rect 12253 7528 12265 7531
rect 10928 7500 12265 7528
rect 10928 7488 10934 7500
rect 12253 7497 12265 7500
rect 12299 7528 12311 7531
rect 12342 7528 12348 7540
rect 12299 7500 12348 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 12802 7528 12808 7540
rect 12759 7500 12808 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 13357 7531 13415 7537
rect 13357 7497 13369 7531
rect 13403 7528 13415 7531
rect 13446 7528 13452 7540
rect 13403 7500 13452 7528
rect 13403 7497 13415 7500
rect 13357 7491 13415 7497
rect 1636 7432 2452 7460
rect 1636 7420 1642 7432
rect 2498 7420 2504 7472
rect 2556 7460 2562 7472
rect 2777 7463 2835 7469
rect 2777 7460 2789 7463
rect 2556 7432 2789 7460
rect 2556 7420 2562 7432
rect 2777 7429 2789 7432
rect 2823 7429 2835 7463
rect 2777 7423 2835 7429
rect 3694 7420 3700 7472
rect 3752 7420 3758 7472
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 5074 7460 5080 7472
rect 4663 7432 5080 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 10778 7460 10784 7472
rect 10367 7432 10784 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 10778 7420 10784 7432
rect 10836 7460 10842 7472
rect 11054 7460 11060 7472
rect 10836 7432 11060 7460
rect 10836 7420 10842 7432
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7392 2283 7395
rect 2271 7364 3280 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 1394 7216 1400 7268
rect 1452 7256 1458 7268
rect 2222 7256 2228 7268
rect 1452 7228 2228 7256
rect 1452 7216 1458 7228
rect 2222 7216 2228 7228
rect 2280 7256 2286 7268
rect 3252 7265 3280 7364
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3712 7392 3740 7420
rect 3568 7364 4108 7392
rect 3568 7352 3574 7364
rect 3748 7327 3806 7333
rect 3748 7293 3760 7327
rect 3794 7324 3806 7327
rect 4080 7324 4108 7364
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4396 7364 4721 7392
rect 4396 7352 4402 7364
rect 4709 7361 4721 7364
rect 4755 7392 4767 7395
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 4755 7364 6285 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 6273 7361 6285 7364
rect 6319 7361 6331 7395
rect 6273 7355 6331 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11422 7392 11428 7404
rect 11195 7364 11428 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11422 7352 11428 7364
rect 11480 7392 11486 7404
rect 12894 7392 12900 7404
rect 11480 7364 12900 7392
rect 11480 7352 11486 7364
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 3794 7296 4016 7324
rect 4080 7296 5641 7324
rect 3794 7293 3806 7296
rect 3748 7287 3806 7293
rect 2317 7259 2375 7265
rect 2317 7256 2329 7259
rect 2280 7228 2329 7256
rect 2280 7216 2286 7228
rect 2317 7225 2329 7228
rect 2363 7225 2375 7259
rect 2317 7219 2375 7225
rect 3237 7259 3295 7265
rect 3237 7225 3249 7259
rect 3283 7256 3295 7259
rect 3835 7259 3893 7265
rect 3835 7256 3847 7259
rect 3283 7228 3847 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 3835 7225 3847 7228
rect 3881 7225 3893 7259
rect 3835 7219 3893 7225
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 3988 7188 4016 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 7147 7296 7481 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7469 7293 7481 7296
rect 7515 7324 7527 7327
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7515 7296 7849 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 7837 7293 7849 7296
rect 7883 7324 7895 7327
rect 7926 7324 7932 7336
rect 7883 7296 7932 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8202 7324 8208 7336
rect 8163 7296 8208 7324
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7324 8447 7327
rect 8662 7324 8668 7336
rect 8435 7296 8668 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 9528 7327 9586 7333
rect 9528 7324 9540 7327
rect 8812 7296 9540 7324
rect 8812 7284 8818 7296
rect 9528 7293 9540 7296
rect 9574 7293 9586 7327
rect 9528 7287 9586 7293
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 11054 7324 11060 7336
rect 10827 7296 11060 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 5074 7265 5080 7268
rect 5071 7256 5080 7265
rect 5035 7228 5080 7256
rect 5071 7219 5080 7228
rect 5074 7216 5080 7219
rect 5132 7216 5138 7268
rect 9401 7259 9459 7265
rect 9401 7225 9413 7259
rect 9447 7256 9459 7259
rect 10796 7256 10824 7287
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7324 11575 7327
rect 12621 7327 12679 7333
rect 12621 7324 12633 7327
rect 11563 7296 12633 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 12621 7293 12633 7296
rect 12667 7324 12679 7327
rect 13372 7324 13400 7491
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 16850 7528 16856 7540
rect 16811 7500 16856 7528
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21434 7531 21492 7537
rect 21434 7528 21446 7531
rect 20772 7500 21446 7528
rect 20772 7488 20778 7500
rect 21434 7497 21446 7500
rect 21480 7528 21492 7531
rect 22281 7531 22339 7537
rect 22281 7528 22293 7531
rect 21480 7500 22293 7528
rect 21480 7497 21492 7500
rect 21434 7491 21492 7497
rect 22281 7497 22293 7500
rect 22327 7497 22339 7531
rect 22281 7491 22339 7497
rect 22462 7488 22468 7540
rect 22520 7528 22526 7540
rect 22649 7531 22707 7537
rect 22649 7528 22661 7531
rect 22520 7500 22661 7528
rect 22520 7488 22526 7500
rect 22649 7497 22661 7500
rect 22695 7497 22707 7531
rect 22649 7491 22707 7497
rect 21545 7463 21603 7469
rect 21545 7460 21557 7463
rect 21100 7432 21557 7460
rect 21100 7404 21128 7432
rect 21545 7429 21557 7432
rect 21591 7460 21603 7463
rect 21591 7432 23704 7460
rect 21591 7429 21603 7432
rect 21545 7423 21603 7429
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 14182 7392 14188 7404
rect 13771 7364 14188 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 14108 7333 14136 7364
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7392 15531 7395
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 15519 7364 15945 7392
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 15933 7361 15945 7364
rect 15979 7392 15991 7395
rect 16482 7392 16488 7404
rect 15979 7364 16488 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 18138 7352 18144 7404
rect 18196 7392 18202 7404
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18196 7364 18797 7392
rect 18196 7352 18202 7364
rect 18785 7361 18797 7364
rect 18831 7392 18843 7395
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18831 7364 19073 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19797 7395 19855 7401
rect 19797 7392 19809 7395
rect 19484 7364 19809 7392
rect 19484 7352 19490 7364
rect 19797 7361 19809 7364
rect 19843 7361 19855 7395
rect 21082 7392 21088 7404
rect 21043 7364 21088 7392
rect 19797 7355 19855 7361
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 21726 7392 21732 7404
rect 21687 7364 21732 7392
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 23566 7392 23572 7404
rect 23523 7364 23572 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 23566 7352 23572 7364
rect 23624 7352 23630 7404
rect 12667 7296 13400 7324
rect 14093 7327 14151 7333
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14274 7324 14280 7336
rect 14235 7296 14280 7324
rect 14093 7287 14151 7293
rect 9447 7228 10824 7256
rect 9447 7225 9459 7228
rect 9401 7219 9459 7225
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 11532 7256 11560 7287
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 14700 7296 18061 7324
rect 14700 7284 14706 7296
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18322 7324 18328 7336
rect 18095 7296 18328 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7324 20499 7327
rect 20714 7324 20720 7336
rect 20487 7296 20720 7324
rect 20487 7293 20499 7296
rect 20441 7287 20499 7293
rect 11882 7256 11888 7268
rect 11020 7228 11560 7256
rect 11795 7228 11888 7256
rect 11020 7216 11026 7228
rect 11882 7216 11888 7228
rect 11940 7256 11946 7268
rect 12437 7259 12495 7265
rect 12437 7256 12449 7259
rect 11940 7228 12449 7256
rect 11940 7216 11946 7228
rect 12437 7225 12449 7228
rect 12483 7256 12495 7259
rect 13722 7256 13728 7268
rect 12483 7228 13728 7256
rect 12483 7225 12495 7228
rect 12437 7219 12495 7225
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 15746 7216 15752 7268
rect 15804 7256 15810 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 15804 7228 15853 7256
rect 15804 7216 15810 7228
rect 15841 7225 15853 7228
rect 15887 7256 15899 7259
rect 16295 7259 16353 7265
rect 16295 7256 16307 7259
rect 15887 7228 16307 7256
rect 15887 7225 15899 7228
rect 15841 7219 15899 7225
rect 16295 7225 16307 7228
rect 16341 7225 16353 7259
rect 16295 7219 16353 7225
rect 4157 7191 4215 7197
rect 4157 7188 4169 7191
rect 3200 7160 4169 7188
rect 3200 7148 3206 7160
rect 4157 7157 4169 7160
rect 4203 7157 4215 7191
rect 7650 7188 7656 7200
rect 7611 7160 7656 7188
rect 4157 7151 4215 7157
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 9631 7191 9689 7197
rect 9631 7188 9643 7191
rect 9180 7160 9643 7188
rect 9180 7148 9186 7160
rect 9631 7157 9643 7160
rect 9677 7157 9689 7191
rect 9631 7151 9689 7157
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 13872 7160 13921 7188
rect 13872 7148 13878 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 16316 7188 16344 7219
rect 17402 7216 17408 7268
rect 17460 7256 17466 7268
rect 18524 7256 18552 7287
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 21266 7324 21272 7336
rect 21227 7296 21272 7324
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 23676 7333 23704 7432
rect 21608 7327 21666 7333
rect 21608 7324 21620 7327
rect 21376 7296 21620 7324
rect 17460 7228 18552 7256
rect 19889 7259 19947 7265
rect 17460 7216 17466 7228
rect 19889 7225 19901 7259
rect 19935 7256 19947 7259
rect 19978 7256 19984 7268
rect 19935 7228 19984 7256
rect 19935 7225 19947 7228
rect 19889 7219 19947 7225
rect 16482 7188 16488 7200
rect 16316 7160 16488 7188
rect 13909 7151 13967 7157
rect 16482 7148 16488 7160
rect 16540 7188 16546 7200
rect 17865 7191 17923 7197
rect 17865 7188 17877 7191
rect 16540 7160 17877 7188
rect 16540 7148 16546 7160
rect 17865 7157 17877 7160
rect 17911 7188 17923 7191
rect 18414 7188 18420 7200
rect 17911 7160 18420 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 19613 7191 19671 7197
rect 19613 7157 19625 7191
rect 19659 7188 19671 7191
rect 19904 7188 19932 7219
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 20809 7259 20867 7265
rect 20809 7225 20821 7259
rect 20855 7256 20867 7259
rect 21174 7256 21180 7268
rect 20855 7228 21180 7256
rect 20855 7225 20867 7228
rect 20809 7219 20867 7225
rect 21174 7216 21180 7228
rect 21232 7256 21238 7268
rect 21376 7256 21404 7296
rect 21608 7293 21620 7296
rect 21654 7293 21666 7327
rect 21608 7287 21666 7293
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7324 23719 7327
rect 24121 7327 24179 7333
rect 24121 7324 24133 7327
rect 23707 7296 24133 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 24121 7293 24133 7296
rect 24167 7293 24179 7327
rect 24121 7287 24179 7293
rect 24670 7284 24676 7336
rect 24728 7333 24734 7336
rect 24728 7327 24766 7333
rect 24754 7324 24766 7327
rect 25133 7327 25191 7333
rect 25133 7324 25145 7327
rect 24754 7296 25145 7324
rect 24754 7293 24766 7296
rect 24728 7287 24766 7293
rect 25133 7293 25145 7296
rect 25179 7293 25191 7327
rect 25133 7287 25191 7293
rect 24728 7284 24734 7287
rect 21232 7228 21404 7256
rect 21232 7216 21238 7228
rect 19659 7160 19932 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 23474 7148 23480 7200
rect 23532 7188 23538 7200
rect 23845 7191 23903 7197
rect 23845 7188 23857 7191
rect 23532 7160 23857 7188
rect 23532 7148 23538 7160
rect 23845 7157 23857 7160
rect 23891 7157 23903 7191
rect 23845 7151 23903 7157
rect 24762 7148 24768 7200
rect 24820 7197 24826 7200
rect 24820 7191 24869 7197
rect 24820 7157 24823 7191
rect 24857 7157 24869 7191
rect 24820 7151 24869 7157
rect 24820 7148 24826 7151
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2593 6987 2651 6993
rect 2593 6984 2605 6987
rect 2280 6956 2605 6984
rect 2280 6944 2286 6956
rect 2593 6953 2605 6956
rect 2639 6953 2651 6987
rect 2593 6947 2651 6953
rect 4801 6987 4859 6993
rect 4801 6953 4813 6987
rect 4847 6984 4859 6987
rect 5074 6984 5080 6996
rect 4847 6956 5080 6984
rect 4847 6953 4859 6956
rect 4801 6947 4859 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6454 6984 6460 6996
rect 6415 6956 6460 6984
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 8570 6944 8576 6996
rect 8628 6944 8634 6996
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 8812 6956 9413 6984
rect 8812 6944 8818 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9401 6947 9459 6953
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17460 6956 17509 6984
rect 17460 6944 17466 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 18141 6987 18199 6993
rect 18141 6953 18153 6987
rect 18187 6984 18199 6987
rect 18322 6984 18328 6996
rect 18187 6956 18328 6984
rect 18187 6953 18199 6956
rect 18141 6947 18199 6953
rect 18322 6944 18328 6956
rect 18380 6984 18386 6996
rect 19242 6984 19248 6996
rect 18380 6956 19248 6984
rect 18380 6944 18386 6956
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 19521 6987 19579 6993
rect 19521 6953 19533 6987
rect 19567 6984 19579 6987
rect 19978 6984 19984 6996
rect 19567 6956 19984 6984
rect 19567 6953 19579 6956
rect 19521 6947 19579 6953
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 20990 6984 20996 6996
rect 20763 6956 20996 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 20990 6944 20996 6956
rect 21048 6984 21054 6996
rect 21174 6984 21180 6996
rect 21048 6956 21180 6984
rect 21048 6944 21054 6956
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 1670 6876 1676 6928
rect 1728 6916 1734 6928
rect 1765 6919 1823 6925
rect 1765 6916 1777 6919
rect 1728 6888 1777 6916
rect 1728 6876 1734 6888
rect 1765 6885 1777 6888
rect 1811 6916 1823 6919
rect 7098 6916 7104 6928
rect 1811 6888 2360 6916
rect 7059 6888 7104 6916
rect 1811 6885 1823 6888
rect 1765 6879 1823 6885
rect 2332 6848 2360 6888
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 8588 6916 8616 6944
rect 8220 6888 8616 6916
rect 13556 6888 13768 6916
rect 2682 6848 2688 6860
rect 2332 6820 2688 6848
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 5169 6851 5227 6857
rect 5169 6848 5181 6851
rect 4396 6820 5181 6848
rect 4396 6808 4402 6820
rect 5169 6817 5181 6820
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6270 6848 6276 6860
rect 5675 6820 6276 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8220 6848 8248 6888
rect 8067 6820 8248 6848
rect 8532 6851 8590 6857
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8532 6817 8544 6851
rect 8578 6848 8590 6851
rect 9674 6848 9680 6860
rect 8578 6820 8800 6848
rect 9635 6820 9680 6848
rect 8578 6817 8590 6820
rect 8532 6811 8590 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2498 6780 2504 6792
rect 1719 6752 2504 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 4948 6752 5733 6780
rect 4948 6740 4954 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7374 6780 7380 6792
rect 7335 6752 7380 6780
rect 7009 6743 7067 6749
rect 2222 6712 2228 6724
rect 2183 6684 2228 6712
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 4028 6684 4261 6712
rect 4028 6672 4034 6684
rect 4249 6681 4261 6684
rect 4295 6681 4307 6715
rect 4249 6675 4307 6681
rect 6825 6715 6883 6721
rect 6825 6681 6837 6715
rect 6871 6712 6883 6715
rect 7024 6712 7052 6743
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 8619 6783 8677 6789
rect 8619 6749 8631 6783
rect 8665 6749 8677 6783
rect 8619 6743 8677 6749
rect 7282 6712 7288 6724
rect 6871 6684 7288 6712
rect 6871 6681 6883 6684
rect 6825 6675 6883 6681
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 8634 6712 8662 6743
rect 8772 6724 8800 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 10318 6848 10324 6860
rect 10279 6820 10324 6848
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 10962 6848 10968 6860
rect 10919 6820 10968 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11112 6820 11621 6848
rect 11112 6808 11118 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11882 6848 11888 6860
rect 11843 6820 11888 6848
rect 11609 6811 11667 6817
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 12676 6820 13093 6848
rect 12676 6808 12682 6820
rect 13081 6817 13093 6820
rect 13127 6848 13139 6851
rect 13446 6848 13452 6860
rect 13127 6820 13452 6848
rect 13127 6817 13139 6820
rect 13081 6811 13139 6817
rect 13446 6808 13452 6820
rect 13504 6848 13510 6860
rect 13556 6848 13584 6888
rect 13504 6820 13584 6848
rect 13633 6851 13691 6857
rect 13504 6808 13510 6820
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13740 6848 13768 6888
rect 14826 6876 14832 6928
rect 14884 6916 14890 6928
rect 14884 6888 15608 6916
rect 14884 6876 14890 6888
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 13740 6820 15301 6848
rect 13633 6811 13691 6817
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 15470 6848 15476 6860
rect 15335 6820 15476 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12802 6780 12808 6792
rect 12492 6752 12808 6780
rect 12492 6740 12498 6752
rect 12802 6740 12808 6752
rect 12860 6780 12866 6792
rect 13648 6780 13676 6811
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15580 6848 15608 6888
rect 18414 6876 18420 6928
rect 18472 6916 18478 6928
rect 18922 6919 18980 6925
rect 18922 6916 18934 6919
rect 18472 6888 18934 6916
rect 18472 6876 18478 6888
rect 18922 6885 18934 6888
rect 18968 6916 18980 6919
rect 19058 6916 19064 6928
rect 18968 6888 19064 6916
rect 18968 6885 18980 6888
rect 18922 6879 18980 6885
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 21082 6916 21088 6928
rect 20995 6888 21088 6916
rect 21082 6876 21088 6888
rect 21140 6916 21146 6928
rect 21140 6888 21680 6916
rect 21140 6876 21146 6888
rect 15580 6820 15792 6848
rect 12860 6752 13676 6780
rect 12860 6740 12866 6752
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14001 6783 14059 6789
rect 14001 6780 14013 6783
rect 13780 6752 14013 6780
rect 13780 6740 13786 6752
rect 14001 6749 14013 6752
rect 14047 6749 14059 6783
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 14001 6743 14059 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15764 6789 15792 6820
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16264 6820 16313 6848
rect 16264 6808 16270 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 16301 6811 16359 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 21652 6848 21680 6888
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 21652 6820 22477 6848
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 22554 6808 22560 6860
rect 22612 6848 22618 6860
rect 22612 6820 22657 6848
rect 22612 6808 22618 6820
rect 23934 6808 23940 6860
rect 23992 6848 23998 6860
rect 24029 6851 24087 6857
rect 24029 6848 24041 6851
rect 23992 6820 24041 6848
rect 23992 6808 23998 6820
rect 24029 6817 24041 6820
rect 24075 6817 24087 6851
rect 24029 6811 24087 6817
rect 25200 6851 25258 6857
rect 25200 6817 25212 6851
rect 25246 6848 25258 6851
rect 25498 6848 25504 6860
rect 25246 6820 25504 6848
rect 25246 6817 25258 6820
rect 25200 6811 25258 6817
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6780 15807 6783
rect 16390 6780 16396 6792
rect 15795 6752 16396 6780
rect 15795 6749 15807 6752
rect 15749 6743 15807 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 17218 6780 17224 6792
rect 17179 6752 17224 6780
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 18601 6783 18659 6789
rect 18601 6749 18613 6783
rect 18647 6780 18659 6783
rect 20990 6780 20996 6792
rect 18647 6752 19932 6780
rect 20951 6752 20996 6780
rect 18647 6749 18659 6752
rect 18601 6743 18659 6749
rect 7392 6684 8662 6712
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 7392 6644 7420 6684
rect 8754 6672 8760 6724
rect 8812 6672 8818 6724
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 12452 6684 15577 6712
rect 12452 6656 12480 6684
rect 15565 6681 15577 6684
rect 15611 6712 15623 6715
rect 15838 6712 15844 6724
rect 15611 6684 15844 6712
rect 15611 6681 15623 6684
rect 15565 6675 15623 6681
rect 15838 6672 15844 6684
rect 15896 6712 15902 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 15896 6684 16681 6712
rect 15896 6672 15902 6684
rect 16669 6681 16681 6684
rect 16715 6712 16727 6715
rect 17129 6715 17187 6721
rect 17129 6712 17141 6715
rect 16715 6684 17141 6712
rect 16715 6681 16727 6684
rect 16669 6675 16727 6681
rect 17129 6681 17141 6684
rect 17175 6681 17187 6715
rect 17129 6675 17187 6681
rect 19904 6656 19932 6752
rect 20990 6740 20996 6752
rect 21048 6740 21054 6792
rect 21269 6783 21327 6789
rect 21269 6749 21281 6783
rect 21315 6780 21327 6783
rect 22094 6780 22100 6792
rect 21315 6752 22100 6780
rect 21315 6749 21327 6752
rect 21269 6743 21327 6749
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 21284 6712 21312 6743
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 20772 6684 21312 6712
rect 20772 6672 20778 6684
rect 3016 6616 7420 6644
rect 8389 6647 8447 6653
rect 3016 6604 3022 6616
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8570 6644 8576 6656
rect 8435 6616 8576 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 11514 6644 11520 6656
rect 11475 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6644 11578 6656
rect 12434 6644 12440 6656
rect 11572 6616 12440 6644
rect 11572 6604 11578 6616
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6644 13694 6656
rect 13771 6647 13829 6653
rect 13771 6644 13783 6647
rect 13688 6616 13783 6644
rect 13688 6604 13694 6616
rect 13771 6613 13783 6616
rect 13817 6613 13829 6647
rect 13771 6607 13829 6613
rect 13909 6647 13967 6653
rect 13909 6613 13921 6647
rect 13955 6644 13967 6647
rect 13998 6644 14004 6656
rect 13955 6616 14004 6644
rect 13955 6613 13967 6616
rect 13909 6607 13967 6613
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14274 6644 14280 6656
rect 14235 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 14826 6644 14832 6656
rect 14783 6616 14832 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15454 6647 15512 6653
rect 15454 6613 15466 6647
rect 15500 6644 15512 6647
rect 17018 6647 17076 6653
rect 17018 6644 17030 6647
rect 15500 6616 17030 6644
rect 15500 6613 15512 6616
rect 15454 6607 15512 6613
rect 17018 6613 17030 6616
rect 17064 6644 17076 6647
rect 17402 6644 17408 6656
rect 17064 6616 17408 6644
rect 17064 6613 17076 6616
rect 17018 6607 17076 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 18104 6616 18429 6644
rect 18104 6604 18110 6616
rect 18417 6613 18429 6616
rect 18463 6613 18475 6647
rect 19886 6644 19892 6656
rect 19847 6616 19892 6644
rect 18417 6607 18475 6613
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21913 6647 21971 6653
rect 21913 6644 21925 6647
rect 21324 6616 21925 6644
rect 21324 6604 21330 6616
rect 21913 6613 21925 6616
rect 21959 6613 21971 6647
rect 21913 6607 21971 6613
rect 23842 6604 23848 6656
rect 23900 6644 23906 6656
rect 24213 6647 24271 6653
rect 24213 6644 24225 6647
rect 23900 6616 24225 6644
rect 23900 6604 23906 6616
rect 24213 6613 24225 6616
rect 24259 6613 24271 6647
rect 24213 6607 24271 6613
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 25271 6647 25329 6653
rect 25271 6644 25283 6647
rect 25188 6616 25283 6644
rect 25188 6604 25194 6616
rect 25271 6613 25283 6616
rect 25317 6613 25329 6647
rect 25271 6607 25329 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 5074 6440 5080 6452
rect 4939 6412 5080 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 7190 6440 7196 6452
rect 7151 6412 7196 6440
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 10226 6440 10232 6452
rect 9815 6412 10232 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 11882 6440 11888 6452
rect 11747 6412 11888 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 12492 6412 12725 6440
rect 12492 6400 12498 6412
rect 12713 6409 12725 6412
rect 12759 6409 12771 6443
rect 17589 6443 17647 6449
rect 17589 6440 17601 6443
rect 12713 6403 12771 6409
rect 12912 6412 17601 6440
rect 2593 6375 2651 6381
rect 2593 6341 2605 6375
rect 2639 6372 2651 6375
rect 2682 6372 2688 6384
rect 2639 6344 2688 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 5902 6372 5908 6384
rect 5863 6344 5908 6372
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 10321 6375 10379 6381
rect 10321 6341 10333 6375
rect 10367 6372 10379 6375
rect 10778 6372 10784 6384
rect 10367 6344 10784 6372
rect 10367 6341 10379 6344
rect 10321 6335 10379 6341
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 6641 6307 6699 6313
rect 3660 6276 6592 6304
rect 3660 6264 3666 6276
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3694 6236 3700 6248
rect 3375 6208 3700 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4706 6236 4712 6248
rect 4203 6208 4712 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4706 6196 4712 6208
rect 4764 6236 4770 6248
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4764 6208 4997 6236
rect 4764 6196 4770 6208
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 6564 6236 6592 6276
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 6687 6276 7297 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7285 6273 7297 6276
rect 7331 6304 7343 6307
rect 7650 6304 7656 6316
rect 7331 6276 7656 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 6564 6208 8493 6236
rect 4985 6199 5043 6205
rect 8481 6205 8493 6208
rect 8527 6236 8539 6239
rect 8754 6236 8760 6248
rect 8527 6208 8760 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 10428 6245 10456 6344
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 11606 6332 11612 6384
rect 11664 6372 11670 6384
rect 11790 6372 11796 6384
rect 11664 6344 11796 6372
rect 11664 6332 11670 6344
rect 11790 6332 11796 6344
rect 11848 6372 11854 6384
rect 12253 6375 12311 6381
rect 12253 6372 12265 6375
rect 11848 6344 12265 6372
rect 11848 6332 11854 6344
rect 12253 6341 12265 6344
rect 12299 6372 12311 6375
rect 12912 6372 12940 6412
rect 17589 6409 17601 6412
rect 17635 6409 17647 6443
rect 17589 6403 17647 6409
rect 17770 6400 17776 6452
rect 17828 6440 17834 6452
rect 18506 6440 18512 6452
rect 17828 6412 18512 6440
rect 17828 6400 17834 6412
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19300 6412 19441 6440
rect 19300 6400 19306 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 20993 6443 21051 6449
rect 20993 6409 21005 6443
rect 21039 6440 21051 6443
rect 21082 6440 21088 6452
rect 21039 6412 21088 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 21342 6443 21400 6449
rect 21342 6440 21354 6443
rect 21192 6412 21354 6440
rect 12299 6344 12940 6372
rect 12299 6341 12311 6344
rect 12253 6335 12311 6341
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12820 6313 12848 6344
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 14277 6375 14335 6381
rect 14277 6372 14289 6375
rect 14056 6344 14289 6372
rect 14056 6332 14062 6344
rect 14277 6341 14289 6344
rect 14323 6372 14335 6375
rect 14458 6372 14464 6384
rect 14323 6344 14464 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 14458 6332 14464 6344
rect 14516 6372 14522 6384
rect 14826 6372 14832 6384
rect 14516 6344 14832 6372
rect 14516 6332 14522 6344
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 17218 6372 17224 6384
rect 15672 6344 17224 6372
rect 15672 6316 15700 6344
rect 17218 6332 17224 6344
rect 17276 6372 17282 6384
rect 17405 6375 17463 6381
rect 17405 6372 17417 6375
rect 17276 6344 17417 6372
rect 17276 6332 17282 6344
rect 17405 6341 17417 6344
rect 17451 6341 17463 6375
rect 17405 6335 17463 6341
rect 17865 6375 17923 6381
rect 17865 6341 17877 6375
rect 17911 6372 17923 6375
rect 18322 6372 18328 6384
rect 17911 6344 18328 6372
rect 17911 6341 17923 6344
rect 17865 6335 17923 6341
rect 18322 6332 18328 6344
rect 18380 6332 18386 6384
rect 21192 6372 21220 6412
rect 21342 6409 21354 6412
rect 21388 6440 21400 6443
rect 22186 6440 22192 6452
rect 21388 6412 22192 6440
rect 21388 6409 21400 6412
rect 21342 6403 21400 6409
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 22612 6412 22937 6440
rect 22612 6400 22618 6412
rect 22925 6409 22937 6412
rect 22971 6409 22983 6443
rect 22925 6403 22983 6409
rect 23934 6400 23940 6452
rect 23992 6440 23998 6452
rect 24121 6443 24179 6449
rect 24121 6440 24133 6443
rect 23992 6412 24133 6440
rect 23992 6400 23998 6412
rect 24121 6409 24133 6412
rect 24167 6409 24179 6443
rect 24121 6403 24179 6409
rect 18524 6344 21220 6372
rect 21453 6375 21511 6381
rect 12584 6307 12642 6313
rect 12584 6304 12596 6307
rect 12492 6276 12596 6304
rect 12492 6264 12498 6276
rect 12584 6273 12596 6276
rect 12630 6273 12642 6307
rect 12584 6267 12642 6273
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 12894 6264 12900 6316
rect 12952 6304 12958 6316
rect 12952 6276 12997 6304
rect 12952 6264 12958 6276
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13780 6276 14381 6304
rect 13780 6264 13786 6276
rect 14369 6273 14381 6276
rect 14415 6304 14427 6307
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 14415 6276 15301 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 15289 6273 15301 6276
rect 15335 6304 15347 6307
rect 15654 6304 15660 6316
rect 15335 6276 15660 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16485 6307 16543 6313
rect 16485 6304 16497 6307
rect 16264 6276 16497 6304
rect 16264 6264 16270 6276
rect 16485 6273 16497 6276
rect 16531 6273 16543 6307
rect 18414 6304 18420 6316
rect 18375 6276 18420 6304
rect 16485 6267 16543 6273
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 9068 6239 9126 6245
rect 9068 6236 9080 6239
rect 8864 6208 9080 6236
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6137 1731 6171
rect 2222 6168 2228 6180
rect 2183 6140 2228 6168
rect 1673 6131 1731 6137
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 1688 6100 1716 6131
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 5306 6171 5364 6177
rect 5306 6168 5318 6171
rect 5132 6140 5318 6168
rect 5132 6128 5138 6140
rect 5306 6137 5318 6140
rect 5352 6137 5364 6171
rect 6270 6168 6276 6180
rect 6231 6140 6276 6168
rect 5306 6131 5364 6137
rect 6270 6128 6276 6140
rect 6328 6128 6334 6180
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 7606 6171 7664 6177
rect 7606 6168 7618 6171
rect 7248 6140 7618 6168
rect 7248 6128 7254 6140
rect 7606 6137 7618 6140
rect 7652 6137 7664 6171
rect 7606 6131 7664 6137
rect 1544 6072 1716 6100
rect 1544 6060 1550 6072
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2314 6100 2320 6112
rect 2096 6072 2320 6100
rect 2096 6060 2102 6072
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 2498 6060 2504 6112
rect 2556 6100 2562 6112
rect 2961 6103 3019 6109
rect 2961 6100 2973 6103
rect 2556 6072 2973 6100
rect 2556 6060 2562 6072
rect 2961 6069 2973 6072
rect 3007 6100 3019 6103
rect 3786 6100 3792 6112
rect 3007 6072 3792 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 4396 6072 4445 6100
rect 4396 6060 4402 6072
rect 4433 6069 4445 6072
rect 4479 6069 4491 6103
rect 8202 6100 8208 6112
rect 8163 6072 8208 6100
rect 4433 6063 4491 6069
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 8864 6109 8892 6208
rect 9068 6205 9080 6208
rect 9114 6205 9126 6239
rect 9068 6199 9126 6205
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6205 10471 6239
rect 10962 6236 10968 6248
rect 10923 6208 10968 6236
rect 10413 6199 10471 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14148 6239 14206 6245
rect 14148 6236 14160 6239
rect 13688 6208 14160 6236
rect 13688 6196 13694 6208
rect 14148 6205 14160 6208
rect 14194 6236 14206 6239
rect 18138 6236 18144 6248
rect 14194 6208 14964 6236
rect 18106 6208 18144 6236
rect 14194 6205 14206 6208
rect 14148 6199 14206 6205
rect 12437 6171 12495 6177
rect 12437 6137 12449 6171
rect 12483 6168 12495 6171
rect 12526 6168 12532 6180
rect 12483 6140 12532 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 13504 6140 14013 6168
rect 13504 6128 13510 6140
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14001 6131 14059 6137
rect 14737 6171 14795 6177
rect 14737 6137 14749 6171
rect 14783 6168 14795 6171
rect 14826 6168 14832 6180
rect 14783 6140 14832 6168
rect 14783 6137 14795 6140
rect 14737 6131 14795 6137
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 14936 6112 14964 6208
rect 18138 6196 18144 6208
rect 18196 6245 18202 6248
rect 18196 6239 18254 6245
rect 18196 6205 18208 6239
rect 18242 6236 18254 6239
rect 18524 6236 18552 6344
rect 21453 6341 21465 6375
rect 21499 6372 21511 6375
rect 21634 6372 21640 6384
rect 21499 6344 21640 6372
rect 21499 6341 21511 6344
rect 21453 6335 21511 6341
rect 21634 6332 21640 6344
rect 21692 6372 21698 6384
rect 22281 6375 22339 6381
rect 22281 6372 22293 6375
rect 21692 6344 22293 6372
rect 21692 6332 21698 6344
rect 22281 6341 22293 6344
rect 22327 6372 22339 6375
rect 23474 6372 23480 6384
rect 22327 6344 23480 6372
rect 22327 6341 22339 6344
rect 22281 6335 22339 6341
rect 23474 6332 23480 6344
rect 23532 6332 23538 6384
rect 24854 6372 24860 6384
rect 24815 6344 24860 6372
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 19886 6264 19892 6316
rect 19944 6304 19950 6316
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 19944 6276 20177 6304
rect 19944 6264 19950 6276
rect 20165 6273 20177 6276
rect 20211 6273 20223 6307
rect 21542 6304 21548 6316
rect 21455 6276 21548 6304
rect 20165 6267 20223 6273
rect 21542 6264 21548 6276
rect 21600 6304 21606 6316
rect 22557 6307 22615 6313
rect 22557 6304 22569 6307
rect 21600 6276 22569 6304
rect 21600 6264 21606 6276
rect 22557 6273 22569 6276
rect 22603 6273 22615 6307
rect 22557 6267 22615 6273
rect 18242 6208 18552 6236
rect 18242 6205 18254 6208
rect 18196 6199 18254 6205
rect 18196 6196 18202 6199
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 19518 6236 19524 6248
rect 19300 6208 19524 6236
rect 19300 6196 19306 6208
rect 19518 6196 19524 6208
rect 19576 6236 19582 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19576 6208 19625 6236
rect 19576 6196 19582 6208
rect 19613 6205 19625 6208
rect 19659 6205 19671 6239
rect 20070 6236 20076 6248
rect 20031 6208 20076 6236
rect 19613 6199 19671 6205
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 20714 6196 20720 6248
rect 20772 6236 20778 6248
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 20772 6208 21189 6236
rect 20772 6196 20778 6208
rect 21177 6205 21189 6208
rect 21223 6236 21235 6239
rect 21266 6236 21272 6248
rect 21223 6208 21272 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 24670 6236 24676 6248
rect 24631 6208 24676 6236
rect 24670 6196 24676 6208
rect 24728 6236 24734 6248
rect 25133 6239 25191 6245
rect 25133 6236 25145 6239
rect 24728 6208 25145 6236
rect 24728 6196 24734 6208
rect 25133 6205 25145 6208
rect 25179 6205 25191 6239
rect 25133 6199 25191 6205
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16574 6168 16580 6180
rect 16347 6140 16580 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 17126 6168 17132 6180
rect 17087 6140 17132 6168
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 18046 6168 18052 6180
rect 18007 6140 18052 6168
rect 18046 6128 18052 6140
rect 18104 6128 18110 6180
rect 9214 6109 9220 6112
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8812 6072 8861 6100
rect 8812 6060 8818 6072
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 8849 6063 8907 6069
rect 9171 6103 9220 6109
rect 9171 6069 9183 6103
rect 9217 6069 9220 6103
rect 9171 6063 9220 6069
rect 9214 6060 9220 6063
rect 9272 6060 9278 6112
rect 10686 6100 10692 6112
rect 10647 6072 10692 6100
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 12066 6100 12072 6112
rect 11480 6072 12072 6100
rect 11480 6060 11486 6072
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13722 6100 13728 6112
rect 13683 6072 13728 6100
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 14976 6072 15761 6100
rect 14976 6060 14982 6072
rect 15749 6069 15761 6072
rect 15795 6100 15807 6103
rect 17402 6100 17408 6112
rect 15795 6072 17408 6100
rect 15795 6069 15807 6072
rect 15749 6063 15807 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 17589 6103 17647 6109
rect 17589 6069 17601 6103
rect 17635 6100 17647 6103
rect 17954 6100 17960 6112
rect 17635 6072 17960 6100
rect 17635 6069 17647 6072
rect 17589 6063 17647 6069
rect 17954 6060 17960 6072
rect 18012 6100 18018 6112
rect 18598 6100 18604 6112
rect 18012 6072 18604 6100
rect 18012 6060 18018 6072
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 23658 6100 23664 6112
rect 23619 6072 23664 6100
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 25498 6100 25504 6112
rect 25459 6072 25504 6100
rect 25498 6060 25504 6072
rect 25556 6060 25562 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1544 5868 1593 5896
rect 1544 5856 1550 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 1670 5856 1676 5908
rect 1728 5896 1734 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 1728 5868 2973 5896
rect 1728 5856 1734 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3970 5896 3976 5908
rect 3559 5868 3976 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4120 5868 4261 5896
rect 4120 5856 4126 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4706 5896 4712 5908
rect 4667 5868 4712 5896
rect 4249 5859 4307 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 4816 5868 5825 5896
rect 1210 5788 1216 5840
rect 1268 5828 1274 5840
rect 2133 5831 2191 5837
rect 2133 5828 2145 5831
rect 1268 5800 2145 5828
rect 1268 5788 1274 5800
rect 2133 5797 2145 5800
rect 2179 5828 2191 5831
rect 2682 5828 2688 5840
rect 2179 5800 2688 5828
rect 2179 5797 2191 5800
rect 2133 5791 2191 5797
rect 2682 5788 2688 5800
rect 2740 5828 2746 5840
rect 4816 5828 4844 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 7098 5896 7104 5908
rect 7059 5868 7104 5896
rect 5813 5859 5871 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8018 5856 8024 5908
rect 8076 5856 8082 5908
rect 12526 5896 12532 5908
rect 12487 5868 12532 5896
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 14458 5896 14464 5908
rect 14419 5868 14464 5896
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 14918 5896 14924 5908
rect 14875 5868 14924 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15838 5896 15844 5908
rect 15799 5868 15844 5896
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 16574 5856 16580 5908
rect 16632 5896 16638 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 16632 5868 17049 5896
rect 16632 5856 16638 5868
rect 17037 5865 17049 5868
rect 17083 5896 17095 5899
rect 17862 5896 17868 5908
rect 17083 5868 17868 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18506 5856 18512 5908
rect 18564 5896 18570 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 18564 5868 19625 5896
rect 18564 5856 18570 5868
rect 19613 5865 19625 5868
rect 19659 5896 19671 5899
rect 20070 5896 20076 5908
rect 19659 5868 20076 5896
rect 19659 5865 19671 5868
rect 19613 5859 19671 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 20898 5896 20904 5908
rect 20763 5868 20904 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 22005 5899 22063 5905
rect 22005 5865 22017 5899
rect 22051 5896 22063 5899
rect 22186 5896 22192 5908
rect 22051 5868 22192 5896
rect 22051 5865 22063 5868
rect 22005 5859 22063 5865
rect 22186 5856 22192 5868
rect 22244 5856 22250 5908
rect 22554 5896 22560 5908
rect 22515 5868 22560 5896
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 2740 5800 4844 5828
rect 2740 5788 2746 5800
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 5214 5831 5272 5837
rect 5214 5828 5226 5831
rect 5132 5800 5226 5828
rect 5132 5788 5138 5800
rect 5214 5797 5226 5800
rect 5260 5797 5272 5831
rect 7006 5828 7012 5840
rect 5214 5791 5272 5797
rect 6723 5800 7012 5828
rect 4890 5760 4896 5772
rect 4851 5732 4896 5760
rect 4890 5720 4896 5732
rect 4948 5760 4954 5772
rect 6546 5760 6552 5772
rect 4948 5732 6552 5760
rect 4948 5720 4954 5732
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 6723 5769 6751 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 8036 5828 8064 5856
rect 9858 5828 9864 5840
rect 8036 5800 9352 5828
rect 9819 5800 9864 5828
rect 6708 5763 6766 5769
rect 6708 5729 6720 5763
rect 6754 5729 6766 5763
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 6708 5723 6766 5729
rect 6794 5732 7665 5760
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2222 5692 2228 5704
rect 2087 5664 2228 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2222 5652 2228 5664
rect 2280 5692 2286 5704
rect 2774 5692 2780 5704
rect 2280 5664 2780 5692
rect 2280 5652 2286 5664
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 4338 5652 4344 5704
rect 4396 5692 4402 5704
rect 6794 5692 6822 5732
rect 7653 5729 7665 5732
rect 7699 5760 7711 5763
rect 8018 5760 8024 5772
rect 7699 5732 8024 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 8128 5692 8156 5723
rect 4396 5664 6822 5692
rect 7668 5664 8156 5692
rect 9324 5692 9352 5800
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11241 5831 11299 5837
rect 11241 5828 11253 5831
rect 11204 5800 11253 5828
rect 11204 5788 11210 5800
rect 11241 5797 11253 5800
rect 11287 5828 11299 5831
rect 12066 5828 12072 5840
rect 11287 5800 12072 5828
rect 11287 5797 11299 5800
rect 11241 5791 11299 5797
rect 12066 5788 12072 5800
rect 12124 5828 12130 5840
rect 16482 5837 16488 5840
rect 16479 5828 16488 5837
rect 12124 5800 12848 5828
rect 16443 5800 16488 5828
rect 12124 5788 12130 5800
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9582 5760 9588 5772
rect 9456 5732 9588 5760
rect 9456 5720 9462 5732
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 12434 5760 12440 5772
rect 11440 5732 12440 5760
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9324 5664 9781 5692
rect 4396 5652 4402 5664
rect 7668 5636 7696 5664
rect 2314 5584 2320 5636
rect 2372 5624 2378 5636
rect 2593 5627 2651 5633
rect 2593 5624 2605 5627
rect 2372 5596 2605 5624
rect 2372 5584 2378 5596
rect 2593 5593 2605 5596
rect 2639 5593 2651 5627
rect 2593 5587 2651 5593
rect 7650 5584 7656 5636
rect 7708 5584 7714 5636
rect 6638 5516 6644 5568
rect 6696 5556 6702 5568
rect 6779 5559 6837 5565
rect 6779 5556 6791 5559
rect 6696 5528 6791 5556
rect 6696 5516 6702 5528
rect 6779 5525 6791 5528
rect 6825 5525 6837 5559
rect 7466 5556 7472 5568
rect 7427 5528 7472 5556
rect 6779 5519 6837 5525
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 9600 5556 9628 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 11149 5695 11207 5701
rect 11149 5661 11161 5695
rect 11195 5692 11207 5695
rect 11238 5692 11244 5704
rect 11195 5664 11244 5692
rect 11195 5661 11207 5664
rect 11149 5655 11207 5661
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10060 5624 10088 5655
rect 11238 5652 11244 5664
rect 11296 5692 11302 5704
rect 11440 5701 11468 5732
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 12820 5769 12848 5800
rect 16479 5791 16488 5800
rect 16482 5788 16488 5791
rect 16540 5788 16546 5840
rect 17402 5828 17408 5840
rect 17315 5800 17408 5828
rect 17402 5788 17408 5800
rect 17460 5828 17466 5840
rect 18156 5828 18184 5856
rect 17460 5800 18184 5828
rect 18666 5831 18724 5837
rect 17460 5788 17466 5800
rect 18666 5797 18678 5831
rect 18712 5828 18724 5831
rect 19058 5828 19064 5840
rect 18712 5800 19064 5828
rect 18712 5797 18724 5800
rect 18666 5791 18724 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 12986 5760 12992 5772
rect 12851 5732 12992 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20680 5732 20913 5760
rect 20680 5720 20686 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 21818 5760 21824 5772
rect 21499 5732 21824 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 21818 5720 21824 5732
rect 21876 5760 21882 5772
rect 22094 5760 22100 5772
rect 21876 5732 22100 5760
rect 21876 5720 21882 5732
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 22370 5720 22376 5772
rect 22428 5760 22434 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22428 5732 22477 5760
rect 22428 5720 22434 5732
rect 22465 5729 22477 5732
rect 22511 5729 22523 5763
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22465 5723 22523 5729
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 24026 5760 24032 5772
rect 23987 5732 24032 5760
rect 24026 5720 24032 5732
rect 24084 5720 24090 5772
rect 25130 5760 25136 5772
rect 25091 5732 25136 5760
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 11388 5695 11468 5701
rect 11388 5692 11400 5695
rect 11296 5664 11400 5692
rect 11296 5652 11302 5664
rect 11388 5661 11400 5664
rect 11434 5664 11468 5695
rect 11606 5692 11612 5704
rect 11567 5664 11612 5692
rect 11434 5661 11446 5664
rect 11388 5655 11446 5661
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 12894 5652 12900 5704
rect 12952 5692 12958 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 12952 5664 13185 5692
rect 12952 5652 12958 5664
rect 13173 5661 13185 5664
rect 13219 5692 13231 5695
rect 13722 5692 13728 5704
rect 13219 5664 13728 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13722 5652 13728 5664
rect 13780 5692 13786 5704
rect 14001 5695 14059 5701
rect 14001 5692 14013 5695
rect 13780 5664 14013 5692
rect 13780 5652 13786 5664
rect 14001 5661 14013 5664
rect 14047 5661 14059 5695
rect 14001 5655 14059 5661
rect 16850 5652 16856 5704
rect 16908 5692 16914 5704
rect 17770 5692 17776 5704
rect 16908 5664 17776 5692
rect 16908 5652 16914 5664
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 18414 5692 18420 5704
rect 18371 5664 18420 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 18414 5652 18420 5664
rect 18472 5692 18478 5704
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 18472 5664 21373 5692
rect 18472 5652 18478 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 9732 5596 10088 5624
rect 10781 5627 10839 5633
rect 9732 5584 9738 5596
rect 10781 5593 10793 5627
rect 10827 5624 10839 5627
rect 10962 5624 10968 5636
rect 10827 5596 10968 5624
rect 10827 5593 10839 5596
rect 10781 5587 10839 5593
rect 10962 5584 10968 5596
rect 11020 5624 11026 5636
rect 12802 5624 12808 5636
rect 11020 5596 12808 5624
rect 11020 5584 11026 5596
rect 12802 5584 12808 5596
rect 12860 5624 12866 5636
rect 13265 5627 13323 5633
rect 13265 5624 13277 5627
rect 12860 5596 13277 5624
rect 12860 5584 12866 5596
rect 13265 5593 13277 5596
rect 13311 5593 13323 5627
rect 25314 5624 25320 5636
rect 25275 5596 25320 5624
rect 13265 5587 13323 5593
rect 25314 5584 25320 5596
rect 25372 5584 25378 5636
rect 10134 5556 10140 5568
rect 9600 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 11514 5556 11520 5568
rect 11475 5528 11520 5556
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11698 5556 11704 5568
rect 11659 5528 11704 5556
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 12943 5559 13001 5565
rect 12943 5556 12955 5559
rect 12492 5528 12955 5556
rect 12492 5516 12498 5528
rect 12943 5525 12955 5528
rect 12989 5525 13001 5559
rect 12943 5519 13001 5525
rect 13081 5559 13139 5565
rect 13081 5525 13093 5559
rect 13127 5556 13139 5559
rect 13446 5556 13452 5568
rect 13127 5528 13452 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13446 5516 13452 5528
rect 13504 5556 13510 5568
rect 14458 5556 14464 5568
rect 13504 5528 14464 5556
rect 13504 5516 13510 5528
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 19242 5556 19248 5568
rect 19203 5528 19248 5556
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19978 5556 19984 5568
rect 19939 5528 19984 5556
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 24210 5556 24216 5568
rect 24171 5528 24216 5556
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 2777 5355 2835 5361
rect 2777 5352 2789 5355
rect 2740 5324 2789 5352
rect 2740 5312 2746 5324
rect 2777 5321 2789 5324
rect 2823 5321 2835 5355
rect 2777 5315 2835 5321
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5074 5352 5080 5364
rect 5031 5324 5080 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7248 5324 7389 5352
rect 7248 5312 7254 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 7392 5284 7420 5315
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 8076 5324 8769 5352
rect 8076 5312 8082 5324
rect 8757 5321 8769 5324
rect 8803 5321 8815 5355
rect 8757 5315 8815 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9398 5352 9404 5364
rect 8987 5324 9404 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 8772 5284 8800 5315
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 11011 5355 11069 5361
rect 11011 5352 11023 5355
rect 10284 5324 11023 5352
rect 10284 5312 10290 5324
rect 11011 5321 11023 5324
rect 11057 5321 11069 5355
rect 11011 5315 11069 5321
rect 11425 5355 11483 5361
rect 11425 5321 11437 5355
rect 11471 5352 11483 5355
rect 11606 5352 11612 5364
rect 11471 5324 11612 5352
rect 11471 5321 11483 5324
rect 11425 5315 11483 5321
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14792 5324 15025 5352
rect 14792 5312 14798 5324
rect 15013 5321 15025 5324
rect 15059 5321 15071 5355
rect 15013 5315 15071 5321
rect 15473 5355 15531 5361
rect 15473 5321 15485 5355
rect 15519 5352 15531 5355
rect 16114 5352 16120 5364
rect 15519 5324 16120 5352
rect 15519 5321 15531 5324
rect 15473 5315 15531 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 16482 5352 16488 5364
rect 16255 5324 16488 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 18601 5355 18659 5361
rect 18601 5321 18613 5355
rect 18647 5352 18659 5355
rect 19058 5352 19064 5364
rect 18647 5324 19064 5352
rect 18647 5321 18659 5324
rect 18601 5315 18659 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19518 5312 19524 5364
rect 19576 5352 19582 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 19576 5324 20453 5352
rect 19576 5312 19582 5324
rect 20441 5321 20453 5324
rect 20487 5352 20499 5355
rect 20622 5352 20628 5364
rect 20487 5324 20628 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22152 5324 22477 5352
rect 22152 5312 22158 5324
rect 22465 5321 22477 5324
rect 22511 5352 22523 5355
rect 22922 5352 22928 5364
rect 22511 5324 22928 5352
rect 22511 5321 22523 5324
rect 22465 5315 22523 5321
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 24026 5312 24032 5364
rect 24084 5352 24090 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 24084 5324 24685 5352
rect 24084 5312 24090 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 25130 5352 25136 5364
rect 25091 5324 25136 5352
rect 24673 5315 24731 5321
rect 25130 5312 25136 5324
rect 25188 5312 25194 5364
rect 11146 5284 11152 5296
rect 7392 5256 7788 5284
rect 8772 5256 11152 5284
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3694 5216 3700 5228
rect 3559 5188 3700 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3694 5176 3700 5188
rect 3752 5216 3758 5228
rect 5905 5219 5963 5225
rect 3752 5188 5488 5216
rect 3752 5176 3758 5188
rect 3896 5157 3924 5188
rect 5460 5157 5488 5188
rect 5905 5185 5917 5219
rect 5951 5216 5963 5219
rect 7466 5216 7472 5228
rect 5951 5188 7472 5216
rect 5951 5185 5963 5188
rect 5905 5179 5963 5185
rect 7466 5176 7472 5188
rect 7524 5216 7530 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 7524 5188 7573 5216
rect 7524 5176 7530 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5117 4215 5151
rect 4157 5111 4215 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5534 5148 5540 5160
rect 5491 5120 5540 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 1946 5040 1952 5092
rect 2004 5080 2010 5092
rect 2004 5052 2049 5080
rect 2004 5040 2010 5052
rect 3694 5040 3700 5092
rect 3752 5080 3758 5092
rect 4172 5080 4200 5111
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 5767 5120 6316 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 5258 5080 5264 5092
rect 3752 5052 5264 5080
rect 3752 5040 3758 5052
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 6288 5089 6316 5120
rect 6273 5083 6331 5089
rect 6273 5049 6285 5083
rect 6319 5080 6331 5083
rect 7650 5080 7656 5092
rect 6319 5052 7656 5080
rect 6319 5049 6331 5052
rect 6273 5043 6331 5049
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 7760 5080 7788 5256
rect 11146 5244 11152 5256
rect 11204 5284 11210 5296
rect 13170 5284 13176 5296
rect 11204 5256 13176 5284
rect 11204 5244 11210 5256
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8772 5188 9137 5216
rect 8772 5160 8800 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9674 5216 9680 5228
rect 9635 5188 9680 5216
rect 9125 5179 9183 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11238 5216 11244 5228
rect 10827 5188 11244 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 8754 5108 8760 5160
rect 8812 5108 8818 5160
rect 10940 5151 10998 5157
rect 10940 5117 10952 5151
rect 10986 5148 10998 5151
rect 11054 5148 11060 5160
rect 10986 5120 11060 5148
rect 10986 5117 10998 5120
rect 10940 5111 10998 5117
rect 11054 5108 11060 5120
rect 11112 5148 11118 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11112 5120 11713 5148
rect 11112 5108 11118 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 12360 5148 12388 5256
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 18874 5284 18880 5296
rect 18835 5256 18880 5284
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 20073 5287 20131 5293
rect 20073 5253 20085 5287
rect 20119 5284 20131 5287
rect 20119 5256 21772 5284
rect 20119 5253 20131 5256
rect 20073 5247 20131 5253
rect 16022 5176 16028 5228
rect 16080 5216 16086 5228
rect 16485 5219 16543 5225
rect 16485 5216 16497 5219
rect 16080 5188 16497 5216
rect 16080 5176 16086 5188
rect 16485 5185 16497 5188
rect 16531 5216 16543 5219
rect 16758 5216 16764 5228
rect 16531 5188 16764 5216
rect 16531 5185 16543 5188
rect 16485 5179 16543 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 17126 5176 17132 5188
rect 17184 5216 17190 5228
rect 19521 5219 19579 5225
rect 19521 5216 19533 5219
rect 17184 5188 19533 5216
rect 17184 5176 17190 5188
rect 19521 5185 19533 5188
rect 19567 5216 19579 5219
rect 19978 5216 19984 5228
rect 19567 5188 19984 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 21082 5216 21088 5228
rect 21043 5188 21088 5216
rect 21082 5176 21088 5188
rect 21140 5176 21146 5228
rect 21744 5225 21772 5256
rect 22370 5244 22376 5296
rect 22428 5284 22434 5296
rect 23017 5287 23075 5293
rect 23017 5284 23029 5287
rect 22428 5256 23029 5284
rect 22428 5244 22434 5256
rect 23017 5253 23029 5256
rect 23063 5253 23075 5287
rect 23017 5247 23075 5253
rect 25409 5287 25467 5293
rect 25409 5253 25421 5287
rect 25455 5284 25467 5287
rect 26694 5284 26700 5296
rect 25455 5256 26700 5284
rect 25455 5253 25467 5256
rect 25409 5247 25467 5253
rect 26694 5244 26700 5256
rect 26752 5244 26758 5296
rect 21729 5219 21787 5225
rect 21729 5185 21741 5219
rect 21775 5216 21787 5219
rect 21910 5216 21916 5228
rect 21775 5188 21916 5216
rect 21775 5185 21787 5188
rect 21729 5179 21787 5185
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12360 5120 12449 5148
rect 11701 5111 11759 5117
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12860 5120 12909 5148
rect 12860 5108 12866 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 14182 5148 14188 5160
rect 14143 5120 14188 5148
rect 12897 5111 12955 5117
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 14826 5148 14832 5160
rect 14599 5120 14832 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 7882 5083 7940 5089
rect 7882 5080 7894 5083
rect 7760 5052 7894 5080
rect 7882 5049 7894 5052
rect 7928 5049 7940 5083
rect 7882 5043 7940 5049
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 9401 5083 9459 5089
rect 9401 5080 9413 5083
rect 8352 5052 9413 5080
rect 8352 5040 8358 5052
rect 1673 5015 1731 5021
rect 1673 4981 1685 5015
rect 1719 5012 1731 5015
rect 1964 5012 1992 5040
rect 9324 5024 9352 5052
rect 9401 5049 9413 5052
rect 9447 5049 9459 5083
rect 9401 5043 9459 5049
rect 9493 5083 9551 5089
rect 9493 5049 9505 5083
rect 9539 5080 9551 5083
rect 9582 5080 9588 5092
rect 9539 5052 9588 5080
rect 9539 5049 9551 5052
rect 9493 5043 9551 5049
rect 9582 5040 9588 5052
rect 9640 5040 9646 5092
rect 9858 5040 9864 5092
rect 9916 5080 9922 5092
rect 10413 5083 10471 5089
rect 10413 5080 10425 5083
rect 9916 5052 10425 5080
rect 9916 5040 9922 5052
rect 10413 5049 10425 5052
rect 10459 5080 10471 5083
rect 10778 5080 10784 5092
rect 10459 5052 10784 5080
rect 10459 5049 10471 5052
rect 10413 5043 10471 5049
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 13170 5080 13176 5092
rect 13131 5052 13176 5080
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 13909 5083 13967 5089
rect 13909 5049 13921 5083
rect 13955 5080 13967 5083
rect 14568 5080 14596 5111
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 23753 5151 23811 5157
rect 23753 5117 23765 5151
rect 23799 5117 23811 5151
rect 23753 5111 23811 5117
rect 14734 5080 14740 5092
rect 13955 5052 14596 5080
rect 14695 5052 14740 5080
rect 13955 5049 13967 5052
rect 13909 5043 13967 5049
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 15841 5083 15899 5089
rect 15841 5049 15853 5083
rect 15887 5080 15899 5083
rect 16574 5080 16580 5092
rect 15887 5052 16580 5080
rect 15887 5049 15899 5052
rect 15841 5043 15899 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 19242 5040 19248 5092
rect 19300 5080 19306 5092
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 19300 5052 19349 5080
rect 19300 5040 19306 5052
rect 19337 5049 19349 5052
rect 19383 5080 19395 5083
rect 19613 5083 19671 5089
rect 19613 5080 19625 5083
rect 19383 5052 19625 5080
rect 19383 5049 19395 5052
rect 19337 5043 19395 5049
rect 19613 5049 19625 5052
rect 19659 5080 19671 5083
rect 19978 5080 19984 5092
rect 19659 5052 19984 5080
rect 19659 5049 19671 5052
rect 19613 5043 19671 5049
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 21177 5083 21235 5089
rect 21177 5049 21189 5083
rect 21223 5049 21235 5083
rect 23658 5080 23664 5092
rect 23619 5052 23664 5080
rect 21177 5043 21235 5049
rect 3878 5012 3884 5024
rect 1719 4984 1992 5012
rect 3839 4984 3884 5012
rect 1719 4981 1731 4984
rect 1673 4975 1731 4981
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 8481 5015 8539 5021
rect 8481 4981 8493 5015
rect 8527 5012 8539 5015
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8527 4984 8953 5012
rect 8527 4981 8539 4984
rect 8481 4975 8539 4981
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 8941 4975 8999 4981
rect 9306 4972 9312 5024
rect 9364 4972 9370 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12894 5012 12900 5024
rect 12032 4984 12900 5012
rect 12032 4972 12038 4984
rect 12894 4972 12900 4984
rect 12952 5012 12958 5024
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 12952 4984 13461 5012
rect 12952 4972 12958 4984
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 13449 4975 13507 4981
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 20898 5012 20904 5024
rect 20859 4984 20904 5012
rect 20898 4972 20904 4984
rect 20956 5012 20962 5024
rect 21192 5012 21220 5043
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 20956 4984 21220 5012
rect 20956 4972 20962 4984
rect 21910 4972 21916 5024
rect 21968 5012 21974 5024
rect 22557 5015 22615 5021
rect 22557 5012 22569 5015
rect 21968 4984 22569 5012
rect 21968 4972 21974 4984
rect 22557 4981 22569 4984
rect 22603 4981 22615 5015
rect 22557 4975 22615 4981
rect 23477 5015 23535 5021
rect 23477 4981 23489 5015
rect 23523 5012 23535 5015
rect 23768 5012 23796 5111
rect 24118 5108 24124 5160
rect 24176 5148 24182 5160
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 24176 5120 25237 5148
rect 24176 5108 24182 5120
rect 25225 5117 25237 5120
rect 25271 5148 25283 5151
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25271 5120 25789 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 23842 5012 23848 5024
rect 23523 4984 23848 5012
rect 23523 4981 23535 4984
rect 23477 4975 23535 4981
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2832 4780 3249 4808
rect 2832 4768 2838 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3694 4808 3700 4820
rect 3655 4780 3700 4808
rect 3237 4771 3295 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 4706 4808 4712 4820
rect 4667 4780 4712 4808
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5592 4780 5641 4808
rect 5592 4768 5598 4780
rect 5629 4777 5641 4780
rect 5675 4777 5687 4811
rect 9306 4808 9312 4820
rect 9267 4780 9312 4808
rect 5629 4771 5687 4777
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10134 4808 10140 4820
rect 9999 4780 10140 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11514 4808 11520 4820
rect 11379 4780 11520 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13446 4808 13452 4820
rect 12943 4780 13452 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 2406 4740 2412 4752
rect 2367 4712 2412 4740
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6365 4743 6423 4749
rect 6365 4740 6377 4743
rect 6328 4712 6377 4740
rect 6328 4700 6334 4712
rect 6365 4709 6377 4712
rect 6411 4740 6423 4743
rect 6730 4740 6736 4752
rect 6411 4712 6736 4740
rect 6411 4709 6423 4712
rect 6365 4703 6423 4709
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 7926 4740 7932 4752
rect 7887 4712 7932 4740
rect 7926 4700 7932 4712
rect 7984 4700 7990 4752
rect 10407 4743 10465 4749
rect 10407 4709 10419 4743
rect 10453 4740 10465 4743
rect 10778 4740 10784 4752
rect 10453 4712 10784 4740
rect 10453 4709 10465 4712
rect 10407 4703 10465 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 11146 4700 11152 4752
rect 11204 4740 11210 4752
rect 11609 4743 11667 4749
rect 11609 4740 11621 4743
rect 11204 4712 11621 4740
rect 11204 4700 11210 4712
rect 11609 4709 11621 4712
rect 11655 4709 11667 4743
rect 11609 4703 11667 4709
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 12912 4740 12940 4771
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 14240 4780 14381 4808
rect 14240 4768 14246 4780
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 16390 4808 16396 4820
rect 16351 4780 16396 4808
rect 14369 4771 14427 4777
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 16758 4808 16764 4820
rect 16719 4780 16764 4808
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 18414 4808 18420 4820
rect 18375 4780 18420 4808
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 19797 4811 19855 4817
rect 19797 4777 19809 4811
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 20990 4808 20996 4820
rect 20763 4780 20996 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 12124 4712 12940 4740
rect 17129 4743 17187 4749
rect 12124 4700 12130 4712
rect 17129 4709 17141 4743
rect 17175 4740 17187 4743
rect 17494 4740 17500 4752
rect 17175 4712 17500 4740
rect 17175 4709 17187 4712
rect 17129 4703 17187 4709
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 19058 4700 19064 4752
rect 19116 4740 19122 4752
rect 19198 4743 19256 4749
rect 19198 4740 19210 4743
rect 19116 4712 19210 4740
rect 19116 4700 19122 4712
rect 19198 4709 19210 4712
rect 19244 4709 19256 4743
rect 19812 4740 19840 4771
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 19812 4712 21097 4740
rect 19198 4703 19256 4709
rect 21085 4709 21097 4712
rect 21131 4740 21143 4743
rect 21634 4740 21640 4752
rect 21131 4712 21640 4740
rect 21131 4709 21143 4712
rect 21085 4703 21143 4709
rect 21634 4700 21640 4712
rect 21692 4740 21698 4752
rect 21692 4712 22692 4740
rect 21692 4700 21698 4712
rect 4338 4632 4344 4684
rect 4396 4672 4402 4684
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 4396 4644 4629 4672
rect 4396 4632 4402 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 5258 4672 5264 4684
rect 5215 4644 5264 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10134 4672 10140 4684
rect 10091 4644 10140 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10134 4632 10140 4644
rect 10192 4672 10198 4684
rect 10686 4672 10692 4684
rect 10192 4644 10692 4672
rect 10192 4632 10198 4644
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 11790 4672 11796 4684
rect 11751 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 13998 4672 14004 4684
rect 13959 4644 14004 4672
rect 13998 4632 14004 4644
rect 14056 4672 14062 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 14056 4644 15301 4672
rect 14056 4632 14062 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15838 4672 15844 4684
rect 15799 4644 15844 4672
rect 15289 4635 15347 4641
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 18874 4672 18880 4684
rect 18835 4644 18880 4672
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 22664 4681 22692 4712
rect 22649 4675 22707 4681
rect 22649 4641 22661 4675
rect 22695 4641 22707 4675
rect 24670 4672 24676 4684
rect 24631 4644 24676 4672
rect 22649 4635 22707 4641
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2498 4604 2504 4616
rect 2363 4576 2504 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3050 4604 3056 4616
rect 3007 4576 3056 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4604 6331 4607
rect 6362 4604 6368 4616
rect 6319 4576 6368 4604
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6963 4576 7297 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7285 4573 7297 4576
rect 7331 4604 7343 4607
rect 7834 4604 7840 4616
rect 7331 4576 7840 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8754 4604 8760 4616
rect 8527 4576 8760 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 11974 4564 11980 4616
rect 12032 4604 12038 4616
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 12032 4576 12173 4604
rect 12032 4564 12038 4576
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 12584 4576 13369 4604
rect 12584 4564 12590 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 17034 4604 17040 4616
rect 16995 4576 17040 4604
rect 13357 4567 13415 4573
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17276 4576 17325 4604
rect 17276 4564 17282 4576
rect 17313 4573 17325 4576
rect 17359 4604 17371 4607
rect 17678 4604 17684 4616
rect 17359 4576 17684 4604
rect 17359 4573 17371 4576
rect 17313 4567 17371 4573
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 20864 4576 21005 4604
rect 20864 4564 20870 4576
rect 20993 4573 21005 4576
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 21637 4607 21695 4613
rect 21637 4573 21649 4607
rect 21683 4604 21695 4607
rect 21726 4604 21732 4616
rect 21683 4576 21732 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 21726 4564 21732 4576
rect 21784 4564 21790 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22465 4607 22523 4613
rect 22465 4604 22477 4607
rect 22244 4576 22477 4604
rect 22244 4564 22250 4576
rect 22465 4573 22477 4576
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 10686 4536 10692 4548
rect 10100 4508 10692 4536
rect 10100 4496 10106 4508
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 10962 4536 10968 4548
rect 10923 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 15378 4536 15384 4548
rect 15339 4508 15384 4536
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 7650 4468 7656 4480
rect 7611 4440 7656 4468
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 11882 4468 11888 4480
rect 11296 4440 11888 4468
rect 11296 4428 11302 4440
rect 11882 4428 11888 4440
rect 11940 4477 11946 4480
rect 11940 4471 11989 4477
rect 11940 4437 11943 4471
rect 11977 4437 11989 4471
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 11940 4431 11989 4437
rect 11940 4428 11946 4431
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12492 4440 12537 4468
rect 12492 4428 12498 4440
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 13044 4440 13185 4468
rect 13044 4428 13050 4440
rect 13173 4437 13185 4440
rect 13219 4437 13231 4471
rect 14826 4468 14832 4480
rect 14787 4440 14832 4468
rect 13173 4431 13231 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 24118 4428 24124 4480
rect 24176 4468 24182 4480
rect 24305 4471 24363 4477
rect 24305 4468 24317 4471
rect 24176 4440 24317 4468
rect 24176 4428 24182 4440
rect 24305 4437 24317 4440
rect 24351 4437 24363 4471
rect 24305 4431 24363 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2406 4264 2412 4276
rect 2271 4236 2412 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 3878 4264 3884 4276
rect 3839 4236 3884 4264
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4338 4264 4344 4276
rect 4299 4236 4344 4264
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4709 4267 4767 4273
rect 4709 4233 4721 4267
rect 4755 4264 4767 4267
rect 5074 4264 5080 4276
rect 4755 4236 5080 4264
rect 4755 4233 4767 4236
rect 4709 4227 4767 4233
rect 5074 4224 5080 4236
rect 5132 4224 5138 4276
rect 6270 4264 6276 4276
rect 6231 4236 6276 4264
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6420 4236 6561 4264
rect 6420 4224 6426 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7248 4236 7573 4264
rect 7248 4224 7254 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 7561 4227 7619 4233
rect 10965 4267 11023 4273
rect 10965 4233 10977 4267
rect 11011 4264 11023 4267
rect 12066 4264 12072 4276
rect 11011 4236 12072 4264
rect 11011 4233 11023 4236
rect 10965 4227 11023 4233
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2590 4128 2596 4140
rect 2455 4100 2596 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3896 4128 3924 4224
rect 7576 4196 7604 4227
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 19058 4264 19064 4276
rect 19019 4236 19064 4264
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 21634 4264 21640 4276
rect 21595 4236 21640 4264
rect 21634 4224 21640 4236
rect 21692 4264 21698 4276
rect 22741 4267 22799 4273
rect 22741 4264 22753 4267
rect 21692 4236 22753 4264
rect 21692 4224 21698 4236
rect 22741 4233 22753 4236
rect 22787 4233 22799 4267
rect 22741 4227 22799 4233
rect 7576 4168 7880 4196
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 3896 4100 4813 4128
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7742 4128 7748 4140
rect 7331 4100 7748 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 1872 3964 2513 3992
rect 1872 3936 1900 3964
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 2590 3952 2596 4004
rect 2648 3992 2654 4004
rect 3329 3995 3387 4001
rect 3329 3992 3341 3995
rect 2648 3964 3341 3992
rect 2648 3952 2654 3964
rect 3329 3961 3341 3964
rect 3375 3961 3387 3995
rect 3329 3955 3387 3961
rect 5074 3952 5080 4004
rect 5132 4001 5138 4004
rect 5132 3995 5180 4001
rect 5132 3961 5134 3995
rect 5168 3961 5180 3995
rect 7852 3992 7880 4168
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 14884 4168 15148 4196
rect 14884 4156 14890 4168
rect 9030 4128 9036 4140
rect 8991 4100 9036 4128
rect 9030 4088 9036 4100
rect 9088 4128 9094 4140
rect 9585 4131 9643 4137
rect 9585 4128 9597 4131
rect 9088 4100 9597 4128
rect 9088 4088 9094 4100
rect 9585 4097 9597 4100
rect 9631 4097 9643 4131
rect 9858 4128 9864 4140
rect 9819 4100 9864 4128
rect 9585 4091 9643 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 12710 4128 12716 4140
rect 12623 4100 12716 4128
rect 12710 4088 12716 4100
rect 12768 4128 12774 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 12768 4100 14013 4128
rect 12768 4088 12774 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 15120 4128 15148 4168
rect 16390 4156 16396 4208
rect 16448 4196 16454 4208
rect 16448 4168 16528 4196
rect 16448 4156 16454 4168
rect 16500 4128 16528 4168
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 18932 4168 19288 4196
rect 18932 4156 18938 4168
rect 19260 4128 19288 4168
rect 19978 4156 19984 4208
rect 20036 4196 20042 4208
rect 20036 4168 20668 4196
rect 20036 4156 20042 4168
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 15120 4100 15332 4128
rect 16500 4100 16896 4128
rect 19260 4100 19441 4128
rect 14001 4091 14059 4097
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 10778 4060 10784 4072
rect 10643 4032 10784 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11146 4069 11152 4072
rect 11124 4063 11152 4069
rect 11124 4029 11136 4063
rect 11204 4060 11210 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11204 4032 11529 4060
rect 11124 4023 11152 4029
rect 11146 4020 11152 4023
rect 11204 4020 11210 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 14918 4060 14924 4072
rect 14700 4032 14924 4060
rect 14700 4020 14706 4032
rect 14918 4020 14924 4032
rect 14976 4060 14982 4072
rect 15304 4069 15332 4100
rect 16868 4069 16896 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 20070 4128 20076 4140
rect 20031 4100 20076 4128
rect 19429 4091 19487 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20640 4128 20668 4168
rect 20990 4128 20996 4140
rect 20640 4100 20996 4128
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 21361 4131 21419 4137
rect 21361 4097 21373 4131
rect 21407 4128 21419 4131
rect 21726 4128 21732 4140
rect 21407 4100 21732 4128
rect 21407 4097 21419 4100
rect 21361 4091 21419 4097
rect 21726 4088 21732 4100
rect 21784 4088 21790 4140
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22152 4100 22232 4128
rect 22152 4088 22158 4100
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14976 4032 15117 4060
rect 14976 4020 14982 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4029 15347 4063
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 15289 4023 15347 4029
rect 15488 4032 16221 4060
rect 8066 3995 8124 4001
rect 8066 3992 8078 3995
rect 7852 3964 8078 3992
rect 5132 3955 5180 3961
rect 8066 3961 8078 3964
rect 8112 3961 8124 3995
rect 9398 3992 9404 4004
rect 9311 3964 9404 3992
rect 8066 3955 8124 3961
rect 5132 3952 5138 3955
rect 9398 3952 9404 3964
rect 9456 3992 9462 4004
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 9456 3964 9689 3992
rect 9456 3952 9462 3964
rect 9677 3961 9689 3964
rect 9723 3961 9735 3995
rect 9677 3955 9735 3961
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12299 3964 12817 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12805 3961 12817 3964
rect 12851 3992 12863 3995
rect 13170 3992 13176 4004
rect 12851 3964 13176 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 13357 3995 13415 4001
rect 13357 3961 13369 3995
rect 13403 3992 13415 3995
rect 13446 3992 13452 4004
rect 13403 3964 13452 3992
rect 13403 3961 13415 3964
rect 13357 3955 13415 3961
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 15120 3992 15148 4023
rect 15488 3992 15516 4032
rect 16209 4029 16221 4032
rect 16255 4060 16267 4063
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 16255 4032 16405 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 16853 4063 16911 4069
rect 16853 4029 16865 4063
rect 16899 4029 16911 4063
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 16853 4023 16911 4029
rect 17052 4032 17785 4060
rect 15120 3964 15516 3992
rect 15565 3995 15623 4001
rect 15565 3961 15577 3995
rect 15611 3992 15623 3995
rect 15746 3992 15752 4004
rect 15611 3964 15752 3992
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 15746 3952 15752 3964
rect 15804 3952 15810 4004
rect 16408 3992 16436 4023
rect 17052 3992 17080 4032
rect 17773 4029 17785 4032
rect 17819 4060 17831 4063
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17819 4032 18061 4060
rect 17819 4029 17831 4032
rect 17773 4023 17831 4029
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 22204 4069 22232 4100
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18380 4032 18521 4060
rect 18380 4020 18386 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 22189 4063 22247 4069
rect 22189 4029 22201 4063
rect 22235 4029 22247 4063
rect 23753 4063 23811 4069
rect 23753 4060 23765 4063
rect 22189 4023 22247 4029
rect 23492 4032 23765 4060
rect 16408 3964 17080 3992
rect 17129 3995 17187 4001
rect 17129 3961 17141 3995
rect 17175 3992 17187 3995
rect 17678 3992 17684 4004
rect 17175 3964 17684 3992
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 20714 3992 20720 4004
rect 20675 3964 20720 3992
rect 20714 3952 20720 3964
rect 20772 3952 20778 4004
rect 20809 3995 20867 4001
rect 20809 3961 20821 3995
rect 20855 3961 20867 3995
rect 22002 3992 22008 4004
rect 20809 3955 20867 3961
rect 21468 3964 22008 3992
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 8662 3924 8668 3936
rect 8623 3896 8668 3924
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 11195 3927 11253 3933
rect 11195 3893 11207 3927
rect 11241 3924 11253 3927
rect 11330 3924 11336 3936
rect 11241 3896 11336 3924
rect 11241 3893 11253 3896
rect 11195 3887 11253 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 13725 3927 13783 3933
rect 13725 3893 13737 3927
rect 13771 3924 13783 3927
rect 13998 3924 14004 3936
rect 13771 3896 14004 3924
rect 13771 3893 13783 3896
rect 13725 3887 13783 3893
rect 13998 3884 14004 3896
rect 14056 3924 14062 3936
rect 14737 3927 14795 3933
rect 14737 3924 14749 3927
rect 14056 3896 14749 3924
rect 14056 3884 14062 3896
rect 14737 3893 14749 3896
rect 14783 3924 14795 3927
rect 14826 3924 14832 3936
rect 14783 3896 14832 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 17494 3924 17500 3936
rect 17455 3896 17500 3924
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 18138 3924 18144 3936
rect 18099 3896 18144 3924
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3924 19671 3927
rect 19978 3924 19984 3936
rect 19659 3896 19984 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20533 3927 20591 3933
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 20824 3924 20852 3955
rect 21468 3924 21496 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 23492 3936 23520 4032
rect 23753 4029 23765 4032
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 23934 4020 23940 4072
rect 23992 4020 23998 4072
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 25225 4063 25283 4069
rect 25225 4060 25237 4063
rect 24820 4032 25237 4060
rect 24820 4020 24826 4032
rect 25225 4029 25237 4032
rect 25271 4060 25283 4063
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 25271 4032 25789 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 23658 3952 23664 4004
rect 23716 3992 23722 4004
rect 23952 3992 23980 4020
rect 23716 3964 23980 3992
rect 23716 3952 23722 3964
rect 20579 3896 21496 3924
rect 22373 3927 22431 3933
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 22373 3893 22385 3927
rect 22419 3924 22431 3927
rect 22646 3924 22652 3936
rect 22419 3896 22652 3924
rect 22419 3893 22431 3896
rect 22373 3887 22431 3893
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 23474 3924 23480 3936
rect 23435 3896 23480 3924
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24670 3924 24676 3936
rect 24631 3896 24676 3924
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 25130 3884 25136 3936
rect 25188 3924 25194 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 25188 3896 25421 3924
rect 25188 3884 25194 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2406 3720 2412 3732
rect 2363 3692 2412 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3720 4767 3723
rect 5258 3720 5264 3732
rect 4755 3692 5264 3720
rect 4755 3689 4767 3692
rect 4709 3683 4767 3689
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 6086 3720 6092 3732
rect 6047 3692 6092 3720
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 8110 3720 8116 3732
rect 7616 3692 8116 3720
rect 7616 3680 7622 3692
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 10134 3720 10140 3732
rect 8904 3692 9996 3720
rect 10095 3692 10140 3720
rect 8904 3680 8910 3692
rect 1949 3655 2007 3661
rect 1949 3621 1961 3655
rect 1995 3652 2007 3655
rect 2498 3652 2504 3664
rect 1995 3624 2504 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 2498 3612 2504 3624
rect 2556 3612 2562 3664
rect 2593 3655 2651 3661
rect 2593 3621 2605 3655
rect 2639 3652 2651 3655
rect 3234 3652 3240 3664
rect 2639 3624 3240 3652
rect 2639 3621 2651 3624
rect 2593 3615 2651 3621
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 5074 3612 5080 3664
rect 5132 3661 5138 3664
rect 5132 3655 5180 3661
rect 5132 3621 5134 3655
rect 5168 3621 5180 3655
rect 5132 3615 5180 3621
rect 6457 3655 6515 3661
rect 6457 3621 6469 3655
rect 6503 3652 6515 3655
rect 6638 3652 6644 3664
rect 6503 3624 6644 3652
rect 6503 3621 6515 3624
rect 6457 3615 6515 3621
rect 5132 3612 5138 3615
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 9815 3655 9873 3661
rect 9815 3652 9827 3655
rect 6788 3624 6833 3652
rect 8128 3624 9827 3652
rect 6788 3612 6794 3624
rect 8128 3596 8156 3624
rect 9815 3621 9827 3624
rect 9861 3621 9873 3655
rect 9968 3652 9996 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11974 3720 11980 3732
rect 10836 3692 11165 3720
rect 11935 3692 11980 3720
rect 10836 3680 10842 3692
rect 10502 3652 10508 3664
rect 9968 3624 10508 3652
rect 9815 3615 9873 3621
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 11137 3661 11165 3692
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 12618 3720 12624 3732
rect 12483 3692 12624 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 12802 3720 12808 3732
rect 12763 3692 12808 3720
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13265 3723 13323 3729
rect 13265 3689 13277 3723
rect 13311 3720 13323 3723
rect 13538 3720 13544 3732
rect 13311 3692 13544 3720
rect 13311 3689 13323 3692
rect 13265 3683 13323 3689
rect 11122 3655 11180 3661
rect 11122 3621 11134 3655
rect 11168 3652 11180 3655
rect 11514 3652 11520 3664
rect 11168 3624 11520 3652
rect 11168 3621 11180 3624
rect 11122 3615 11180 3621
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 1464 3587 1522 3593
rect 1464 3553 1476 3587
rect 1510 3584 1522 3587
rect 2314 3584 2320 3596
rect 1510 3556 2320 3584
rect 1510 3553 1522 3556
rect 1464 3547 1522 3553
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 4801 3587 4859 3593
rect 4801 3584 4813 3587
rect 4764 3556 4813 3584
rect 4764 3544 4770 3556
rect 4801 3553 4813 3556
rect 4847 3553 4859 3587
rect 8110 3584 8116 3596
rect 8023 3556 8116 3584
rect 4801 3547 4859 3553
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 9712 3587 9770 3593
rect 9712 3584 9724 3587
rect 8812 3556 9724 3584
rect 8812 3544 8818 3556
rect 9712 3553 9724 3556
rect 9758 3553 9770 3587
rect 9712 3547 9770 3553
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 10870 3584 10876 3596
rect 10827 3556 10876 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 13372 3593 13400 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 13872 3692 14289 3720
rect 13872 3680 13878 3692
rect 14277 3689 14289 3692
rect 14323 3720 14335 3723
rect 15378 3720 15384 3732
rect 14323 3692 15384 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 17034 3720 17040 3732
rect 16995 3692 17040 3720
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 17678 3720 17684 3732
rect 17639 3692 17684 3720
rect 17678 3680 17684 3692
rect 17736 3720 17742 3732
rect 19337 3723 19395 3729
rect 17736 3692 18460 3720
rect 17736 3680 17742 3692
rect 13719 3655 13777 3661
rect 13719 3621 13731 3655
rect 13765 3652 13777 3655
rect 14918 3652 14924 3664
rect 13765 3624 13860 3652
rect 14879 3624 14924 3652
rect 13765 3621 13777 3624
rect 13719 3615 13777 3621
rect 13832 3596 13860 3624
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 16090 3655 16148 3661
rect 16090 3621 16102 3655
rect 16136 3652 16148 3655
rect 16482 3652 16488 3664
rect 16136 3624 16488 3652
rect 16136 3621 16148 3624
rect 16090 3615 16148 3621
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 18141 3655 18199 3661
rect 18141 3621 18153 3655
rect 18187 3652 18199 3655
rect 18322 3652 18328 3664
rect 18187 3624 18328 3652
rect 18187 3621 18199 3624
rect 18141 3615 18199 3621
rect 18322 3612 18328 3624
rect 18380 3612 18386 3664
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 13814 3544 13820 3596
rect 13872 3544 13878 3596
rect 18432 3593 18460 3692
rect 19337 3689 19349 3723
rect 19383 3720 19395 3723
rect 19518 3720 19524 3732
rect 19383 3692 19524 3720
rect 19383 3689 19395 3692
rect 19337 3683 19395 3689
rect 19518 3680 19524 3692
rect 19576 3720 19582 3732
rect 20070 3720 20076 3732
rect 19576 3692 20076 3720
rect 19576 3680 19582 3692
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20714 3720 20720 3732
rect 20627 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3720 20778 3732
rect 21910 3720 21916 3732
rect 20772 3692 21916 3720
rect 20772 3680 20778 3692
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 24305 3723 24363 3729
rect 24305 3720 24317 3723
rect 24084 3692 24317 3720
rect 24084 3680 24090 3692
rect 24305 3689 24317 3692
rect 24351 3689 24363 3723
rect 24305 3683 24363 3689
rect 18779 3655 18837 3661
rect 18779 3621 18791 3655
rect 18825 3652 18837 3655
rect 19058 3652 19064 3664
rect 18825 3624 19064 3652
rect 18825 3621 18837 3624
rect 18779 3615 18837 3621
rect 19058 3612 19064 3624
rect 19116 3612 19122 3664
rect 20898 3652 20904 3664
rect 20859 3624 20904 3652
rect 20898 3612 20904 3624
rect 20956 3612 20962 3664
rect 18417 3587 18475 3593
rect 18417 3553 18429 3587
rect 18463 3553 18475 3587
rect 20990 3584 20996 3596
rect 20951 3556 20996 3584
rect 18417 3547 18475 3553
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 22554 3584 22560 3596
rect 22515 3556 22560 3584
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 24026 3544 24032 3596
rect 24084 3584 24090 3596
rect 24121 3587 24179 3593
rect 24121 3584 24133 3587
rect 24084 3556 24133 3584
rect 24084 3544 24090 3556
rect 24121 3553 24133 3556
rect 24167 3553 24179 3587
rect 24121 3547 24179 3553
rect 382 3476 388 3528
rect 440 3516 446 3528
rect 1302 3516 1308 3528
rect 440 3488 1308 3516
rect 440 3476 446 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 2332 3516 2360 3544
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 2332 3488 3433 3516
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 7282 3516 7288 3528
rect 7243 3488 7288 3516
rect 3421 3479 3479 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 7926 3516 7932 3528
rect 7883 3488 7932 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 7926 3476 7932 3488
rect 7984 3516 7990 3528
rect 8662 3516 8668 3528
rect 7984 3488 8668 3516
rect 7984 3476 7990 3488
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 15746 3516 15752 3528
rect 15707 3488 15752 3516
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 22462 3516 22468 3528
rect 22423 3488 22468 3516
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 3053 3451 3111 3457
rect 3053 3417 3065 3451
rect 3099 3448 3111 3451
rect 5721 3451 5779 3457
rect 3099 3420 3924 3448
rect 3099 3417 3111 3420
rect 3053 3411 3111 3417
rect 3896 3392 3924 3420
rect 5721 3417 5733 3451
rect 5767 3448 5779 3451
rect 6178 3448 6184 3460
rect 5767 3420 6184 3448
rect 5767 3417 5779 3420
rect 5721 3411 5779 3417
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 11698 3448 11704 3460
rect 11659 3420 11704 3448
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 1535 3383 1593 3389
rect 1535 3349 1547 3383
rect 1581 3380 1593 3383
rect 2130 3380 2136 3392
rect 1581 3352 2136 3380
rect 1581 3349 1593 3352
rect 1535 3343 1593 3349
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 3878 3380 3884 3392
rect 3839 3352 3884 3380
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 8294 3380 8300 3392
rect 8255 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 16666 3380 16672 3392
rect 16627 3352 16672 3380
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 19610 3380 19616 3392
rect 19571 3352 19616 3380
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 3234 3176 3240 3188
rect 3195 3148 3240 3176
rect 3234 3136 3240 3148
rect 3292 3176 3298 3188
rect 3418 3176 3424 3188
rect 3292 3148 3424 3176
rect 3292 3136 3298 3148
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5169 3179 5227 3185
rect 5169 3176 5181 3179
rect 4764 3148 5181 3176
rect 4764 3136 4770 3148
rect 5169 3145 5181 3148
rect 5215 3145 5227 3179
rect 5534 3176 5540 3188
rect 5495 3148 5540 3176
rect 5169 3139 5227 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 9953 3179 10011 3185
rect 9953 3145 9965 3179
rect 9999 3176 10011 3179
rect 10870 3176 10876 3188
rect 9999 3148 10876 3176
rect 9999 3145 10011 3148
rect 9953 3139 10011 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11882 3176 11888 3188
rect 11843 3148 11888 3176
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12526 3176 12532 3188
rect 12299 3148 12532 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 15013 3179 15071 3185
rect 15013 3176 15025 3179
rect 14792 3148 15025 3176
rect 14792 3136 14798 3148
rect 15013 3145 15025 3148
rect 15059 3145 15071 3179
rect 15013 3139 15071 3145
rect 15657 3179 15715 3185
rect 15657 3145 15669 3179
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 4893 3111 4951 3117
rect 4893 3077 4905 3111
rect 4939 3108 4951 3111
rect 5074 3108 5080 3120
rect 4939 3080 5080 3108
rect 4939 3077 4951 3080
rect 4893 3071 4951 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 11054 3108 11060 3120
rect 11015 3080 11060 3108
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3878 3040 3884 3052
rect 3007 3012 3884 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 7975 3012 8493 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8481 3009 8493 3012
rect 8527 3040 8539 3043
rect 8570 3040 8576 3052
rect 8527 3012 8576 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8754 3000 8760 3012
rect 8812 3040 8818 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 8812 3012 9505 3040
rect 8812 3000 8818 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 10502 3040 10508 3052
rect 10463 3012 10508 3040
rect 9493 3003 9551 3009
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 14752 3040 14780 3136
rect 15672 3108 15700 3139
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 15804 3148 17417 3176
rect 15804 3136 15810 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 17405 3139 17463 3145
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19518 3176 19524 3188
rect 19479 3148 19524 3176
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 20036 3148 20637 3176
rect 20036 3136 20042 3148
rect 20625 3145 20637 3148
rect 20671 3176 20683 3179
rect 22554 3176 22560 3188
rect 20671 3148 21312 3176
rect 22515 3148 22560 3176
rect 20671 3145 20683 3148
rect 20625 3139 20683 3145
rect 16117 3111 16175 3117
rect 16117 3108 16129 3111
rect 13863 3012 14780 3040
rect 15488 3080 16129 3108
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 5350 2972 5356 2984
rect 5311 2944 5356 2972
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2972 6331 2975
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6319 2944 6653 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 6641 2941 6653 2944
rect 6687 2972 6699 2975
rect 6730 2972 6736 2984
rect 6687 2944 6736 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 6730 2932 6736 2944
rect 6788 2972 6794 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 6788 2944 7481 2972
rect 6788 2932 6794 2944
rect 7469 2941 7481 2944
rect 7515 2972 7527 2975
rect 8202 2972 8208 2984
rect 7515 2944 8208 2972
rect 7515 2941 7527 2944
rect 7469 2935 7527 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12526 2972 12532 2984
rect 12483 2944 12532 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 12621 2975 12679 2981
rect 12621 2941 12633 2975
rect 12667 2972 12679 2975
rect 13262 2972 13268 2984
rect 12667 2944 13268 2972
rect 12667 2941 12679 2944
rect 12621 2935 12679 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14608 2944 14749 2972
rect 14608 2932 14614 2944
rect 14737 2941 14749 2944
rect 14783 2972 14795 2975
rect 15378 2972 15384 2984
rect 14783 2944 15384 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 2314 2904 2320 2916
rect 1811 2876 2320 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 2314 2864 2320 2876
rect 2372 2864 2378 2916
rect 2406 2864 2412 2916
rect 2464 2904 2470 2916
rect 3697 2907 3755 2913
rect 2464 2876 2509 2904
rect 2464 2864 2470 2876
rect 3697 2873 3709 2907
rect 3743 2904 3755 2907
rect 3970 2904 3976 2916
rect 3743 2876 3976 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4522 2904 4528 2916
rect 4483 2876 4528 2904
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2904 8355 2907
rect 8570 2904 8576 2916
rect 8343 2876 8576 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 10597 2907 10655 2913
rect 10597 2873 10609 2907
rect 10643 2904 10655 2907
rect 11698 2904 11704 2916
rect 10643 2876 11704 2904
rect 10643 2873 10655 2876
rect 10597 2867 10655 2873
rect 2133 2839 2191 2845
rect 2133 2805 2145 2839
rect 2179 2836 2191 2839
rect 2424 2836 2452 2864
rect 7098 2836 7104 2848
rect 2179 2808 2452 2836
rect 7059 2808 7104 2836
rect 2179 2805 2191 2808
rect 2133 2799 2191 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 10612 2836 10640 2867
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 13814 2904 13820 2916
rect 13771 2876 13820 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 11514 2836 11520 2848
rect 10367 2808 10640 2836
rect 11427 2808 11520 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 11514 2796 11520 2808
rect 11572 2836 11578 2848
rect 13740 2836 13768 2867
rect 13814 2864 13820 2876
rect 13872 2904 13878 2916
rect 14179 2907 14237 2913
rect 14179 2904 14191 2907
rect 13872 2876 14191 2904
rect 13872 2864 13878 2876
rect 14179 2873 14191 2876
rect 14225 2904 14237 2907
rect 15488 2904 15516 3080
rect 16117 3077 16129 3080
rect 16163 3108 16175 3111
rect 16482 3108 16488 3120
rect 16163 3080 16488 3108
rect 16163 3077 16175 3080
rect 16117 3071 16175 3077
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 19610 3068 19616 3120
rect 19668 3108 19674 3120
rect 19668 3080 19748 3108
rect 19668 3068 19674 3080
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 15712 3012 16221 3040
rect 15712 3000 15718 3012
rect 16209 3009 16221 3012
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 17368 3012 18153 3040
rect 17368 3000 17374 3012
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18141 3003 18199 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19720 3049 19748 3080
rect 21284 3049 21312 3148
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23566 3176 23572 3188
rect 23523 3148 23572 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 24084 3148 24685 3176
rect 24084 3136 24090 3148
rect 24673 3145 24685 3148
rect 24719 3145 24731 3179
rect 24673 3139 24731 3145
rect 24210 3068 24216 3120
rect 24268 3108 24274 3120
rect 25409 3111 25467 3117
rect 25409 3108 25421 3111
rect 24268 3080 25421 3108
rect 24268 3068 24274 3080
rect 25409 3077 25421 3080
rect 25455 3077 25467 3111
rect 25409 3071 25467 3077
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 17175 2944 17908 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 14225 2876 15516 2904
rect 14225 2873 14237 2876
rect 14179 2867 14237 2873
rect 16482 2864 16488 2916
rect 16540 2913 16546 2916
rect 16540 2907 16588 2913
rect 16540 2873 16542 2907
rect 16576 2873 16588 2907
rect 16540 2867 16588 2873
rect 16540 2864 16546 2867
rect 17880 2845 17908 2944
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 23624 2944 23765 2972
rect 23624 2932 23630 2944
rect 23753 2941 23765 2944
rect 23799 2941 23811 2975
rect 25222 2972 25228 2984
rect 25183 2944 25228 2972
rect 23753 2935 23811 2941
rect 25222 2932 25228 2944
rect 25280 2972 25286 2984
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 25280 2944 25789 2972
rect 25280 2932 25286 2944
rect 25777 2941 25789 2944
rect 25823 2941 25835 2975
rect 25777 2935 25835 2941
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 19797 2907 19855 2913
rect 18288 2876 18333 2904
rect 18288 2864 18294 2876
rect 19797 2873 19809 2907
rect 19843 2873 19855 2907
rect 19797 2867 19855 2873
rect 20349 2907 20407 2913
rect 20349 2873 20361 2907
rect 20395 2873 20407 2907
rect 20349 2867 20407 2873
rect 21085 2907 21143 2913
rect 21085 2873 21097 2907
rect 21131 2904 21143 2907
rect 21358 2904 21364 2916
rect 21131 2876 21364 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 11572 2808 13768 2836
rect 17865 2839 17923 2845
rect 11572 2796 11578 2808
rect 17865 2805 17877 2839
rect 17911 2836 17923 2839
rect 18248 2836 18276 2864
rect 17911 2808 18276 2836
rect 17911 2805 17923 2808
rect 17865 2799 17923 2805
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 19812 2836 19840 2867
rect 19576 2808 19840 2836
rect 20364 2836 20392 2867
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 21913 2907 21971 2913
rect 21913 2873 21925 2907
rect 21959 2873 21971 2907
rect 21913 2867 21971 2873
rect 21450 2836 21456 2848
rect 20364 2808 21456 2836
rect 19576 2796 19582 2808
rect 21450 2796 21456 2808
rect 21508 2836 21514 2848
rect 21928 2836 21956 2867
rect 23290 2864 23296 2916
rect 23348 2904 23354 2916
rect 23661 2907 23719 2913
rect 23661 2904 23673 2907
rect 23348 2876 23673 2904
rect 23348 2864 23354 2876
rect 23661 2873 23673 2876
rect 23707 2873 23719 2907
rect 23661 2867 23719 2873
rect 21508 2808 21956 2836
rect 21508 2796 21514 2808
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 3510 2632 3516 2644
rect 2363 2604 3516 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 2608 2573 2636 2604
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9214 2632 9220 2644
rect 9171 2604 9220 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2533 2651 2567
rect 2593 2527 2651 2533
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 3326 2564 3332 2576
rect 3191 2536 3332 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 3326 2524 3332 2536
rect 3384 2524 3390 2576
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4246 2564 4252 2576
rect 3927 2536 4252 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 6733 2567 6791 2573
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 7098 2564 7104 2576
rect 6779 2536 7104 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 1394 2456 1400 2508
rect 1452 2505 1458 2508
rect 1452 2499 1490 2505
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1452 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 6086 2496 6092 2508
rect 5675 2468 6092 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 1452 2456 1458 2459
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 9140 2496 9168 2595
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 9490 2592 9496 2604
rect 9548 2632 9554 2644
rect 13630 2632 13636 2644
rect 9548 2604 10456 2632
rect 9548 2592 9554 2604
rect 10428 2573 10456 2604
rect 12912 2604 13636 2632
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2533 10471 2567
rect 10413 2527 10471 2533
rect 10502 2524 10508 2576
rect 10560 2564 10566 2576
rect 10560 2536 10605 2564
rect 10560 2524 10566 2536
rect 11514 2524 11520 2576
rect 11572 2564 11578 2576
rect 12250 2564 12256 2576
rect 11572 2536 12256 2564
rect 11572 2524 11578 2536
rect 12250 2524 12256 2536
rect 12308 2524 12314 2576
rect 12912 2573 12940 2604
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 13814 2632 13820 2644
rect 13775 2604 13820 2632
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 19797 2635 19855 2641
rect 18187 2604 18552 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 18524 2576 18552 2604
rect 19797 2601 19809 2635
rect 19843 2632 19855 2635
rect 20438 2632 20444 2644
rect 19843 2604 20444 2632
rect 19843 2601 19855 2604
rect 19797 2595 19855 2601
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 12897 2567 12955 2573
rect 12897 2564 12909 2567
rect 12483 2536 12909 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 12897 2533 12909 2536
rect 12943 2533 12955 2567
rect 13446 2564 13452 2576
rect 13407 2536 13452 2564
rect 12897 2527 12955 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 15194 2524 15200 2576
rect 15252 2564 15258 2576
rect 15611 2567 15669 2573
rect 15611 2564 15623 2567
rect 15252 2536 15623 2564
rect 15252 2524 15258 2536
rect 15611 2533 15623 2536
rect 15657 2533 15669 2567
rect 15611 2527 15669 2533
rect 16393 2567 16451 2573
rect 16393 2533 16405 2567
rect 16439 2564 16451 2567
rect 16666 2564 16672 2576
rect 16439 2536 16672 2564
rect 16439 2533 16451 2536
rect 16393 2527 16451 2533
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 17218 2564 17224 2576
rect 17179 2536 17224 2564
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2564 17831 2567
rect 18046 2564 18052 2576
rect 17819 2536 18052 2564
rect 17819 2533 17831 2536
rect 17773 2527 17831 2533
rect 18046 2524 18052 2536
rect 18104 2564 18110 2576
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 18104 2536 18429 2564
rect 18104 2524 18110 2536
rect 18417 2533 18429 2536
rect 18463 2533 18475 2567
rect 18417 2527 18475 2533
rect 18506 2524 18512 2576
rect 18564 2564 18570 2576
rect 18564 2536 18609 2564
rect 18564 2524 18570 2536
rect 8527 2468 9168 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14312 2499 14370 2505
rect 14312 2496 14324 2499
rect 14148 2468 14324 2496
rect 14148 2456 14154 2468
rect 14312 2465 14324 2468
rect 14358 2496 14370 2499
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14358 2468 14749 2496
rect 14358 2465 14370 2468
rect 14312 2459 14370 2465
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 19904 2505 19932 2604
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 20990 2632 20996 2644
rect 20951 2604 20996 2632
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 23382 2632 23388 2644
rect 23343 2604 23388 2632
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 15508 2499 15566 2505
rect 15508 2496 15520 2499
rect 15436 2468 15520 2496
rect 15436 2456 15442 2468
rect 15508 2465 15520 2468
rect 15554 2496 15566 2499
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15554 2468 15945 2496
rect 15554 2465 15566 2468
rect 15508 2459 15566 2465
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 20530 2456 20536 2508
rect 20588 2496 20594 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 20588 2468 21281 2496
rect 20588 2456 20594 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 22741 2499 22799 2505
rect 22741 2465 22753 2499
rect 22787 2496 22799 2499
rect 23400 2496 23428 2592
rect 23842 2496 23848 2508
rect 22787 2468 23428 2496
rect 23755 2468 23848 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 23842 2456 23848 2468
rect 23900 2496 23906 2508
rect 24121 2499 24179 2505
rect 24121 2496 24133 2499
rect 23900 2468 24133 2496
rect 23900 2456 23906 2468
rect 24121 2465 24133 2468
rect 24167 2465 24179 2499
rect 24121 2459 24179 2465
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2096 2400 2513 2428
rect 2096 2388 2102 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 4154 2428 4160 2440
rect 3559 2400 4160 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4522 2428 4528 2440
rect 4483 2400 4528 2428
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7282 2428 7288 2440
rect 7243 2400 7288 2428
rect 7009 2391 7067 2397
rect 1535 2363 1593 2369
rect 1535 2329 1547 2363
rect 1581 2360 1593 2363
rect 2682 2360 2688 2372
rect 1581 2332 2688 2360
rect 1581 2329 1593 2332
rect 1535 2323 1593 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 6270 2360 6276 2372
rect 6231 2332 6276 2360
rect 6270 2320 6276 2332
rect 6328 2360 6334 2372
rect 7024 2360 7052 2391
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 11974 2428 11980 2440
rect 8628 2400 11376 2428
rect 11935 2400 11980 2428
rect 8628 2388 8634 2400
rect 10962 2360 10968 2372
rect 6328 2332 7052 2360
rect 10923 2332 10968 2360
rect 6328 2320 6334 2332
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 11348 2360 11376 2400
rect 11974 2388 11980 2400
rect 12032 2428 12038 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12032 2400 12817 2428
rect 12032 2388 12038 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 16577 2431 16635 2437
rect 16577 2428 16589 2431
rect 12805 2391 12863 2397
rect 15304 2400 16589 2428
rect 12158 2360 12164 2372
rect 11348 2332 12164 2360
rect 12158 2320 12164 2332
rect 12216 2320 12222 2372
rect 15304 2304 15332 2400
rect 16577 2397 16589 2400
rect 16623 2397 16635 2431
rect 18782 2428 18788 2440
rect 18743 2400 18788 2428
rect 16577 2391 16635 2397
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 21174 2428 21180 2440
rect 21135 2400 21180 2428
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 24026 2428 24032 2440
rect 23987 2400 24032 2428
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 25590 2428 25596 2440
rect 25551 2400 25596 2428
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 20073 2363 20131 2369
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 21082 2360 21088 2372
rect 20119 2332 21088 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 8662 2292 8668 2304
rect 8623 2264 8668 2292
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2292 10287 2295
rect 10502 2292 10508 2304
rect 10275 2264 10508 2292
rect 10275 2261 10287 2264
rect 10229 2255 10287 2261
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 14415 2295 14473 2301
rect 14415 2292 14427 2295
rect 13872 2264 14427 2292
rect 13872 2252 13878 2264
rect 14415 2261 14427 2264
rect 14461 2261 14473 2295
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 14415 2255 14473 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 20530 2292 20536 2304
rect 20491 2264 20536 2292
rect 20530 2252 20536 2264
rect 20588 2252 20594 2304
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 21968 2264 22937 2292
rect 21968 2252 21974 2264
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 6730 552 6736 604
rect 6788 592 6794 604
rect 7006 592 7012 604
rect 6788 564 7012 592
rect 6788 552 6794 564
rect 7006 552 7012 564
rect 7064 552 7070 604
rect 11422 552 11428 604
rect 11480 592 11486 604
rect 12342 592 12348 604
rect 11480 564 12348 592
rect 11480 552 11486 564
rect 12342 552 12348 564
rect 12400 552 12406 604
rect 14734 552 14740 604
rect 14792 592 14798 604
rect 14826 592 14832 604
rect 14792 564 14832 592
rect 14792 552 14798 564
rect 14826 552 14832 564
rect 14884 552 14890 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1492 24259 1544 24268
rect 1492 24225 1510 24259
rect 1510 24225 1544 24259
rect 1492 24216 1544 24225
rect 1768 24012 1820 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1492 23808 1544 23860
rect 1400 23647 1452 23656
rect 1400 23613 1444 23647
rect 1444 23613 1452 23647
rect 1400 23604 1452 23613
rect 1860 23468 1912 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22516 1636 22568
rect 2504 22380 2556 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21471 1544 21480
rect 1492 21437 1510 21471
rect 1510 21437 1544 21471
rect 1492 21428 1544 21437
rect 1584 21292 1636 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1400 20995 1452 21004
rect 1400 20961 1444 20995
rect 1444 20961 1452 20995
rect 1400 20952 1452 20961
rect 1676 20748 1728 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20544 1452 20596
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1492 19907 1544 19916
rect 1492 19873 1510 19907
rect 1510 19873 1544 19907
rect 1492 19864 1544 19873
rect 2596 19660 2648 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1492 19456 1544 19508
rect 1952 19320 2004 19372
rect 3332 19320 3384 19372
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 5540 18776 5592 18828
rect 6276 18572 6328 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 5540 18368 5592 18420
rect 1584 18164 1636 18216
rect 1492 18028 1544 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1400 17731 1452 17740
rect 1400 17697 1444 17731
rect 1444 17697 1452 17731
rect 1400 17688 1452 17697
rect 2964 17688 3016 17740
rect 11152 17731 11204 17740
rect 11152 17697 11196 17731
rect 11196 17697 11204 17731
rect 11152 17688 11204 17697
rect 2412 17552 2464 17604
rect 2136 17527 2188 17536
rect 2136 17493 2145 17527
rect 2145 17493 2179 17527
rect 2179 17493 2188 17527
rect 2136 17484 2188 17493
rect 2596 17484 2648 17536
rect 12164 17484 12216 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 11152 17323 11204 17332
rect 11152 17289 11161 17323
rect 11161 17289 11195 17323
rect 11195 17289 11204 17323
rect 11152 17280 11204 17289
rect 2136 17119 2188 17128
rect 2136 17085 2145 17119
rect 2145 17085 2179 17119
rect 2179 17085 2188 17119
rect 2136 17076 2188 17085
rect 3516 17076 3568 17128
rect 2044 17051 2096 17060
rect 2044 17017 2053 17051
rect 2053 17017 2087 17051
rect 2087 17017 2096 17051
rect 2044 17008 2096 17017
rect 1400 16940 1452 16992
rect 2964 16940 3016 16992
rect 3240 16940 3292 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3884 16668 3936 16720
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 1676 16532 1728 16584
rect 4344 16600 4396 16652
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 3884 16056 3936 16108
rect 1676 15852 1728 15904
rect 2228 15895 2280 15904
rect 2228 15861 2237 15895
rect 2237 15861 2271 15895
rect 2271 15861 2280 15895
rect 2228 15852 2280 15861
rect 2596 15895 2648 15904
rect 2596 15861 2605 15895
rect 2605 15861 2639 15895
rect 2639 15861 2648 15895
rect 2596 15852 2648 15861
rect 3424 15852 3476 15904
rect 4252 15852 4304 15904
rect 4988 15852 5040 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1216 15648 1268 15700
rect 1860 15648 1912 15700
rect 1860 15512 1912 15564
rect 4620 15555 4672 15564
rect 4620 15521 4629 15555
rect 4629 15521 4663 15555
rect 4663 15521 4672 15555
rect 4620 15512 4672 15521
rect 10140 15512 10192 15564
rect 15476 15512 15528 15564
rect 4528 15487 4580 15496
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 6184 15444 6236 15496
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2136 15308 2188 15317
rect 10692 15308 10744 15360
rect 16304 15308 16356 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 10140 15104 10192 15156
rect 15476 15104 15528 15156
rect 1400 14900 1452 14952
rect 4068 14900 4120 14952
rect 5264 14900 5316 14952
rect 6092 14832 6144 14884
rect 1860 14764 1912 14816
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5080 14764 5132 14816
rect 8024 14764 8076 14816
rect 9956 14900 10008 14952
rect 9128 14764 9180 14816
rect 10140 14764 10192 14816
rect 11520 14764 11572 14816
rect 12348 14764 12400 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2688 14424 2740 14476
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 5448 14467 5500 14476
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 8944 14424 8996 14476
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 11888 14424 11940 14476
rect 15568 14467 15620 14476
rect 15568 14433 15612 14467
rect 15612 14433 15620 14467
rect 15568 14424 15620 14433
rect 5172 14356 5224 14408
rect 7380 14356 7432 14408
rect 1400 14288 1452 14340
rect 1768 14220 1820 14272
rect 2780 14220 2832 14272
rect 5264 14220 5316 14272
rect 5540 14220 5592 14272
rect 8852 14220 8904 14272
rect 11428 14220 11480 14272
rect 11980 14220 12032 14272
rect 15936 14220 15988 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1124 14016 1176 14068
rect 1492 14016 1544 14068
rect 3056 14016 3108 14068
rect 3792 14059 3844 14068
rect 3792 14025 3801 14059
rect 3801 14025 3835 14059
rect 3835 14025 3844 14059
rect 3792 14016 3844 14025
rect 4528 14016 4580 14068
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 7012 14016 7064 14068
rect 3148 13948 3200 14000
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 5264 13948 5316 14000
rect 7472 14016 7524 14068
rect 10508 14016 10560 14068
rect 10876 14016 10928 14068
rect 7288 13948 7340 14000
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 7472 13812 7524 13864
rect 4160 13744 4212 13796
rect 4528 13787 4580 13796
rect 4528 13753 4537 13787
rect 4537 13753 4571 13787
rect 4571 13753 4580 13787
rect 4528 13744 4580 13753
rect 5448 13744 5500 13796
rect 8300 13812 8352 13864
rect 10692 13948 10744 14000
rect 12900 14016 12952 14068
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 12716 13948 12768 14000
rect 9036 13880 9088 13932
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 9864 13812 9916 13864
rect 8760 13744 8812 13796
rect 11888 13812 11940 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13636 13812 13688 13864
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 10784 13744 10836 13796
rect 1768 13676 1820 13728
rect 2136 13676 2188 13728
rect 7104 13719 7156 13728
rect 7104 13685 7113 13719
rect 7113 13685 7147 13719
rect 7147 13685 7156 13719
rect 7104 13676 7156 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 4160 13472 4212 13524
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 2136 13447 2188 13456
rect 2136 13413 2145 13447
rect 2145 13413 2179 13447
rect 2179 13413 2188 13447
rect 2136 13404 2188 13413
rect 5540 13447 5592 13456
rect 5540 13413 5549 13447
rect 5549 13413 5583 13447
rect 5583 13413 5592 13447
rect 5540 13404 5592 13413
rect 7012 13404 7064 13456
rect 4160 13379 4212 13388
rect 4160 13345 4178 13379
rect 4178 13345 4212 13379
rect 4160 13336 4212 13345
rect 1216 13268 1268 13320
rect 1124 13200 1176 13252
rect 2320 13200 2372 13252
rect 8668 13336 8720 13388
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 11796 13379 11848 13388
rect 9680 13336 9732 13345
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 14004 13379 14056 13388
rect 5172 13268 5224 13320
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 11152 13268 11204 13320
rect 14004 13345 14013 13379
rect 14013 13345 14047 13379
rect 14047 13345 14056 13379
rect 14004 13336 14056 13345
rect 15384 13379 15436 13388
rect 15384 13345 15428 13379
rect 15428 13345 15436 13379
rect 15384 13336 15436 13345
rect 13452 13268 13504 13320
rect 3056 13175 3108 13184
rect 3056 13141 3065 13175
rect 3065 13141 3099 13175
rect 3099 13141 3108 13175
rect 3056 13132 3108 13141
rect 4896 13175 4948 13184
rect 4896 13141 4905 13175
rect 4905 13141 4939 13175
rect 4939 13141 4948 13175
rect 4896 13132 4948 13141
rect 9772 13132 9824 13184
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 13360 13132 13412 13184
rect 14648 13132 14700 13184
rect 16396 13132 16448 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1768 12928 1820 12980
rect 2136 12928 2188 12980
rect 1216 12860 1268 12912
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 5540 12928 5592 12980
rect 6920 12928 6972 12980
rect 7196 12928 7248 12980
rect 11520 12928 11572 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 14004 12928 14056 12980
rect 15384 12928 15436 12980
rect 2688 12860 2740 12912
rect 5448 12903 5500 12912
rect 5448 12869 5457 12903
rect 5457 12869 5491 12903
rect 5491 12869 5500 12903
rect 5448 12860 5500 12869
rect 7012 12860 7064 12912
rect 8668 12903 8720 12912
rect 8668 12869 8677 12903
rect 8677 12869 8711 12903
rect 8711 12869 8720 12903
rect 8668 12860 8720 12869
rect 10876 12860 10928 12912
rect 3056 12792 3108 12844
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 5356 12792 5408 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 7748 12792 7800 12844
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 14556 12792 14608 12844
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 10232 12724 10284 12776
rect 10876 12724 10928 12776
rect 12808 12724 12860 12776
rect 14096 12724 14148 12776
rect 16028 12767 16080 12776
rect 16028 12733 16072 12767
rect 16072 12733 16080 12767
rect 16028 12724 16080 12733
rect 1124 12656 1176 12708
rect 1676 12656 1728 12708
rect 1768 12656 1820 12708
rect 4620 12656 4672 12708
rect 1216 12588 1268 12640
rect 1400 12588 1452 12640
rect 5172 12656 5224 12708
rect 7656 12699 7708 12708
rect 7656 12665 7665 12699
rect 7665 12665 7699 12699
rect 7699 12665 7708 12699
rect 7656 12656 7708 12665
rect 7748 12699 7800 12708
rect 7748 12665 7757 12699
rect 7757 12665 7791 12699
rect 7791 12665 7800 12699
rect 7748 12656 7800 12665
rect 10416 12656 10468 12708
rect 11152 12656 11204 12708
rect 13176 12699 13228 12708
rect 13176 12665 13185 12699
rect 13185 12665 13219 12699
rect 13219 12665 13228 12699
rect 13176 12656 13228 12665
rect 13544 12656 13596 12708
rect 5908 12588 5960 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 10048 12588 10100 12640
rect 11520 12588 11572 12640
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 16212 12588 16264 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 5908 12427 5960 12436
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 7196 12384 7248 12436
rect 8668 12384 8720 12436
rect 9680 12384 9732 12436
rect 9772 12384 9824 12436
rect 12532 12384 12584 12436
rect 14188 12384 14240 12436
rect 2044 12316 2096 12368
rect 2688 12359 2740 12368
rect 2688 12325 2697 12359
rect 2697 12325 2731 12359
rect 2731 12325 2740 12359
rect 2688 12316 2740 12325
rect 5172 12316 5224 12368
rect 7012 12316 7064 12368
rect 11060 12316 11112 12368
rect 11612 12359 11664 12368
rect 11612 12325 11621 12359
rect 11621 12325 11655 12359
rect 11655 12325 11664 12359
rect 11612 12316 11664 12325
rect 13176 12359 13228 12368
rect 13176 12325 13185 12359
rect 13185 12325 13219 12359
rect 13219 12325 13228 12359
rect 13176 12316 13228 12325
rect 9772 12291 9824 12300
rect 9772 12257 9781 12291
rect 9781 12257 9815 12291
rect 9815 12257 9824 12291
rect 9772 12248 9824 12257
rect 15384 12291 15436 12300
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 2136 12180 2188 12232
rect 6092 12180 6144 12232
rect 7104 12180 7156 12232
rect 7472 12180 7524 12232
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9588 12180 9640 12232
rect 10876 12180 10928 12232
rect 11336 12180 11388 12232
rect 12164 12180 12216 12232
rect 13728 12180 13780 12232
rect 12348 12112 12400 12164
rect 14004 12112 14056 12164
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 2872 12044 2924 12096
rect 3424 12044 3476 12096
rect 7840 12044 7892 12096
rect 10876 12044 10928 12096
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 2136 11840 2188 11892
rect 6092 11883 6144 11892
rect 6092 11849 6101 11883
rect 6101 11849 6135 11883
rect 6135 11849 6144 11883
rect 6092 11840 6144 11849
rect 9772 11883 9824 11892
rect 9772 11849 9781 11883
rect 9781 11849 9815 11883
rect 9815 11849 9824 11883
rect 9772 11840 9824 11849
rect 11612 11840 11664 11892
rect 12624 11840 12676 11892
rect 13176 11840 13228 11892
rect 13728 11840 13780 11892
rect 15384 11840 15436 11892
rect 11428 11772 11480 11824
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 7012 11704 7064 11756
rect 7656 11704 7708 11756
rect 7932 11704 7984 11756
rect 10048 11704 10100 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 1676 11636 1728 11688
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2872 11611 2924 11620
rect 2872 11577 2881 11611
rect 2881 11577 2915 11611
rect 2915 11577 2924 11611
rect 2872 11568 2924 11577
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 12532 11679 12584 11688
rect 5172 11611 5224 11620
rect 5172 11577 5175 11611
rect 5175 11577 5209 11611
rect 5209 11577 5224 11611
rect 5172 11568 5224 11577
rect 7196 11611 7248 11620
rect 7196 11577 7205 11611
rect 7205 11577 7239 11611
rect 7239 11577 7248 11611
rect 7196 11568 7248 11577
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 9404 11611 9456 11620
rect 7288 11568 7340 11577
rect 9404 11577 9413 11611
rect 9413 11577 9447 11611
rect 9447 11577 9456 11611
rect 9404 11568 9456 11577
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 12532 11645 12541 11679
rect 12541 11645 12575 11679
rect 12575 11645 12584 11679
rect 12532 11636 12584 11645
rect 10692 11568 10744 11620
rect 12900 11568 12952 11620
rect 13360 11568 13412 11620
rect 12624 11500 12676 11552
rect 16120 11568 16172 11620
rect 16304 11611 16356 11620
rect 16304 11577 16313 11611
rect 16313 11577 16347 11611
rect 16347 11577 16356 11611
rect 16304 11568 16356 11577
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11296 1728 11348
rect 2504 11296 2556 11348
rect 5540 11296 5592 11348
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 7472 11339 7524 11348
rect 7472 11305 7481 11339
rect 7481 11305 7515 11339
rect 7515 11305 7524 11339
rect 7472 11296 7524 11305
rect 10048 11296 10100 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 12992 11296 13044 11348
rect 13452 11296 13504 11348
rect 13636 11296 13688 11348
rect 4252 11228 4304 11280
rect 5172 11271 5224 11280
rect 5172 11237 5175 11271
rect 5175 11237 5209 11271
rect 5209 11237 5224 11271
rect 5172 11228 5224 11237
rect 1676 11160 1728 11212
rect 2044 11160 2096 11212
rect 2872 11160 2924 11212
rect 3516 11160 3568 11212
rect 7564 11228 7616 11280
rect 7288 11160 7340 11212
rect 9404 11228 9456 11280
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 10784 11228 10836 11280
rect 10876 11228 10928 11280
rect 3332 11092 3384 11144
rect 4160 11092 4212 11144
rect 5448 11092 5500 11144
rect 8484 11092 8536 11144
rect 10876 11092 10928 11144
rect 2136 11024 2188 11076
rect 6736 11067 6788 11076
rect 6736 11033 6745 11067
rect 6745 11033 6779 11067
rect 6779 11033 6788 11067
rect 6736 11024 6788 11033
rect 10048 11024 10100 11076
rect 12164 11228 12216 11280
rect 13820 11271 13872 11280
rect 13820 11237 13829 11271
rect 13829 11237 13863 11271
rect 13863 11237 13872 11271
rect 13820 11228 13872 11237
rect 14832 11228 14884 11280
rect 16304 11228 16356 11280
rect 16120 11160 16172 11212
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 18512 11203 18564 11212
rect 16948 11160 17000 11169
rect 18512 11169 18530 11203
rect 18530 11169 18564 11203
rect 18512 11160 18564 11169
rect 14004 11135 14056 11144
rect 11704 11067 11756 11076
rect 11704 11033 11713 11067
rect 11713 11033 11747 11067
rect 11747 11033 11756 11067
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 14740 11092 14792 11144
rect 11704 11024 11756 11033
rect 12992 11024 13044 11076
rect 14556 11024 14608 11076
rect 20168 11024 20220 11076
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 10784 10956 10836 11008
rect 11152 10956 11204 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 3700 10752 3752 10804
rect 4068 10752 4120 10804
rect 5172 10752 5224 10804
rect 5448 10752 5500 10804
rect 7564 10752 7616 10804
rect 9404 10752 9456 10804
rect 10692 10752 10744 10804
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11796 10752 11848 10804
rect 12440 10752 12492 10804
rect 12808 10752 12860 10804
rect 13728 10752 13780 10804
rect 14832 10752 14884 10804
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 1216 10616 1268 10668
rect 1400 10616 1452 10668
rect 2504 10616 2556 10668
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 1952 10523 2004 10532
rect 1952 10489 1961 10523
rect 1961 10489 1995 10523
rect 1995 10489 2004 10523
rect 1952 10480 2004 10489
rect 2504 10523 2556 10532
rect 2504 10489 2513 10523
rect 2513 10489 2547 10523
rect 2547 10489 2556 10523
rect 2504 10480 2556 10489
rect 3516 10548 3568 10600
rect 5172 10591 5224 10600
rect 4068 10480 4120 10532
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 2872 10455 2924 10464
rect 2872 10421 2881 10455
rect 2881 10421 2915 10455
rect 2915 10421 2924 10455
rect 2872 10412 2924 10421
rect 3424 10412 3476 10464
rect 4804 10412 4856 10464
rect 8760 10548 8812 10600
rect 9220 10548 9272 10600
rect 7656 10480 7708 10532
rect 12164 10684 12216 10736
rect 12348 10684 12400 10736
rect 13176 10684 13228 10736
rect 16488 10727 16540 10736
rect 16488 10693 16497 10727
rect 16497 10693 16531 10727
rect 16531 10693 16540 10727
rect 16488 10684 16540 10693
rect 13544 10616 13596 10668
rect 13820 10548 13872 10600
rect 16856 10548 16908 10600
rect 13176 10523 13228 10532
rect 6460 10412 6512 10464
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 12440 10412 12492 10464
rect 13176 10489 13185 10523
rect 13185 10489 13219 10523
rect 13219 10489 13228 10523
rect 13176 10480 13228 10489
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 15752 10412 15804 10464
rect 17684 10480 17736 10532
rect 18512 10480 18564 10532
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2044 10208 2096 10260
rect 3516 10208 3568 10260
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 4896 10208 4948 10260
rect 5540 10208 5592 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 12440 10208 12492 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 13544 10208 13596 10260
rect 2688 10140 2740 10192
rect 7104 10140 7156 10192
rect 3424 10072 3476 10124
rect 5080 10072 5132 10124
rect 5264 10072 5316 10124
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 3516 10047 3568 10056
rect 3516 10013 3525 10047
rect 3525 10013 3559 10047
rect 3559 10013 3568 10047
rect 3516 10004 3568 10013
rect 4160 10004 4212 10056
rect 6184 10072 6236 10124
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 10692 10140 10744 10192
rect 10968 10140 11020 10192
rect 12164 10140 12216 10192
rect 14004 10140 14056 10192
rect 14740 10208 14792 10260
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 15384 10140 15436 10192
rect 16488 10140 16540 10192
rect 8760 10072 8812 10124
rect 9312 10072 9364 10124
rect 10876 10072 10928 10124
rect 17500 10140 17552 10192
rect 17776 10072 17828 10124
rect 19064 10115 19116 10124
rect 19064 10081 19073 10115
rect 19073 10081 19107 10115
rect 19107 10081 19116 10115
rect 19064 10072 19116 10081
rect 23480 10072 23532 10124
rect 8576 10004 8628 10056
rect 13452 10047 13504 10056
rect 2780 9936 2832 9988
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 15752 10004 15804 10056
rect 16488 10004 16540 10056
rect 17960 10004 18012 10056
rect 13820 9936 13872 9988
rect 1768 9868 1820 9920
rect 2872 9868 2924 9920
rect 3240 9868 3292 9920
rect 9220 9868 9272 9920
rect 11428 9868 11480 9920
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 24124 9868 24176 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2320 9664 2372 9716
rect 2688 9707 2740 9716
rect 2688 9673 2697 9707
rect 2697 9673 2731 9707
rect 2731 9673 2740 9707
rect 2688 9664 2740 9673
rect 2872 9664 2924 9716
rect 1584 9596 1636 9648
rect 1216 9528 1268 9580
rect 2044 9596 2096 9648
rect 3240 9596 3292 9648
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3516 9460 3568 9512
rect 6460 9664 6512 9716
rect 5540 9596 5592 9648
rect 7104 9664 7156 9716
rect 9220 9707 9272 9716
rect 9220 9673 9229 9707
rect 9229 9673 9263 9707
rect 9263 9673 9272 9707
rect 9220 9664 9272 9673
rect 10876 9664 10928 9716
rect 12164 9664 12216 9716
rect 14004 9664 14056 9716
rect 15384 9664 15436 9716
rect 6920 9596 6972 9648
rect 7380 9596 7432 9648
rect 4804 9528 4856 9580
rect 7380 9460 7432 9512
rect 7932 9460 7984 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 8668 9460 8720 9512
rect 10968 9596 11020 9648
rect 17500 9664 17552 9716
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 19064 9707 19116 9716
rect 19064 9673 19073 9707
rect 19073 9673 19107 9707
rect 19107 9673 19116 9707
rect 19064 9664 19116 9673
rect 23480 9707 23532 9716
rect 23480 9673 23489 9707
rect 23489 9673 23523 9707
rect 23523 9673 23532 9707
rect 23480 9664 23532 9673
rect 11704 9528 11756 9580
rect 13820 9528 13872 9580
rect 2044 9392 2096 9444
rect 2136 9392 2188 9444
rect 2504 9392 2556 9444
rect 2688 9392 2740 9444
rect 3884 9435 3936 9444
rect 3884 9401 3893 9435
rect 3893 9401 3927 9435
rect 3927 9401 3936 9435
rect 3884 9392 3936 9401
rect 5080 9435 5132 9444
rect 5080 9401 5083 9435
rect 5083 9401 5117 9435
rect 5117 9401 5132 9435
rect 5080 9392 5132 9401
rect 9312 9392 9364 9444
rect 12716 9460 12768 9512
rect 13084 9460 13136 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 14188 9460 14240 9512
rect 16396 9596 16448 9648
rect 20168 9596 20220 9648
rect 20444 9596 20496 9648
rect 14924 9460 14976 9512
rect 17224 9460 17276 9512
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 19156 9460 19208 9512
rect 21272 9503 21324 9512
rect 21272 9469 21290 9503
rect 21290 9469 21324 9503
rect 21272 9460 21324 9469
rect 23664 9503 23716 9512
rect 23664 9469 23708 9503
rect 23708 9469 23716 9503
rect 23664 9460 23716 9469
rect 15568 9435 15620 9444
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 15568 9392 15620 9401
rect 2964 9324 3016 9376
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 6184 9324 6236 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 17868 9392 17920 9444
rect 20352 9435 20404 9444
rect 20352 9401 20361 9435
rect 20361 9401 20395 9435
rect 20395 9401 20404 9435
rect 20352 9392 20404 9401
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 18236 9324 18288 9376
rect 21548 9324 21600 9376
rect 24032 9324 24084 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 3884 9120 3936 9172
rect 1124 9052 1176 9104
rect 2044 9052 2096 9104
rect 2504 9052 2556 9104
rect 2780 9052 2832 9104
rect 8392 9120 8444 9172
rect 9588 9120 9640 9172
rect 10784 9163 10836 9172
rect 10784 9129 10793 9163
rect 10793 9129 10827 9163
rect 10827 9129 10836 9163
rect 10784 9120 10836 9129
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 5080 9052 5132 9104
rect 10232 9052 10284 9104
rect 10876 9052 10928 9104
rect 10968 9052 11020 9104
rect 11152 9052 11204 9104
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 11888 9052 11940 9104
rect 13452 9052 13504 9104
rect 14096 9052 14148 9104
rect 16580 9095 16632 9104
rect 16580 9061 16589 9095
rect 16589 9061 16623 9095
rect 16623 9061 16632 9095
rect 16580 9052 16632 9061
rect 16764 9120 16816 9172
rect 18972 9120 19024 9172
rect 19156 9163 19208 9172
rect 19156 9129 19165 9163
rect 19165 9129 19199 9163
rect 19199 9129 19208 9163
rect 19156 9120 19208 9129
rect 17224 9095 17276 9104
rect 17224 9061 17233 9095
rect 17233 9061 17267 9095
rect 17267 9061 17276 9095
rect 17224 9052 17276 9061
rect 18328 9052 18380 9104
rect 11704 8984 11756 9036
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 13360 9027 13412 9036
rect 13360 8993 13369 9027
rect 13369 8993 13403 9027
rect 13403 8993 13412 9027
rect 13360 8984 13412 8993
rect 21916 9027 21968 9036
rect 21916 8993 21960 9027
rect 21960 8993 21968 9027
rect 21916 8984 21968 8993
rect 2688 8916 2740 8968
rect 3148 8916 3200 8968
rect 6276 8916 6328 8968
rect 8484 8916 8536 8968
rect 9220 8916 9272 8968
rect 10692 8916 10744 8968
rect 10968 8916 11020 8968
rect 13728 8916 13780 8968
rect 15936 8916 15988 8968
rect 17868 8916 17920 8968
rect 19616 8959 19668 8968
rect 6000 8848 6052 8900
rect 7380 8848 7432 8900
rect 9588 8848 9640 8900
rect 11520 8848 11572 8900
rect 17960 8848 18012 8900
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 1860 8780 1912 8832
rect 2044 8780 2096 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 12440 8780 12492 8832
rect 13176 8780 13228 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 22008 8780 22060 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2320 8576 2372 8628
rect 2872 8576 2924 8628
rect 5356 8576 5408 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 10232 8576 10284 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 12900 8619 12952 8628
rect 8392 8508 8444 8560
rect 9128 8508 9180 8560
rect 9404 8508 9456 8560
rect 10692 8508 10744 8560
rect 10876 8551 10928 8560
rect 10876 8517 10885 8551
rect 10885 8517 10919 8551
rect 10919 8517 10928 8551
rect 10876 8508 10928 8517
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 4068 8440 4120 8492
rect 5448 8440 5500 8492
rect 6000 8440 6052 8492
rect 6920 8440 6972 8492
rect 7748 8440 7800 8492
rect 9220 8440 9272 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 4160 8415 4212 8424
rect 4160 8381 4169 8415
rect 4169 8381 4203 8415
rect 4203 8381 4212 8415
rect 4160 8372 4212 8381
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 10784 8372 10836 8424
rect 2320 8304 2372 8356
rect 3332 8304 3384 8356
rect 4344 8347 4396 8356
rect 4344 8313 4353 8347
rect 4353 8313 4387 8347
rect 4387 8313 4396 8347
rect 4344 8304 4396 8313
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 7104 8304 7156 8356
rect 7656 8304 7708 8356
rect 10232 8304 10284 8356
rect 11520 8304 11572 8356
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 13268 8619 13320 8628
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 14004 8576 14056 8628
rect 12808 8551 12860 8560
rect 12808 8517 12832 8551
rect 12832 8517 12860 8551
rect 12808 8508 12860 8517
rect 12440 8440 12492 8492
rect 16580 8576 16632 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18328 8576 18380 8628
rect 20352 8576 20404 8628
rect 20812 8576 20864 8628
rect 15752 8508 15804 8560
rect 16764 8551 16816 8560
rect 15568 8440 15620 8492
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 14280 8372 14332 8424
rect 14832 8372 14884 8424
rect 5080 8236 5132 8288
rect 7196 8236 7248 8288
rect 13544 8304 13596 8356
rect 16764 8517 16773 8551
rect 16773 8517 16807 8551
rect 16807 8517 16816 8551
rect 16764 8508 16816 8517
rect 18420 8508 18472 8560
rect 21272 8551 21324 8560
rect 21272 8517 21281 8551
rect 21281 8517 21315 8551
rect 21315 8517 21324 8551
rect 21272 8508 21324 8517
rect 17224 8440 17276 8492
rect 19340 8440 19392 8492
rect 19616 8440 19668 8492
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 16304 8372 16356 8424
rect 22100 8372 22152 8424
rect 10784 8236 10836 8288
rect 12440 8236 12492 8288
rect 19156 8304 19208 8356
rect 20812 8347 20864 8356
rect 20812 8313 20821 8347
rect 20821 8313 20855 8347
rect 20855 8313 20864 8347
rect 20812 8304 20864 8313
rect 21456 8304 21508 8356
rect 21916 8347 21968 8356
rect 21916 8313 21925 8347
rect 21925 8313 21959 8347
rect 21959 8313 21968 8347
rect 21916 8304 21968 8313
rect 23296 8304 23348 8356
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2044 8032 2096 8084
rect 2688 8032 2740 8084
rect 4068 8032 4120 8084
rect 5540 8032 5592 8084
rect 6828 8032 6880 8084
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 9588 8032 9640 8084
rect 11888 8032 11940 8084
rect 13360 8032 13412 8084
rect 15568 8032 15620 8084
rect 1584 7964 1636 8016
rect 2228 7964 2280 8016
rect 2780 8007 2832 8016
rect 2780 7973 2789 8007
rect 2789 7973 2823 8007
rect 2823 7973 2832 8007
rect 5080 8007 5132 8016
rect 2780 7964 2832 7973
rect 5080 7973 5083 8007
rect 5083 7973 5117 8007
rect 5117 7973 5132 8007
rect 5080 7964 5132 7973
rect 9312 7964 9364 8016
rect 10048 7964 10100 8016
rect 19156 8032 19208 8084
rect 19340 8075 19392 8084
rect 19340 8041 19349 8075
rect 19349 8041 19383 8075
rect 19383 8041 19392 8075
rect 19340 8032 19392 8041
rect 19432 8032 19484 8084
rect 20720 8075 20772 8084
rect 20720 8041 20729 8075
rect 20729 8041 20763 8075
rect 20763 8041 20772 8075
rect 20720 8032 20772 8041
rect 16672 8007 16724 8016
rect 4896 7896 4948 7948
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 7932 7939 7984 7948
rect 7932 7905 7941 7939
rect 7941 7905 7975 7939
rect 7975 7905 7984 7939
rect 7932 7896 7984 7905
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 8576 7896 8628 7948
rect 10784 7896 10836 7948
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3240 7828 3292 7880
rect 8300 7828 8352 7880
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 16672 7964 16724 7973
rect 16856 7964 16908 8016
rect 17960 7964 18012 8016
rect 18420 7964 18472 8016
rect 11704 7828 11756 7837
rect 2412 7760 2464 7812
rect 2688 7760 2740 7812
rect 1860 7692 1912 7744
rect 9864 7760 9916 7812
rect 10048 7760 10100 7812
rect 10692 7760 10744 7812
rect 10876 7803 10928 7812
rect 10876 7769 10885 7803
rect 10885 7769 10919 7803
rect 10919 7769 10928 7803
rect 10876 7760 10928 7769
rect 11060 7803 11112 7812
rect 11060 7769 11069 7803
rect 11069 7769 11103 7803
rect 11103 7769 11112 7803
rect 11060 7760 11112 7769
rect 12348 7760 12400 7812
rect 12900 7896 12952 7948
rect 16304 7896 16356 7948
rect 20996 7939 21048 7948
rect 20996 7905 21005 7939
rect 21005 7905 21039 7939
rect 21039 7905 21048 7939
rect 20996 7896 21048 7905
rect 22468 7939 22520 7948
rect 22468 7905 22477 7939
rect 22477 7905 22511 7939
rect 22511 7905 22520 7939
rect 22468 7896 22520 7905
rect 23572 7939 23624 7948
rect 23572 7905 23590 7939
rect 23590 7905 23624 7939
rect 23572 7896 23624 7905
rect 13360 7828 13412 7880
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 16856 7828 16908 7880
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 20812 7828 20864 7880
rect 17040 7760 17092 7812
rect 5540 7692 5592 7744
rect 11244 7692 11296 7744
rect 13176 7735 13228 7744
rect 13176 7701 13185 7735
rect 13185 7701 13219 7735
rect 13219 7701 13228 7735
rect 13176 7692 13228 7701
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 21272 7692 21324 7744
rect 22192 7692 22244 7744
rect 23388 7692 23440 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2228 7488 2280 7540
rect 1584 7420 1636 7472
rect 4896 7488 4948 7540
rect 9404 7488 9456 7540
rect 10876 7488 10928 7540
rect 12348 7488 12400 7540
rect 12808 7488 12860 7540
rect 2504 7420 2556 7472
rect 3700 7420 3752 7472
rect 5080 7420 5132 7472
rect 10784 7420 10836 7472
rect 11060 7420 11112 7472
rect 1400 7216 1452 7268
rect 2228 7216 2280 7268
rect 3516 7352 3568 7404
rect 4344 7352 4396 7404
rect 11428 7352 11480 7404
rect 12900 7352 12952 7404
rect 3148 7148 3200 7200
rect 7932 7284 7984 7336
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 8668 7284 8720 7336
rect 8760 7284 8812 7336
rect 5080 7259 5132 7268
rect 5080 7225 5083 7259
rect 5083 7225 5117 7259
rect 5117 7225 5132 7259
rect 5080 7216 5132 7225
rect 11060 7284 11112 7336
rect 13452 7488 13504 7540
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 20720 7488 20772 7540
rect 22468 7488 22520 7540
rect 14188 7352 14240 7404
rect 16488 7352 16540 7404
rect 18144 7352 18196 7404
rect 19432 7352 19484 7404
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 21732 7395 21784 7404
rect 21732 7361 21741 7395
rect 21741 7361 21775 7395
rect 21775 7361 21784 7395
rect 21732 7352 21784 7361
rect 23572 7352 23624 7404
rect 14280 7327 14332 7336
rect 10968 7216 11020 7268
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 14648 7284 14700 7336
rect 18328 7284 18380 7336
rect 11888 7259 11940 7268
rect 11888 7225 11897 7259
rect 11897 7225 11931 7259
rect 11931 7225 11940 7259
rect 11888 7216 11940 7225
rect 13728 7216 13780 7268
rect 15752 7216 15804 7268
rect 7656 7191 7708 7200
rect 7656 7157 7665 7191
rect 7665 7157 7699 7191
rect 7699 7157 7708 7191
rect 7656 7148 7708 7157
rect 9128 7148 9180 7200
rect 13820 7148 13872 7200
rect 17408 7216 17460 7268
rect 20720 7284 20772 7336
rect 21272 7327 21324 7336
rect 21272 7293 21281 7327
rect 21281 7293 21315 7327
rect 21315 7293 21324 7327
rect 21272 7284 21324 7293
rect 16488 7148 16540 7200
rect 18420 7148 18472 7200
rect 19984 7216 20036 7268
rect 21180 7216 21232 7268
rect 24676 7327 24728 7336
rect 24676 7293 24720 7327
rect 24720 7293 24728 7327
rect 24676 7284 24728 7293
rect 23480 7148 23532 7200
rect 24768 7148 24820 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2228 6944 2280 6996
rect 5080 6944 5132 6996
rect 6460 6987 6512 6996
rect 6460 6953 6469 6987
rect 6469 6953 6503 6987
rect 6503 6953 6512 6987
rect 6460 6944 6512 6953
rect 8576 6944 8628 6996
rect 8760 6944 8812 6996
rect 17408 6944 17460 6996
rect 18328 6944 18380 6996
rect 19248 6944 19300 6996
rect 19984 6944 20036 6996
rect 20996 6944 21048 6996
rect 21180 6944 21232 6996
rect 1676 6876 1728 6928
rect 7104 6919 7156 6928
rect 7104 6885 7113 6919
rect 7113 6885 7147 6919
rect 7147 6885 7156 6919
rect 7104 6876 7156 6885
rect 2688 6808 2740 6860
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4344 6808 4396 6860
rect 6276 6808 6328 6860
rect 9680 6851 9732 6860
rect 2504 6740 2556 6792
rect 4896 6740 4948 6792
rect 7380 6783 7432 6792
rect 2228 6715 2280 6724
rect 2228 6681 2237 6715
rect 2237 6681 2271 6715
rect 2271 6681 2280 6715
rect 2228 6672 2280 6681
rect 3976 6672 4028 6724
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 7288 6672 7340 6724
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 10968 6808 11020 6860
rect 11060 6808 11112 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12624 6808 12676 6860
rect 13452 6808 13504 6860
rect 14832 6876 14884 6928
rect 12440 6740 12492 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 15476 6808 15528 6860
rect 18420 6876 18472 6928
rect 19064 6876 19116 6928
rect 21088 6919 21140 6928
rect 21088 6885 21097 6919
rect 21097 6885 21131 6919
rect 21131 6885 21140 6919
rect 21088 6876 21140 6885
rect 12808 6740 12860 6749
rect 13728 6740 13780 6792
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 16212 6808 16264 6860
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 22560 6851 22612 6860
rect 22560 6817 22569 6851
rect 22569 6817 22603 6851
rect 22603 6817 22612 6851
rect 22560 6808 22612 6817
rect 23940 6808 23992 6860
rect 25504 6808 25556 6860
rect 16396 6740 16448 6792
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 20996 6783 21048 6792
rect 2964 6604 3016 6656
rect 8760 6672 8812 6724
rect 15844 6672 15896 6724
rect 20996 6749 21005 6783
rect 21005 6749 21039 6783
rect 21039 6749 21048 6783
rect 20996 6740 21048 6749
rect 20720 6672 20772 6724
rect 22100 6740 22152 6792
rect 8576 6604 8628 6656
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 12440 6604 12492 6656
rect 13636 6604 13688 6656
rect 14004 6604 14056 6656
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 14832 6604 14884 6656
rect 17408 6604 17460 6656
rect 18052 6604 18104 6656
rect 19892 6647 19944 6656
rect 19892 6613 19901 6647
rect 19901 6613 19935 6647
rect 19935 6613 19944 6647
rect 19892 6604 19944 6613
rect 21272 6604 21324 6656
rect 23848 6604 23900 6656
rect 25136 6604 25188 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 5080 6400 5132 6452
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 10232 6400 10284 6452
rect 11888 6400 11940 6452
rect 12440 6400 12492 6452
rect 2688 6332 2740 6384
rect 5908 6375 5960 6384
rect 5908 6341 5917 6375
rect 5917 6341 5951 6375
rect 5951 6341 5960 6375
rect 5908 6332 5960 6341
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 3608 6264 3660 6316
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 4712 6196 4764 6248
rect 7656 6264 7708 6316
rect 8760 6196 8812 6248
rect 10784 6332 10836 6384
rect 11612 6332 11664 6384
rect 11796 6332 11848 6384
rect 17776 6400 17828 6452
rect 18512 6443 18564 6452
rect 18512 6409 18521 6443
rect 18521 6409 18555 6443
rect 18555 6409 18564 6443
rect 18512 6400 18564 6409
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 19248 6400 19300 6452
rect 21088 6400 21140 6452
rect 12440 6264 12492 6316
rect 14004 6332 14056 6384
rect 14464 6332 14516 6384
rect 14832 6332 14884 6384
rect 17224 6332 17276 6384
rect 18328 6375 18380 6384
rect 18328 6341 18337 6375
rect 18337 6341 18371 6375
rect 18371 6341 18380 6375
rect 18328 6332 18380 6341
rect 22192 6400 22244 6452
rect 22560 6400 22612 6452
rect 23940 6400 23992 6452
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 13728 6264 13780 6316
rect 15660 6264 15712 6316
rect 16212 6264 16264 6316
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 2228 6171 2280 6180
rect 1492 6060 1544 6112
rect 2228 6137 2237 6171
rect 2237 6137 2271 6171
rect 2271 6137 2280 6171
rect 2228 6128 2280 6137
rect 5080 6128 5132 6180
rect 6276 6171 6328 6180
rect 6276 6137 6285 6171
rect 6285 6137 6319 6171
rect 6319 6137 6328 6171
rect 6276 6128 6328 6137
rect 7196 6128 7248 6180
rect 2044 6060 2096 6112
rect 2320 6060 2372 6112
rect 2504 6060 2556 6112
rect 3792 6060 3844 6112
rect 4344 6060 4396 6112
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8760 6060 8812 6112
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 13636 6196 13688 6248
rect 12532 6128 12584 6180
rect 13452 6128 13504 6180
rect 14832 6128 14884 6180
rect 18144 6196 18196 6248
rect 21640 6332 21692 6384
rect 23480 6332 23532 6384
rect 24860 6375 24912 6384
rect 24860 6341 24869 6375
rect 24869 6341 24903 6375
rect 24903 6341 24912 6375
rect 24860 6332 24912 6341
rect 19892 6264 19944 6316
rect 21548 6307 21600 6316
rect 21548 6273 21557 6307
rect 21557 6273 21591 6307
rect 21591 6273 21600 6307
rect 21548 6264 21600 6273
rect 19248 6196 19300 6248
rect 19524 6196 19576 6248
rect 20076 6239 20128 6248
rect 20076 6205 20085 6239
rect 20085 6205 20119 6239
rect 20119 6205 20128 6239
rect 20076 6196 20128 6205
rect 20720 6196 20772 6248
rect 21272 6196 21324 6248
rect 24676 6239 24728 6248
rect 24676 6205 24685 6239
rect 24685 6205 24719 6239
rect 24719 6205 24728 6239
rect 24676 6196 24728 6205
rect 16580 6171 16632 6180
rect 16580 6137 16589 6171
rect 16589 6137 16623 6171
rect 16623 6137 16632 6171
rect 16580 6128 16632 6137
rect 17132 6171 17184 6180
rect 17132 6137 17141 6171
rect 17141 6137 17175 6171
rect 17175 6137 17184 6171
rect 17132 6128 17184 6137
rect 18052 6171 18104 6180
rect 18052 6137 18061 6171
rect 18061 6137 18095 6171
rect 18095 6137 18104 6171
rect 18052 6128 18104 6137
rect 9220 6060 9272 6112
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10692 6060 10744 6069
rect 11428 6060 11480 6112
rect 12072 6060 12124 6112
rect 13728 6103 13780 6112
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 13728 6060 13780 6069
rect 14924 6060 14976 6112
rect 17408 6060 17460 6112
rect 17960 6060 18012 6112
rect 18604 6060 18656 6112
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 23664 6103 23716 6112
rect 23664 6069 23673 6103
rect 23673 6069 23707 6103
rect 23707 6069 23716 6103
rect 23664 6060 23716 6069
rect 25504 6103 25556 6112
rect 25504 6069 25513 6103
rect 25513 6069 25547 6103
rect 25547 6069 25556 6103
rect 25504 6060 25556 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1492 5856 1544 5908
rect 1676 5856 1728 5908
rect 3976 5856 4028 5908
rect 4068 5856 4120 5908
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 1216 5788 1268 5840
rect 2688 5788 2740 5840
rect 7104 5899 7156 5908
rect 7104 5865 7113 5899
rect 7113 5865 7147 5899
rect 7147 5865 7156 5899
rect 7104 5856 7156 5865
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 8024 5856 8076 5908
rect 12532 5899 12584 5908
rect 12532 5865 12541 5899
rect 12541 5865 12575 5899
rect 12575 5865 12584 5899
rect 12532 5856 12584 5865
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 14924 5856 14976 5908
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 16580 5856 16632 5908
rect 17868 5856 17920 5908
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 18512 5856 18564 5908
rect 20076 5856 20128 5908
rect 20904 5856 20956 5908
rect 22192 5856 22244 5908
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 5080 5788 5132 5840
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 6552 5720 6604 5772
rect 7012 5788 7064 5840
rect 9864 5831 9916 5840
rect 2228 5652 2280 5704
rect 2780 5652 2832 5704
rect 4344 5652 4396 5704
rect 8024 5720 8076 5772
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 11152 5788 11204 5840
rect 12072 5788 12124 5840
rect 16488 5831 16540 5840
rect 9404 5720 9456 5772
rect 9588 5720 9640 5772
rect 2320 5584 2372 5636
rect 7656 5584 7708 5636
rect 6644 5516 6696 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 9680 5584 9732 5636
rect 11244 5652 11296 5704
rect 12440 5720 12492 5772
rect 16488 5797 16491 5831
rect 16491 5797 16525 5831
rect 16525 5797 16540 5831
rect 16488 5788 16540 5797
rect 17408 5831 17460 5840
rect 17408 5797 17417 5831
rect 17417 5797 17451 5831
rect 17451 5797 17460 5831
rect 17408 5788 17460 5797
rect 19064 5788 19116 5840
rect 12992 5720 13044 5772
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 20628 5720 20680 5772
rect 21824 5720 21876 5772
rect 22100 5720 22152 5772
rect 22376 5720 22428 5772
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 24032 5763 24084 5772
rect 24032 5729 24041 5763
rect 24041 5729 24075 5763
rect 24075 5729 24084 5763
rect 24032 5720 24084 5729
rect 25136 5763 25188 5772
rect 25136 5729 25145 5763
rect 25145 5729 25179 5763
rect 25179 5729 25188 5763
rect 25136 5720 25188 5729
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 12900 5652 12952 5704
rect 13728 5652 13780 5704
rect 16856 5652 16908 5704
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 18420 5652 18472 5704
rect 10968 5584 11020 5636
rect 12808 5584 12860 5636
rect 25320 5627 25372 5636
rect 25320 5593 25329 5627
rect 25329 5593 25363 5627
rect 25363 5593 25372 5627
rect 25320 5584 25372 5593
rect 10140 5516 10192 5568
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 12440 5516 12492 5568
rect 13452 5516 13504 5568
rect 14464 5516 14516 5568
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 19984 5559 20036 5568
rect 19984 5525 19993 5559
rect 19993 5525 20027 5559
rect 20027 5525 20036 5559
rect 19984 5516 20036 5525
rect 24216 5559 24268 5568
rect 24216 5525 24225 5559
rect 24225 5525 24259 5559
rect 24259 5525 24268 5559
rect 24216 5516 24268 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2688 5312 2740 5364
rect 5080 5312 5132 5364
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 7196 5312 7248 5364
rect 8024 5312 8076 5364
rect 9404 5312 9456 5364
rect 10232 5312 10284 5364
rect 11612 5312 11664 5364
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 14740 5312 14792 5364
rect 16120 5312 16172 5364
rect 16488 5312 16540 5364
rect 19064 5312 19116 5364
rect 19524 5312 19576 5364
rect 20628 5312 20680 5364
rect 22100 5355 22152 5364
rect 22100 5321 22109 5355
rect 22109 5321 22143 5355
rect 22143 5321 22152 5355
rect 22100 5312 22152 5321
rect 22928 5312 22980 5364
rect 24032 5312 24084 5364
rect 25136 5355 25188 5364
rect 25136 5321 25145 5355
rect 25145 5321 25179 5355
rect 25179 5321 25188 5355
rect 25136 5312 25188 5321
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3700 5176 3752 5228
rect 7472 5176 7524 5228
rect 1952 5083 2004 5092
rect 1952 5049 1961 5083
rect 1961 5049 1995 5083
rect 1995 5049 2004 5083
rect 1952 5040 2004 5049
rect 3700 5040 3752 5092
rect 5540 5108 5592 5160
rect 5264 5040 5316 5092
rect 7656 5040 7708 5092
rect 11152 5244 11204 5296
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 11244 5176 11296 5228
rect 8760 5108 8812 5160
rect 11060 5108 11112 5160
rect 13176 5244 13228 5296
rect 18880 5287 18932 5296
rect 18880 5253 18889 5287
rect 18889 5253 18923 5287
rect 18923 5253 18932 5287
rect 18880 5244 18932 5253
rect 16028 5176 16080 5228
rect 16764 5176 16816 5228
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 19984 5176 20036 5228
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 22376 5244 22428 5296
rect 26700 5244 26752 5296
rect 21916 5176 21968 5228
rect 12808 5108 12860 5160
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 8300 5040 8352 5092
rect 9588 5040 9640 5092
rect 9864 5040 9916 5092
rect 10784 5040 10836 5092
rect 13176 5083 13228 5092
rect 13176 5049 13185 5083
rect 13185 5049 13219 5083
rect 13219 5049 13228 5083
rect 13176 5040 13228 5049
rect 14832 5108 14884 5160
rect 14740 5083 14792 5092
rect 14740 5049 14749 5083
rect 14749 5049 14783 5083
rect 14783 5049 14792 5083
rect 14740 5040 14792 5049
rect 16580 5083 16632 5092
rect 16580 5049 16589 5083
rect 16589 5049 16623 5083
rect 16623 5049 16632 5083
rect 16580 5040 16632 5049
rect 19248 5040 19300 5092
rect 19984 5040 20036 5092
rect 23664 5083 23716 5092
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 9312 4972 9364 5024
rect 11980 4972 12032 5024
rect 12900 4972 12952 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 20904 5015 20956 5024
rect 20904 4981 20913 5015
rect 20913 4981 20947 5015
rect 20947 4981 20956 5015
rect 23664 5049 23673 5083
rect 23673 5049 23707 5083
rect 23707 5049 23716 5083
rect 23664 5040 23716 5049
rect 20904 4972 20956 4981
rect 21916 4972 21968 5024
rect 24124 5108 24176 5160
rect 23848 4972 23900 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 2780 4768 2832 4820
rect 3700 4811 3752 4820
rect 3700 4777 3709 4811
rect 3709 4777 3743 4811
rect 3743 4777 3752 4811
rect 3700 4768 3752 4777
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 5540 4768 5592 4820
rect 9312 4811 9364 4820
rect 9312 4777 9321 4811
rect 9321 4777 9355 4811
rect 9355 4777 9364 4811
rect 9312 4768 9364 4777
rect 10140 4768 10192 4820
rect 11520 4768 11572 4820
rect 2412 4743 2464 4752
rect 2412 4709 2421 4743
rect 2421 4709 2455 4743
rect 2455 4709 2464 4743
rect 2412 4700 2464 4709
rect 6276 4700 6328 4752
rect 6736 4700 6788 4752
rect 7932 4743 7984 4752
rect 7932 4709 7941 4743
rect 7941 4709 7975 4743
rect 7975 4709 7984 4743
rect 7932 4700 7984 4709
rect 10784 4700 10836 4752
rect 11152 4700 11204 4752
rect 12072 4700 12124 4752
rect 13452 4768 13504 4820
rect 14188 4768 14240 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 16764 4811 16816 4820
rect 16764 4777 16773 4811
rect 16773 4777 16807 4811
rect 16807 4777 16816 4811
rect 16764 4768 16816 4777
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 17500 4700 17552 4752
rect 19064 4700 19116 4752
rect 20996 4768 21048 4820
rect 21640 4700 21692 4752
rect 4344 4632 4396 4684
rect 5264 4632 5316 4684
rect 10140 4632 10192 4684
rect 10692 4632 10744 4684
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 15844 4675 15896 4684
rect 15844 4641 15853 4675
rect 15853 4641 15887 4675
rect 15887 4641 15896 4675
rect 15844 4632 15896 4641
rect 18880 4675 18932 4684
rect 18880 4641 18889 4675
rect 18889 4641 18923 4675
rect 18923 4641 18932 4675
rect 18880 4632 18932 4641
rect 24676 4675 24728 4684
rect 24676 4641 24685 4675
rect 24685 4641 24719 4675
rect 24719 4641 24728 4675
rect 24676 4632 24728 4641
rect 2504 4564 2556 4616
rect 3056 4564 3108 4616
rect 6368 4564 6420 4616
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 8760 4564 8812 4616
rect 11980 4564 12032 4616
rect 12532 4564 12584 4616
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 17224 4564 17276 4616
rect 17684 4564 17736 4616
rect 20812 4564 20864 4616
rect 21732 4564 21784 4616
rect 22192 4564 22244 4616
rect 10048 4496 10100 4548
rect 10692 4496 10744 4548
rect 10968 4539 11020 4548
rect 10968 4505 10977 4539
rect 10977 4505 11011 4539
rect 11011 4505 11020 4539
rect 10968 4496 11020 4505
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 7656 4471 7708 4480
rect 7656 4437 7665 4471
rect 7665 4437 7699 4471
rect 7699 4437 7708 4471
rect 7656 4428 7708 4437
rect 11244 4428 11296 4480
rect 11888 4428 11940 4480
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 12992 4428 13044 4480
rect 14832 4471 14884 4480
rect 14832 4437 14841 4471
rect 14841 4437 14875 4471
rect 14875 4437 14884 4471
rect 14832 4428 14884 4437
rect 24124 4428 24176 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2412 4224 2464 4276
rect 3884 4267 3936 4276
rect 3884 4233 3893 4267
rect 3893 4233 3927 4267
rect 3927 4233 3936 4267
rect 3884 4224 3936 4233
rect 4344 4267 4396 4276
rect 4344 4233 4353 4267
rect 4353 4233 4387 4267
rect 4387 4233 4396 4267
rect 4344 4224 4396 4233
rect 5080 4224 5132 4276
rect 6276 4267 6328 4276
rect 6276 4233 6285 4267
rect 6285 4233 6319 4267
rect 6319 4233 6328 4267
rect 6276 4224 6328 4233
rect 6368 4224 6420 4276
rect 7196 4224 7248 4276
rect 2596 4088 2648 4140
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 12072 4224 12124 4276
rect 19064 4267 19116 4276
rect 19064 4233 19073 4267
rect 19073 4233 19107 4267
rect 19107 4233 19116 4267
rect 19064 4224 19116 4233
rect 21640 4267 21692 4276
rect 21640 4233 21649 4267
rect 21649 4233 21683 4267
rect 21683 4233 21692 4267
rect 21640 4224 21692 4233
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 2596 3952 2648 4004
rect 5080 3952 5132 4004
rect 14832 4156 14884 4208
rect 9036 4131 9088 4140
rect 9036 4097 9045 4131
rect 9045 4097 9079 4131
rect 9079 4097 9088 4131
rect 9036 4088 9088 4097
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 16396 4156 16448 4208
rect 18880 4156 18932 4208
rect 19984 4156 20036 4208
rect 10784 4020 10836 4072
rect 11152 4063 11204 4072
rect 11152 4029 11170 4063
rect 11170 4029 11204 4063
rect 11152 4020 11204 4029
rect 14648 4020 14700 4072
rect 14924 4020 14976 4072
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 20996 4088 21048 4140
rect 21732 4088 21784 4140
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 9404 3995 9456 4004
rect 9404 3961 9413 3995
rect 9413 3961 9447 3995
rect 9447 3961 9456 3995
rect 9404 3952 9456 3961
rect 13176 3952 13228 4004
rect 13452 3952 13504 4004
rect 15752 3952 15804 4004
rect 18328 4020 18380 4072
rect 17684 3952 17736 4004
rect 20720 3995 20772 4004
rect 20720 3961 20729 3995
rect 20729 3961 20763 3995
rect 20763 3961 20772 3995
rect 20720 3952 20772 3961
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 8668 3927 8720 3936
rect 8668 3893 8677 3927
rect 8677 3893 8711 3927
rect 8711 3893 8720 3927
rect 8668 3884 8720 3893
rect 11336 3884 11388 3936
rect 14004 3884 14056 3936
rect 14832 3884 14884 3936
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 17500 3927 17552 3936
rect 17500 3893 17509 3927
rect 17509 3893 17543 3927
rect 17543 3893 17552 3927
rect 17500 3884 17552 3893
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 19984 3884 20036 3936
rect 22008 3952 22060 4004
rect 23940 4020 23992 4072
rect 24768 4020 24820 4072
rect 23664 3952 23716 4004
rect 22652 3884 22704 3936
rect 23480 3927 23532 3936
rect 23480 3893 23489 3927
rect 23489 3893 23523 3927
rect 23523 3893 23532 3927
rect 23480 3884 23532 3893
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 25136 3884 25188 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2412 3680 2464 3732
rect 5264 3680 5316 3732
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 7564 3680 7616 3732
rect 8116 3680 8168 3732
rect 8852 3680 8904 3732
rect 10140 3723 10192 3732
rect 2504 3655 2556 3664
rect 2504 3621 2513 3655
rect 2513 3621 2547 3655
rect 2547 3621 2556 3655
rect 2504 3612 2556 3621
rect 3240 3612 3292 3664
rect 5080 3612 5132 3664
rect 6644 3655 6696 3664
rect 6644 3621 6653 3655
rect 6653 3621 6687 3655
rect 6687 3621 6696 3655
rect 6644 3612 6696 3621
rect 6736 3655 6788 3664
rect 6736 3621 6745 3655
rect 6745 3621 6779 3655
rect 6779 3621 6788 3655
rect 6736 3612 6788 3621
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 10784 3680 10836 3732
rect 11980 3723 12032 3732
rect 10508 3655 10560 3664
rect 10508 3621 10517 3655
rect 10517 3621 10551 3655
rect 10551 3621 10560 3655
rect 10508 3612 10560 3621
rect 11980 3689 11989 3723
rect 11989 3689 12023 3723
rect 12023 3689 12032 3723
rect 11980 3680 12032 3689
rect 12624 3680 12676 3732
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 11520 3612 11572 3664
rect 2320 3544 2372 3596
rect 4712 3544 4764 3596
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 8760 3544 8812 3596
rect 10876 3544 10928 3596
rect 13544 3680 13596 3732
rect 13820 3680 13872 3732
rect 15384 3680 15436 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 17684 3723 17736 3732
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 14924 3655 14976 3664
rect 14924 3621 14933 3655
rect 14933 3621 14967 3655
rect 14967 3621 14976 3655
rect 14924 3612 14976 3621
rect 16488 3612 16540 3664
rect 18328 3612 18380 3664
rect 13820 3544 13872 3596
rect 19524 3680 19576 3732
rect 20076 3680 20128 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 21916 3680 21968 3732
rect 24032 3680 24084 3732
rect 19064 3612 19116 3664
rect 20904 3655 20956 3664
rect 20904 3621 20913 3655
rect 20913 3621 20947 3655
rect 20947 3621 20956 3655
rect 20904 3612 20956 3621
rect 20996 3587 21048 3596
rect 20996 3553 21005 3587
rect 21005 3553 21039 3587
rect 21039 3553 21048 3587
rect 20996 3544 21048 3553
rect 22560 3587 22612 3596
rect 22560 3553 22569 3587
rect 22569 3553 22603 3587
rect 22603 3553 22612 3587
rect 22560 3544 22612 3553
rect 24032 3544 24084 3596
rect 388 3476 440 3528
rect 1308 3476 1360 3528
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 7932 3476 7984 3528
rect 8668 3476 8720 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 6184 3408 6236 3460
rect 11704 3451 11756 3460
rect 11704 3417 11713 3451
rect 11713 3417 11747 3451
rect 11747 3417 11756 3451
rect 11704 3408 11756 3417
rect 2136 3340 2188 3392
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 16672 3383 16724 3392
rect 16672 3349 16681 3383
rect 16681 3349 16715 3383
rect 16715 3349 16724 3383
rect 16672 3340 16724 3349
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 3424 3136 3476 3188
rect 4712 3136 4764 3188
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 10876 3136 10928 3188
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12532 3136 12584 3188
rect 14740 3136 14792 3188
rect 5080 3068 5132 3120
rect 11060 3111 11112 3120
rect 11060 3077 11069 3111
rect 11069 3077 11103 3111
rect 11103 3077 11112 3111
rect 11060 3068 11112 3077
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 8576 3000 8628 3052
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 15752 3136 15804 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 19524 3179 19576 3188
rect 19524 3145 19533 3179
rect 19533 3145 19567 3179
rect 19567 3145 19576 3179
rect 19524 3136 19576 3145
rect 19984 3136 20036 3188
rect 22560 3179 22612 3188
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 6736 2932 6788 2984
rect 8208 2932 8260 2984
rect 12532 2932 12584 2984
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 14556 2932 14608 2984
rect 15384 2932 15436 2984
rect 2320 2907 2372 2916
rect 2320 2873 2329 2907
rect 2329 2873 2363 2907
rect 2363 2873 2372 2907
rect 2320 2864 2372 2873
rect 2412 2907 2464 2916
rect 2412 2873 2421 2907
rect 2421 2873 2455 2907
rect 2455 2873 2464 2907
rect 2412 2864 2464 2873
rect 3976 2907 4028 2916
rect 3976 2873 3985 2907
rect 3985 2873 4019 2907
rect 4019 2873 4028 2907
rect 3976 2864 4028 2873
rect 4528 2907 4580 2916
rect 4528 2873 4537 2907
rect 4537 2873 4571 2907
rect 4571 2873 4580 2907
rect 4528 2864 4580 2873
rect 8576 2907 8628 2916
rect 8576 2873 8585 2907
rect 8585 2873 8619 2907
rect 8619 2873 8628 2907
rect 8576 2864 8628 2873
rect 7104 2839 7156 2848
rect 7104 2805 7113 2839
rect 7113 2805 7147 2839
rect 7147 2805 7156 2839
rect 7104 2796 7156 2805
rect 11704 2864 11756 2916
rect 11520 2839 11572 2848
rect 11520 2805 11529 2839
rect 11529 2805 11563 2839
rect 11563 2805 11572 2839
rect 13820 2864 13872 2916
rect 16488 3068 16540 3120
rect 19616 3068 19668 3120
rect 15660 3000 15712 3052
rect 17316 3000 17368 3052
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 22560 3145 22569 3179
rect 22569 3145 22603 3179
rect 22603 3145 22612 3179
rect 22560 3136 22612 3145
rect 23572 3136 23624 3188
rect 24032 3136 24084 3188
rect 24216 3068 24268 3120
rect 16488 2864 16540 2916
rect 23572 2932 23624 2984
rect 25228 2975 25280 2984
rect 25228 2941 25237 2975
rect 25237 2941 25271 2975
rect 25271 2941 25280 2975
rect 25228 2932 25280 2941
rect 18236 2907 18288 2916
rect 18236 2873 18245 2907
rect 18245 2873 18279 2907
rect 18279 2873 18288 2907
rect 18236 2864 18288 2873
rect 21364 2907 21416 2916
rect 11520 2796 11572 2805
rect 19524 2796 19576 2848
rect 21364 2873 21373 2907
rect 21373 2873 21407 2907
rect 21407 2873 21416 2907
rect 21364 2864 21416 2873
rect 21456 2796 21508 2848
rect 23296 2864 23348 2916
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3516 2592 3568 2644
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 3332 2524 3384 2576
rect 4252 2567 4304 2576
rect 4252 2533 4261 2567
rect 4261 2533 4295 2567
rect 4295 2533 4304 2567
rect 4252 2524 4304 2533
rect 7104 2567 7156 2576
rect 7104 2533 7113 2567
rect 7113 2533 7147 2567
rect 7147 2533 7156 2567
rect 7104 2524 7156 2533
rect 1400 2499 1452 2508
rect 1400 2465 1444 2499
rect 1444 2465 1452 2499
rect 1400 2456 1452 2465
rect 6092 2456 6144 2508
rect 9220 2592 9272 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10508 2567 10560 2576
rect 10508 2533 10517 2567
rect 10517 2533 10551 2567
rect 10551 2533 10560 2567
rect 10508 2524 10560 2533
rect 11520 2524 11572 2576
rect 12256 2524 12308 2576
rect 13636 2592 13688 2644
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 13452 2567 13504 2576
rect 13452 2533 13461 2567
rect 13461 2533 13495 2567
rect 13495 2533 13504 2567
rect 13452 2524 13504 2533
rect 15200 2524 15252 2576
rect 16672 2567 16724 2576
rect 16672 2533 16681 2567
rect 16681 2533 16715 2567
rect 16715 2533 16724 2567
rect 16672 2524 16724 2533
rect 17224 2567 17276 2576
rect 17224 2533 17233 2567
rect 17233 2533 17267 2567
rect 17267 2533 17276 2567
rect 17224 2524 17276 2533
rect 18052 2524 18104 2576
rect 18512 2567 18564 2576
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 14096 2456 14148 2508
rect 15384 2456 15436 2508
rect 20444 2592 20496 2644
rect 20996 2635 21048 2644
rect 20996 2601 21005 2635
rect 21005 2601 21039 2635
rect 21039 2601 21048 2635
rect 20996 2592 21048 2601
rect 23388 2635 23440 2644
rect 23388 2601 23397 2635
rect 23397 2601 23431 2635
rect 23431 2601 23440 2635
rect 23388 2592 23440 2601
rect 20536 2456 20588 2508
rect 23848 2499 23900 2508
rect 23848 2465 23857 2499
rect 23857 2465 23891 2499
rect 23891 2465 23900 2499
rect 23848 2456 23900 2465
rect 2044 2388 2096 2440
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 7288 2431 7340 2440
rect 2688 2320 2740 2372
rect 6276 2363 6328 2372
rect 6276 2329 6285 2363
rect 6285 2329 6319 2363
rect 6319 2329 6328 2363
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 8576 2388 8628 2440
rect 11980 2431 12032 2440
rect 10968 2363 11020 2372
rect 6276 2320 6328 2329
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12164 2320 12216 2372
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 21180 2431 21232 2440
rect 21180 2397 21189 2431
rect 21189 2397 21223 2431
rect 21223 2397 21232 2431
rect 21180 2388 21232 2397
rect 24032 2431 24084 2440
rect 24032 2397 24041 2431
rect 24041 2397 24075 2431
rect 24075 2397 24084 2431
rect 24032 2388 24084 2397
rect 25596 2431 25648 2440
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 21088 2320 21140 2372
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 10508 2252 10560 2304
rect 13820 2252 13872 2304
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 20536 2295 20588 2304
rect 20536 2261 20545 2295
rect 20545 2261 20579 2295
rect 20579 2261 20588 2295
rect 20536 2252 20588 2261
rect 21916 2252 21968 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 6736 552 6788 604
rect 7012 552 7064 604
rect 11428 552 11480 604
rect 12348 552 12400 604
rect 14740 552 14792 604
rect 14832 552 14884 604
<< metal2 >>
rect 1950 27432 2006 27441
rect 1950 27367 2006 27376
rect 1490 26344 1546 26353
rect 1490 26279 1546 26288
rect 1398 25392 1454 25401
rect 1398 25327 1454 25336
rect 1412 23662 1440 25327
rect 1504 24274 1532 26279
rect 1582 24304 1638 24313
rect 1492 24268 1544 24274
rect 1582 24239 1638 24248
rect 1492 24210 1544 24216
rect 1504 23866 1532 24210
rect 1492 23860 1544 23866
rect 1492 23802 1544 23808
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1398 21992 1454 22001
rect 1398 21927 1454 21936
rect 1412 21010 1440 21927
rect 1504 21486 1532 23151
rect 1596 22574 1624 24239
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1584 22568 1636 22574
rect 1584 22510 1636 22516
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1490 21176 1546 21185
rect 1490 21111 1546 21120
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 20602 1440 20946
rect 1400 20596 1452 20602
rect 1400 20538 1452 20544
rect 1504 19922 1532 21111
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1504 19514 1532 19858
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1596 18306 1624 21286
rect 1676 20800 1728 20806
rect 1674 20768 1676 20777
rect 1728 20768 1730 20777
rect 1674 20703 1730 20712
rect 1412 18278 1624 18306
rect 1412 17898 1440 18278
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1412 17870 1532 17898
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1412 16998 1440 17682
rect 1400 16992 1452 16998
rect 1320 16940 1400 16946
rect 1320 16934 1452 16940
rect 1320 16918 1440 16934
rect 1216 15700 1268 15706
rect 1216 15642 1268 15648
rect 1124 14068 1176 14074
rect 1124 14010 1176 14016
rect 1136 13258 1164 14010
rect 1228 13326 1256 15642
rect 1216 13320 1268 13326
rect 1216 13262 1268 13268
rect 1124 13252 1176 13258
rect 1124 13194 1176 13200
rect 1228 12918 1256 13262
rect 1216 12912 1268 12918
rect 1216 12854 1268 12860
rect 1124 12708 1176 12714
rect 1124 12650 1176 12656
rect 1136 9110 1164 12650
rect 1216 12640 1268 12646
rect 1216 12582 1268 12588
rect 1228 10674 1256 12582
rect 1216 10668 1268 10674
rect 1216 10610 1268 10616
rect 1216 9580 1268 9586
rect 1216 9522 1268 9528
rect 1124 9104 1176 9110
rect 1124 9046 1176 9052
rect 1228 5846 1256 9522
rect 1216 5840 1268 5846
rect 1216 5782 1268 5788
rect 1320 3534 1348 16918
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14346 1440 14894
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1412 12646 1440 14282
rect 1504 14074 1532 17870
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1596 13977 1624 18158
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1688 15910 1716 16526
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1582 13968 1638 13977
rect 1492 13932 1544 13938
rect 1582 13903 1638 13912
rect 1492 13874 1544 13880
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 7274 1440 10610
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 1504 6118 1532 13874
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 13530 1624 13806
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1596 12186 1624 13466
rect 1688 12714 1716 15846
rect 1780 14385 1808 24006
rect 1860 23520 1912 23526
rect 1860 23462 1912 23468
rect 1872 15706 1900 23462
rect 1964 19378 1992 27367
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 2504 22432 2556 22438
rect 2504 22374 2556 22380
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2148 17134 2176 17478
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 17060 2096 17066
rect 2044 17002 2096 17008
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1872 14822 1900 15506
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 13841 1808 14214
rect 1766 13832 1822 13841
rect 1766 13767 1822 13776
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 12986 1808 13670
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1780 12714 1808 12922
rect 1676 12708 1728 12714
rect 1676 12650 1728 12656
rect 1768 12708 1820 12714
rect 1768 12650 1820 12656
rect 1780 12345 1808 12650
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1596 12158 1808 12186
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11801 1716 12038
rect 1674 11792 1730 11801
rect 1674 11727 1730 11736
rect 1688 11694 1716 11727
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1674 11520 1730 11529
rect 1596 9761 1624 11494
rect 1674 11455 1730 11464
rect 1688 11354 1716 11455
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1688 10810 1716 11154
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1780 10010 1808 12158
rect 1872 10146 1900 14758
rect 1964 10538 1992 16594
rect 2056 12374 2084 17002
rect 2148 15450 2176 17070
rect 2228 15904 2280 15910
rect 2226 15872 2228 15881
rect 2280 15872 2282 15881
rect 2226 15807 2282 15816
rect 2148 15422 2268 15450
rect 2136 15360 2188 15366
rect 2134 15328 2136 15337
rect 2188 15328 2190 15337
rect 2134 15263 2190 15272
rect 2240 14906 2268 15422
rect 2148 14878 2268 14906
rect 2148 13734 2176 14878
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 2134 13560 2190 13569
rect 2134 13495 2190 13504
rect 2148 13462 2176 13495
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2148 12986 2176 13398
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2134 12472 2190 12481
rect 2134 12407 2190 12416
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2056 11898 2084 12310
rect 2148 12238 2176 12407
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2148 11898 2176 12174
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2042 11248 2098 11257
rect 2042 11183 2044 11192
rect 2096 11183 2098 11192
rect 2044 11154 2096 11160
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1964 10266 1992 10474
rect 2056 10266 2084 11154
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1872 10118 2084 10146
rect 1688 9982 1808 10010
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1596 8022 1624 9590
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1596 7478 1624 7958
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1688 6934 1716 9982
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 6928 1728 6934
rect 1780 6905 1808 9862
rect 2056 9654 2084 10118
rect 2044 9648 2096 9654
rect 1950 9616 2006 9625
rect 2044 9590 2096 9596
rect 1950 9551 2006 9560
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8401 1900 8774
rect 1858 8392 1914 8401
rect 1858 8327 1914 8336
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1676 6870 1728 6876
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1582 6352 1638 6361
rect 1582 6287 1584 6296
rect 1636 6287 1638 6296
rect 1584 6258 1636 6264
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5914 1532 6054
rect 1492 5908 1544 5914
rect 1596 5896 1624 6258
rect 1676 5908 1728 5914
rect 1596 5868 1676 5896
rect 1492 5850 1544 5856
rect 1676 5850 1728 5856
rect 1872 5681 1900 7686
rect 1858 5672 1914 5681
rect 1858 5607 1914 5616
rect 1858 5264 1914 5273
rect 1858 5199 1860 5208
rect 1912 5199 1914 5208
rect 1860 5170 1912 5176
rect 1872 4826 1900 5170
rect 1964 5098 1992 9551
rect 2148 9450 2176 11018
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2056 9110 2084 9386
rect 2134 9344 2190 9353
rect 2134 9279 2190 9288
rect 2148 9178 2176 9279
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 2056 8838 2084 9046
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8090 2084 8774
rect 2148 8498 2176 9114
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2240 8022 2268 14758
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 9722 2360 13194
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2318 9616 2374 9625
rect 2318 9551 2374 9560
rect 2332 8634 2360 9551
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2332 8362 2360 8570
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2240 7546 2268 7958
rect 2424 7818 2452 17546
rect 2516 11354 2544 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 5538 20088 5594 20097
rect 10289 20080 10585 20100
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 5538 20023 5594 20032
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 19417 2636 19654
rect 2594 19408 2650 19417
rect 2594 19343 2650 19352
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 16153 2636 17478
rect 2976 16998 3004 17682
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 2594 16144 2650 16153
rect 2594 16079 2650 16088
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2516 10674 2544 11290
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2516 9450 2544 10474
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2502 9208 2558 9217
rect 2502 9143 2558 9152
rect 2516 9110 2544 9143
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2516 7478 2544 7822
rect 2504 7472 2556 7478
rect 2226 7440 2282 7449
rect 2504 7414 2556 7420
rect 2226 7375 2282 7384
rect 2240 7274 2268 7375
rect 2516 7290 2544 7414
rect 2228 7268 2280 7274
rect 2228 7210 2280 7216
rect 2332 7262 2544 7290
rect 2240 7002 2268 7210
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6186 2268 6666
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1860 3936 1912 3942
rect 1858 3904 1860 3913
rect 1912 3904 1914 3913
rect 1858 3839 1914 3848
rect 388 3528 440 3534
rect 388 3470 440 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 400 480 428 3470
rect 2056 3369 2084 6054
rect 2240 5710 2268 6122
rect 2332 6118 2360 7262
rect 2608 7154 2636 15846
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2700 12918 2728 14418
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2700 12374 2728 12854
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2792 10282 2820 14214
rect 2976 12889 3004 16934
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 14074 3096 14418
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3068 13977 3096 14010
rect 3148 14000 3200 14006
rect 3054 13968 3110 13977
rect 3148 13942 3200 13948
rect 3054 13903 3110 13912
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2962 12880 3018 12889
rect 3068 12850 3096 13126
rect 2962 12815 3018 12824
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11665 2912 12038
rect 3068 11762 3096 12786
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2870 11656 2926 11665
rect 2870 11591 2872 11600
rect 2924 11591 2926 11600
rect 2872 11562 2924 11568
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10470 2912 11154
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2700 10254 2820 10282
rect 2700 10198 2728 10254
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2778 10160 2834 10169
rect 2700 9722 2728 10134
rect 3160 10146 3188 13942
rect 2778 10095 2834 10104
rect 3068 10118 3188 10146
rect 2792 9994 2820 10095
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2700 8974 2728 9386
rect 2792 9194 2820 9930
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9722 2912 9862
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2792 9166 2912 9194
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8090 2728 8910
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 8022 2820 9046
rect 2884 8634 2912 9166
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2424 7126 2636 7154
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2332 5234 2360 5578
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2332 3602 2360 5170
rect 2424 4758 2452 7126
rect 2700 7018 2728 7754
rect 2608 6990 2728 7018
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6118 2544 6734
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2502 4720 2558 4729
rect 2424 4282 2452 4694
rect 2502 4655 2558 4664
rect 2516 4622 2544 4655
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2516 3890 2544 4558
rect 2608 4146 2636 6990
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6390 2728 6802
rect 2976 6662 3004 9318
rect 3068 7721 3096 10118
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3160 8974 3188 9998
rect 3252 9926 3280 16934
rect 3344 11150 3372 19314
rect 4066 19136 4122 19145
rect 4066 19071 4122 19080
rect 4080 17785 4108 19071
rect 5552 18834 5580 20023
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5552 18426 5580 18770
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3436 12102 3464 15846
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3528 11937 3556 17070
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3896 16114 3924 16662
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3698 14920 3754 14929
rect 3698 14855 3754 14864
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3514 11928 3570 11937
rect 3514 11863 3570 11872
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3528 10606 3556 11154
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10130 3464 10406
rect 3528 10266 3556 10542
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3252 7886 3280 9590
rect 3436 9518 3464 10066
rect 3528 10062 3556 10202
rect 3516 10056 3568 10062
rect 3514 10024 3516 10033
rect 3568 10024 3570 10033
rect 3514 9959 3570 9968
rect 3620 9625 3648 14758
rect 3712 13433 3740 14855
rect 3790 14104 3846 14113
rect 3790 14039 3792 14048
rect 3844 14039 3846 14048
rect 3792 14010 3844 14016
rect 3698 13424 3754 13433
rect 3698 13359 3754 13368
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3712 10985 3740 11494
rect 3790 11112 3846 11121
rect 3790 11047 3846 11056
rect 3698 10976 3754 10985
rect 3698 10911 3754 10920
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3054 7712 3110 7721
rect 3054 7647 3110 7656
rect 3344 7313 3372 8298
rect 3712 7478 3740 10746
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3330 7304 3386 7313
rect 3330 7239 3386 7248
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2688 6384 2740 6390
rect 2686 6352 2688 6361
rect 2740 6352 2742 6361
rect 2686 6287 2742 6296
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2700 5370 2728 5782
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2792 4826 2820 5646
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 4185 3096 4558
rect 3054 4176 3110 4185
rect 2596 4140 2648 4146
rect 3054 4111 3056 4120
rect 2596 4082 2648 4088
rect 3108 4111 3110 4120
rect 3056 4082 3108 4088
rect 2608 4010 2636 4082
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 2424 3862 2544 3890
rect 2424 3738 2452 3862
rect 2502 3768 2558 3777
rect 2412 3732 2464 3738
rect 2502 3703 2558 3712
rect 2412 3674 2464 3680
rect 2516 3670 2544 3703
rect 2504 3664 2556 3670
rect 2410 3632 2466 3641
rect 2320 3596 2372 3602
rect 2504 3606 2556 3612
rect 2410 3567 2466 3576
rect 2320 3538 2372 3544
rect 2136 3392 2188 3398
rect 2042 3360 2098 3369
rect 2136 3334 2188 3340
rect 2042 3295 2098 3304
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1122 1184 1178 1193
rect 1122 1119 1178 1128
rect 1136 480 1164 1119
rect 1412 513 1440 2450
rect 2056 2446 2084 3295
rect 2148 3097 2176 3334
rect 2134 3088 2190 3097
rect 2134 3023 2190 3032
rect 2424 2922 2452 3567
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2332 2689 2360 2858
rect 2318 2680 2374 2689
rect 2318 2615 2374 2624
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2686 2408 2742 2417
rect 2686 2343 2688 2352
rect 2740 2343 2742 2352
rect 2688 2314 2740 2320
rect 1950 2000 2006 2009
rect 1950 1935 2006 1944
rect 1398 504 1454 513
rect 386 0 442 480
rect 1122 0 1178 480
rect 1964 480 1992 1935
rect 3160 1306 3188 7142
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3252 3194 3280 3606
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3344 2582 3372 7239
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 2792 1278 3188 1306
rect 2792 480 2820 1278
rect 3436 1057 3464 3130
rect 3528 2650 3556 7346
rect 3804 6633 3832 11047
rect 3896 10849 3924 16050
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3974 13968 4030 13977
rect 3974 13903 4030 13912
rect 3882 10840 3938 10849
rect 3882 10775 3938 10784
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3896 9178 3924 9386
rect 3988 9217 4016 13903
rect 4080 10810 4108 14894
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4172 13530 4200 13738
rect 4264 13569 4292 15846
rect 4250 13560 4306 13569
rect 4160 13524 4212 13530
rect 4250 13495 4306 13504
rect 4160 13466 4212 13472
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12986 4200 13330
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11286 4292 11494
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4068 10668 4120 10674
rect 4172 10656 4200 11086
rect 4120 10628 4200 10656
rect 4068 10610 4120 10616
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 3974 9208 4030 9217
rect 3884 9172 3936 9178
rect 3974 9143 4030 9152
rect 3884 9114 3936 9120
rect 3974 8800 4030 8809
rect 3974 8735 4030 8744
rect 3988 6730 4016 8735
rect 4080 8498 4108 10474
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9382 4200 9998
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4172 8430 4200 9318
rect 4356 8480 4384 16594
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4540 14074 4568 15438
rect 4632 14822 4660 15506
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4540 13802 4568 14010
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4632 12714 4660 14758
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12850 4936 13126
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 10266 4844 10406
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4816 9586 4844 10202
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4264 8452 4384 8480
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4068 8084 4120 8090
rect 4172 8072 4200 8366
rect 4120 8044 4200 8072
rect 4068 8026 4120 8032
rect 4172 7857 4200 8044
rect 4158 7848 4214 7857
rect 4158 7783 4214 7792
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3790 6624 3846 6633
rect 3790 6559 3846 6568
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3620 2530 3648 6258
rect 3700 6248 3752 6254
rect 3976 6248 4028 6254
rect 3700 6190 3752 6196
rect 3974 6216 3976 6225
rect 4028 6216 4030 6225
rect 3712 5234 3740 6190
rect 3974 6151 4030 6160
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3712 4826 3740 5034
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3528 2502 3648 2530
rect 3422 1048 3478 1057
rect 3422 983 3478 992
rect 3528 480 3556 2502
rect 3804 1329 3832 6054
rect 3988 5914 4016 6151
rect 4080 5914 4108 6802
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4282 3924 4966
rect 4264 4729 4292 8452
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7410 4384 8298
rect 4908 7954 4936 10202
rect 5000 10169 5028 15846
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4986 10160 5042 10169
rect 5092 10130 5120 14758
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 13326 5212 14350
rect 5276 14278 5304 14894
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 14006 5304 14214
rect 5460 14074 5488 14418
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12714 5212 13262
rect 5460 12918 5488 13738
rect 5552 13462 5580 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 12986 5580 13398
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5184 11626 5212 12310
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5184 11286 5212 11562
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5184 10810 5212 11222
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5172 10600 5224 10606
rect 5170 10568 5172 10577
rect 5224 10568 5226 10577
rect 5170 10503 5226 10512
rect 5368 10248 5396 12786
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12442 5948 12582
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5538 12336 5594 12345
rect 5538 12271 5594 12280
rect 5552 11354 5580 12271
rect 6104 12238 6132 14826
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6104 11898 6132 12174
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 5724 11688 5776 11694
rect 5722 11656 5724 11665
rect 5776 11656 5778 11665
rect 5722 11591 5778 11600
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10810 5488 11086
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 6196 10418 6224 15438
rect 6104 10390 6224 10418
rect 5540 10260 5592 10266
rect 5368 10220 5540 10248
rect 5540 10202 5592 10208
rect 4986 10095 5042 10104
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5276 10010 5304 10066
rect 5276 9982 5580 10010
rect 5552 9654 5580 9982
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5092 9110 5120 9386
rect 5632 9376 5684 9382
rect 6104 9353 6132 10390
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6196 9382 6224 10066
rect 6184 9376 6236 9382
rect 5632 9318 5684 9324
rect 6090 9344 6146 9353
rect 5644 9217 5672 9318
rect 6184 9318 6236 9324
rect 6090 9279 6146 9288
rect 5630 9208 5686 9217
rect 5630 9143 5686 9152
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5092 8294 5120 9046
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 8362 5396 8570
rect 6012 8498 6040 8842
rect 5448 8492 5500 8498
rect 6000 8492 6052 8498
rect 5500 8452 5580 8480
rect 5448 8434 5500 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8022 5120 8230
rect 5552 8090 5580 8452
rect 6000 8434 6052 8440
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7546 4936 7890
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5092 7478 5120 7958
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5080 7472 5132 7478
rect 5552 7449 5580 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5080 7414 5132 7420
rect 5538 7440 5594 7449
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 5092 7274 5120 7414
rect 5538 7375 5594 7384
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5092 7002 5120 7210
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6118 4384 6802
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4526 6080 4582 6089
rect 4356 5710 4384 6054
rect 4526 6015 4582 6024
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4250 4720 4306 4729
rect 4356 4690 4384 5646
rect 4250 4655 4306 4664
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3974 2952 4030 2961
rect 3974 2887 3976 2896
rect 4028 2887 4030 2896
rect 3976 2858 4028 2864
rect 4080 2553 4108 4519
rect 4356 4282 4384 4626
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4252 3392 4304 3398
rect 4250 3360 4252 3369
rect 4304 3360 4306 3369
rect 4250 3295 4306 3304
rect 4540 2922 4568 6015
rect 4724 5914 4752 6190
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4908 5778 4936 6734
rect 5092 6458 5120 6938
rect 6196 6905 6224 9318
rect 6288 9058 6316 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 10138 18320 10194 18329
rect 10138 18255 10194 18264
rect 9494 16144 9550 16153
rect 9494 16079 9550 16088
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6366 13832 6422 13841
rect 6366 13767 6422 13776
rect 6380 11354 6408 13767
rect 7024 13462 7052 14010
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 13456 7064 13462
rect 6932 13404 7012 13410
rect 6932 13398 7064 13404
rect 6932 13382 7052 13398
rect 6932 12986 6960 13382
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7024 12918 7052 13262
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6918 11792 6974 11801
rect 7024 11762 7052 12310
rect 7116 12238 7144 13670
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7208 12442 7236 12922
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7300 11778 7328 13942
rect 7392 12481 7420 14350
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7484 13870 7512 14010
rect 7472 13864 7524 13870
rect 7470 13832 7472 13841
rect 7524 13832 7526 13841
rect 7470 13767 7526 13776
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7378 12472 7434 12481
rect 7378 12407 7434 12416
rect 7484 12322 7512 12786
rect 7760 12714 7788 12786
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7484 12294 7604 12322
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 6918 11727 6974 11736
rect 7012 11756 7064 11762
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6734 11112 6790 11121
rect 6734 11047 6736 11056
rect 6788 11047 6790 11056
rect 6736 11018 6788 11024
rect 6734 10976 6790 10985
rect 6734 10911 6790 10920
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6472 9722 6500 10406
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6288 9030 6408 9058
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 8634 6316 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 5170 6896 5226 6905
rect 5170 6831 5226 6840
rect 6182 6896 6238 6905
rect 6182 6831 6238 6840
rect 6276 6860 6328 6866
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5092 6186 5120 6394
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5846 5120 6122
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 5092 5370 5120 5782
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4724 3602 4752 4762
rect 5092 4282 5120 5306
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5092 4010 5120 4218
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 3670 5120 3946
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4724 3194 4752 3538
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5092 3126 5120 3606
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4342 2816 4398 2825
rect 4342 2751 4398 2760
rect 4252 2576 4304 2582
rect 3882 2544 3938 2553
rect 3882 2479 3938 2488
rect 4066 2544 4122 2553
rect 4252 2518 4304 2524
rect 4066 2479 4122 2488
rect 3896 1873 3924 2479
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3882 1864 3938 1873
rect 3882 1799 3938 1808
rect 4172 1601 4200 2382
rect 4264 1737 4292 2518
rect 4250 1728 4306 1737
rect 4250 1663 4306 1672
rect 4158 1592 4214 1601
rect 4158 1527 4214 1536
rect 3790 1320 3846 1329
rect 3790 1255 3846 1264
rect 4356 480 4384 2751
rect 4540 2446 4568 2858
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5184 480 5212 6831
rect 6276 6802 6328 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5908 6384 5960 6390
rect 5906 6352 5908 6361
rect 5960 6352 5962 6361
rect 5906 6287 5962 6296
rect 6288 6225 6316 6802
rect 6274 6216 6330 6225
rect 6274 6151 6276 6160
rect 6328 6151 6330 6160
rect 6276 6122 6328 6128
rect 5538 5808 5594 5817
rect 5538 5743 5594 5752
rect 5552 5166 5580 5743
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5276 4729 5304 5034
rect 5552 4826 5580 5102
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6276 4752 6328 4758
rect 5262 4720 5318 4729
rect 6276 4694 6328 4700
rect 5262 4655 5264 4664
rect 5316 4655 5318 4664
rect 5264 4626 5316 4632
rect 5276 3738 5304 4626
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6288 4282 6316 4694
rect 6380 4622 6408 9030
rect 6472 8945 6500 9658
rect 6458 8936 6514 8945
rect 6458 8871 6514 8880
rect 6458 8392 6514 8401
rect 6458 8327 6514 8336
rect 6472 7954 6500 8327
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6472 7002 6500 7890
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5370 6592 5714
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6380 4282 6408 4558
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 6090 3904 6146 3913
rect 5736 3777 5764 3878
rect 6090 3839 6146 3848
rect 5722 3768 5778 3777
rect 5264 3732 5316 3738
rect 6104 3738 6132 3839
rect 5722 3703 5778 3712
rect 6092 3732 6144 3738
rect 5264 3674 5316 3680
rect 6092 3674 6144 3680
rect 5538 3496 5594 3505
rect 5538 3431 5594 3440
rect 5998 3496 6054 3505
rect 5998 3431 6054 3440
rect 5552 3194 5580 3431
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5354 3088 5410 3097
rect 5354 3023 5410 3032
rect 5368 2990 5396 3023
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5368 2650 5396 2926
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5828 2553 5856 2586
rect 5814 2544 5870 2553
rect 5814 2479 5870 2488
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 1442 6040 3431
rect 6104 2514 6132 3674
rect 6656 3670 6684 5510
rect 6748 4758 6776 10911
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 8090 6868 10406
rect 6932 9654 6960 11727
rect 7300 11750 7420 11778
rect 7012 11698 7064 11704
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7208 11529 7236 11562
rect 7194 11520 7250 11529
rect 7194 11455 7250 11464
rect 7300 11218 7328 11562
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7392 10577 7420 11750
rect 7484 11354 7512 12174
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7576 11286 7604 12294
rect 7668 12084 7696 12650
rect 7840 12096 7892 12102
rect 7668 12056 7840 12084
rect 7840 12038 7892 12044
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7576 10810 7604 11222
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7378 10568 7434 10577
rect 7668 10538 7696 11698
rect 7378 10503 7434 10512
rect 7656 10532 7708 10538
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7116 9722 7144 10134
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7392 9654 7420 10503
rect 7656 10474 7708 10480
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7116 8362 7144 8978
rect 7392 8906 7420 9454
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 7116 6934 7144 8298
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7116 5914 7144 6870
rect 7208 6458 7236 8230
rect 7392 6798 7420 8842
rect 7668 8362 7696 10474
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7760 8090 7788 8434
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7208 6186 7236 6394
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7024 5030 7052 5782
rect 7208 5370 7236 6122
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6196 2961 6224 3402
rect 6748 2990 6776 3606
rect 6736 2984 6788 2990
rect 6182 2952 6238 2961
rect 6736 2926 6788 2932
rect 6182 2887 6238 2896
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6196 2145 6224 2887
rect 6274 2408 6330 2417
rect 6274 2343 6276 2352
rect 6328 2343 6330 2352
rect 6276 2314 6328 2320
rect 6182 2136 6238 2145
rect 6182 2071 6238 2080
rect 5920 1414 6040 1442
rect 5920 480 5948 1414
rect 7024 610 7052 4966
rect 7208 4282 7236 5306
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7300 3534 7328 6666
rect 7668 6322 7696 7142
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5234 7512 5510
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7668 5098 7696 5578
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7668 4486 7696 5034
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7668 4321 7696 4422
rect 7654 4312 7710 4321
rect 7654 4247 7710 4256
rect 7760 4146 7788 5850
rect 7852 5545 7880 12038
rect 7944 11762 7972 12786
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7944 9518 7972 10066
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7930 7984 7986 7993
rect 7930 7919 7932 7928
rect 7984 7919 7986 7928
rect 7932 7890 7984 7896
rect 7944 7342 7972 7890
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8036 5914 8064 14758
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8300 13864 8352 13870
rect 8128 13824 8300 13852
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7838 5536 7894 5545
rect 7838 5471 7894 5480
rect 8036 5370 8064 5714
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7852 4457 7880 4558
rect 7838 4448 7894 4457
rect 7838 4383 7894 4392
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2582 7144 2790
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7300 2446 7328 3470
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 6736 604 6788 610
rect 6736 546 6788 552
rect 7012 604 7064 610
rect 7012 546 7064 552
rect 6748 480 6776 546
rect 7576 480 7604 3674
rect 7944 3534 7972 4694
rect 8128 3738 8156 13824
rect 8300 13806 8352 13812
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8772 13530 8800 13738
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8680 13161 8708 13330
rect 8666 13152 8722 13161
rect 8666 13087 8722 13096
rect 8680 12918 8708 13087
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8680 12442 8708 12854
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8496 11150 8524 12174
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10606 8800 10950
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8772 10266 8800 10542
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8390 9616 8446 9625
rect 8390 9551 8446 9560
rect 8404 9518 8432 9551
rect 8588 9518 8616 9998
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8404 9178 8432 9454
rect 8680 9330 8708 9454
rect 8588 9302 8708 9330
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8220 7342 8248 7890
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8128 2650 8156 3538
rect 8220 2990 8248 6054
rect 8312 5098 8340 7822
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8312 1578 8340 3334
rect 8220 1550 8340 1578
rect 8220 1465 8248 1550
rect 8206 1456 8262 1465
rect 8404 1442 8432 8502
rect 8496 1601 8524 8910
rect 8588 7954 8616 9302
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7002 8616 7890
rect 8772 7460 8800 10066
rect 8680 7432 8800 7460
rect 8680 7342 8708 7432
rect 8772 7342 8800 7373
rect 8668 7336 8720 7342
rect 8760 7336 8812 7342
rect 8668 7278 8720 7284
rect 8758 7304 8760 7313
rect 8812 7304 8814 7313
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8680 6882 8708 7278
rect 8758 7239 8814 7248
rect 8772 7002 8800 7239
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8588 6854 8708 6882
rect 8588 6662 8616 6854
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8772 6254 8800 6666
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8760 6112 8812 6118
rect 8758 6080 8760 6089
rect 8812 6080 8814 6089
rect 8758 6015 8814 6024
rect 8760 5160 8812 5166
rect 8758 5128 8760 5137
rect 8812 5128 8814 5137
rect 8758 5063 8814 5072
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8680 3777 8708 3878
rect 8666 3768 8722 3777
rect 8666 3703 8722 3712
rect 8680 3534 8708 3703
rect 8772 3602 8800 4558
rect 8864 3738 8892 14214
rect 8956 13870 8984 14418
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8574 3360 8630 3369
rect 8574 3295 8630 3304
rect 8588 3058 8616 3295
rect 8772 3058 8800 3538
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8588 2446 8616 2858
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 1873 8708 2246
rect 8758 2136 8814 2145
rect 8758 2071 8814 2080
rect 8666 1864 8722 1873
rect 8666 1799 8722 1808
rect 8772 1601 8800 2071
rect 8482 1592 8538 1601
rect 8482 1527 8538 1536
rect 8758 1592 8814 1601
rect 8758 1527 8814 1536
rect 8206 1391 8262 1400
rect 8312 1414 8432 1442
rect 8312 480 8340 1414
rect 8482 1320 8538 1329
rect 8482 1255 8538 1264
rect 8496 1057 8524 1255
rect 8482 1048 8538 1057
rect 8482 983 8538 992
rect 8956 626 8984 13806
rect 9048 4146 9076 13874
rect 9140 8566 9168 14758
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9232 9926 9260 10542
rect 9324 10130 9352 12582
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11286 9444 11562
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9416 10810 9444 11222
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9722 9260 9862
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9232 8498 9260 8910
rect 9324 8634 9352 9386
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 7313 9168 8366
rect 9324 8022 9352 8570
rect 9416 8566 9444 8774
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9416 7546 9444 8502
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9126 7304 9182 7313
rect 9126 7239 9182 7248
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9140 3913 9168 7142
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9126 3904 9182 3913
rect 9126 3839 9182 3848
rect 9232 2650 9260 6054
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9416 5370 9444 5714
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4826 9352 4966
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9416 4010 9444 5306
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9508 2650 9536 16079
rect 10152 15570 10180 18255
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 11150 17776 11206 17785
rect 11150 17711 11152 17720
rect 11204 17711 11206 17720
rect 11152 17682 11204 17688
rect 11164 17338 11192 17682
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10152 15162 10180 15506
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 12782 9720 13330
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9784 12442 9812 13126
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 10985 9628 12174
rect 9586 10976 9642 10985
rect 9586 10911 9642 10920
rect 9586 10024 9642 10033
rect 9586 9959 9642 9968
rect 9600 9178 9628 9959
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8090 9628 8842
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9692 6866 9720 12378
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9784 11898 9812 12242
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9588 5772 9640 5778
rect 9784 5760 9812 11834
rect 9876 7818 9904 13806
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9640 5732 9812 5760
rect 9588 5714 9640 5720
rect 9770 5672 9826 5681
rect 9680 5636 9732 5642
rect 9770 5607 9826 5616
rect 9680 5578 9732 5584
rect 9692 5234 9720 5578
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9586 5128 9642 5137
rect 9586 5063 9588 5072
rect 9640 5063 9642 5072
rect 9588 5034 9640 5040
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9692 2145 9720 5170
rect 9784 2417 9812 5607
rect 9876 5098 9904 5782
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9862 4448 9918 4457
rect 9862 4383 9918 4392
rect 9876 4146 9904 4383
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9770 2408 9826 2417
rect 9770 2343 9826 2352
rect 9678 2136 9734 2145
rect 9678 2071 9734 2080
rect 8956 598 9168 626
rect 9140 480 9168 598
rect 9968 480 9996 14894
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10046 13832 10102 13841
rect 10046 13767 10102 13776
rect 10060 12646 10088 13767
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11354 10088 11698
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10060 8838 10088 11018
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 8022 10088 8774
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 4554 10088 7754
rect 10152 5681 10180 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10520 14074 10548 14418
rect 10704 14090 10732 15302
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10612 14062 10732 14090
rect 10876 14068 10928 14074
rect 10612 13716 10640 14062
rect 10876 14010 10928 14016
rect 10692 14000 10744 14006
rect 10690 13968 10692 13977
rect 10744 13968 10746 13977
rect 10690 13903 10746 13912
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10612 13688 10732 13716
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13410 10732 13688
rect 10796 13530 10824 13738
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10612 13382 10732 13410
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10232 12776 10284 12782
rect 10230 12744 10232 12753
rect 10284 12744 10286 12753
rect 10428 12714 10456 13126
rect 10612 12889 10640 13382
rect 10796 13240 10824 13466
rect 10704 13212 10824 13240
rect 10598 12880 10654 12889
rect 10704 12850 10732 13212
rect 10888 12918 10916 14010
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10876 12912 10928 12918
rect 10796 12872 10876 12900
rect 10598 12815 10654 12824
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10230 12679 10286 12688
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10796 12084 10824 12872
rect 10876 12854 10928 12860
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10888 12594 10916 12718
rect 11164 12714 11192 13262
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 10888 12566 11008 12594
rect 10874 12472 10930 12481
rect 10874 12407 10930 12416
rect 10888 12238 10916 12407
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10876 12096 10928 12102
rect 10796 12056 10876 12084
rect 10876 12038 10928 12044
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10416 11280 10468 11286
rect 10414 11248 10416 11257
rect 10468 11248 10470 11257
rect 10414 11183 10470 11192
rect 10704 10810 10732 11562
rect 10796 11286 10824 11698
rect 10888 11286 10916 12038
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10692 10192 10744 10198
rect 10506 10160 10562 10169
rect 10692 10134 10744 10140
rect 10506 10095 10562 10104
rect 10520 9489 10548 10095
rect 10506 9480 10562 9489
rect 10506 9415 10562 9424
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 8634 10272 9046
rect 10704 8974 10732 10134
rect 10796 9178 10824 10950
rect 10888 10810 10916 11086
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10980 10198 11008 12566
rect 11164 12458 11192 12650
rect 11164 12430 11227 12458
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10968 10192 11020 10198
rect 10874 10160 10930 10169
rect 10968 10134 11020 10140
rect 10874 10095 10876 10104
rect 10928 10095 10930 10104
rect 10876 10066 10928 10072
rect 10888 9722 10916 10066
rect 11072 10010 11100 12310
rect 11199 11778 11227 12430
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11164 11750 11227 11778
rect 11164 11014 11192 11750
rect 11348 11354 11376 12174
rect 11440 11830 11468 14214
rect 11532 13841 11560 14758
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11900 13870 11928 14418
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 13864 11940 13870
rect 11518 13832 11574 13841
rect 11888 13806 11940 13812
rect 11518 13767 11574 13776
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11532 12646 11560 12922
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11334 10704 11390 10713
rect 11334 10639 11390 10648
rect 10980 9982 11100 10010
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10980 9654 11008 9982
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10874 9480 10930 9489
rect 10874 9415 10930 9424
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10244 8362 10272 8570
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7818 10732 8502
rect 10796 8430 10824 9114
rect 10888 9110 10916 9415
rect 10980 9110 11008 9590
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11058 8936 11114 8945
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10784 8424 10836 8430
rect 10782 8392 10784 8401
rect 10836 8392 10838 8401
rect 10782 8327 10838 8336
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7954 10824 8230
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10796 7478 10824 7890
rect 10888 7818 10916 8502
rect 10980 8498 11008 8910
rect 11058 8871 11114 8880
rect 11072 8634 11100 8871
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 7886 11008 8434
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11058 7848 11114 7857
rect 10876 7812 10928 7818
rect 11058 7783 11060 7792
rect 10876 7754 10928 7760
rect 11112 7783 11114 7792
rect 11060 7754 11112 7760
rect 10888 7546 10916 7754
rect 11164 7562 11192 9046
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10980 7534 11192 7562
rect 10784 7472 10836 7478
rect 10980 7426 11008 7534
rect 10784 7414 10836 7420
rect 10888 7398 11008 7426
rect 11060 7472 11112 7478
rect 11112 7432 11192 7460
rect 11060 7414 11112 7420
rect 10888 7154 10916 7398
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10796 7126 10916 7154
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6769 10364 6802
rect 10322 6760 10378 6769
rect 10322 6695 10378 6704
rect 10232 6452 10284 6458
rect 10336 6440 10364 6695
rect 10284 6412 10364 6440
rect 10232 6394 10284 6400
rect 10796 6390 10824 7126
rect 10874 7032 10930 7041
rect 10874 6967 10930 6976
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10138 5672 10194 5681
rect 10138 5607 10194 5616
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10230 5536 10286 5545
rect 10152 4826 10180 5510
rect 10230 5471 10286 5480
rect 10244 5370 10272 5471
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10704 4690 10732 6054
rect 10796 5817 10824 6326
rect 10782 5808 10838 5817
rect 10782 5743 10838 5752
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10796 4865 10824 5034
rect 10782 4856 10838 4865
rect 10782 4791 10838 4800
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10152 3738 10180 4626
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10520 3058 10548 3606
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10520 2310 10548 2518
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10520 1737 10548 2246
rect 10506 1728 10562 1737
rect 10506 1663 10562 1672
rect 10704 480 10732 4490
rect 10796 4078 10824 4694
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10796 3738 10824 4014
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10888 3602 10916 6967
rect 10980 6866 11008 7210
rect 11072 7177 11100 7278
rect 11058 7168 11114 7177
rect 11058 7103 11114 7112
rect 11072 6866 11100 7103
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5642 11008 6190
rect 11164 5846 11192 7432
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11256 5710 11284 7686
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10966 4584 11022 4593
rect 10966 4519 10968 4528
rect 11020 4519 11022 4528
rect 10968 4490 11020 4496
rect 11072 4434 11100 5102
rect 11164 4758 11192 5238
rect 11256 5234 11284 5646
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11256 4486 11284 5170
rect 10980 4406 11100 4434
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10888 3194 10916 3538
rect 10980 3505 11008 4406
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11060 3120 11112 3126
rect 10966 3088 11022 3097
rect 11022 3068 11060 3074
rect 11022 3062 11112 3068
rect 11022 3046 11100 3062
rect 10966 3023 11022 3032
rect 10980 2378 11008 3023
rect 11164 2961 11192 4014
rect 11348 3942 11376 10639
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 9178 11468 9862
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11532 8906 11560 12582
rect 11612 12368 11664 12374
rect 11716 12356 11744 13126
rect 11808 12986 11836 13330
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11664 12328 11744 12356
rect 11612 12310 11664 12316
rect 11624 11898 11652 12310
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 9586 11744 11018
rect 11808 10810 11836 12922
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11900 10169 11928 13806
rect 11886 10160 11942 10169
rect 11808 10118 11886 10146
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 8548 11560 8842
rect 11440 8520 11560 8548
rect 11440 7410 11468 8520
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11532 6662 11560 8298
rect 11716 7886 11744 8978
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11440 610 11468 6054
rect 11532 5574 11560 6598
rect 11808 6390 11836 10118
rect 11886 10095 11942 10104
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11900 8090 11928 9046
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11900 6866 11928 7210
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11900 6458 11928 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11624 5710 11652 6326
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 4826 11560 5510
rect 11624 5370 11652 5646
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11716 4729 11744 5510
rect 11992 5030 12020 14214
rect 12070 12744 12126 12753
rect 12070 12679 12126 12688
rect 12084 6118 12112 12679
rect 12176 12238 12204 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 15474 16688 15530 16697
rect 15474 16623 15530 16632
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15488 15570 15516 16623
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15488 15162 15516 15506
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 13002 12388 14758
rect 15580 14482 15608 15943
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15580 14074 15608 14418
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12452 13161 12480 13806
rect 12438 13152 12494 13161
rect 12438 13087 12494 13096
rect 12360 12974 12480 13002
rect 12452 12356 12480 12974
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12268 12328 12480 12356
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12176 10742 12204 11222
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 10198 12204 10678
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12176 9722 12204 10134
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12084 5370 12112 5782
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11702 4720 11758 4729
rect 11702 4655 11758 4664
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11808 4457 11836 4626
rect 11992 4622 12020 4966
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11888 4480 11940 4486
rect 11794 4448 11850 4457
rect 11888 4422 11940 4428
rect 11794 4383 11850 4392
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 2854 11560 3606
rect 11702 3496 11758 3505
rect 11702 3431 11704 3440
rect 11756 3431 11758 3440
rect 11704 3402 11756 3408
rect 11716 2922 11744 3402
rect 11900 3194 11928 4422
rect 11992 3738 12020 4558
rect 12084 4486 12112 4694
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4282 12112 4422
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 12268 2582 12296 12328
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12360 10742 12388 12106
rect 12544 11694 12572 12378
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12452 10470 12480 10746
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 9625 12572 11630
rect 12636 11558 12664 11834
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12530 9616 12586 9625
rect 12530 9551 12586 9560
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8498 12480 8774
rect 12544 8514 12572 9551
rect 12636 9081 12664 11494
rect 12728 10266 12756 13942
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12820 11354 12848 12718
rect 12912 11762 12940 14010
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 12374 13216 12650
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13188 11898 13216 12310
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13372 11778 13400 13126
rect 13464 12986 13492 13262
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 12900 11756 12952 11762
rect 13280 11750 13400 11778
rect 12952 11716 13032 11744
rect 12900 11698 12952 11704
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12820 10810 12848 11290
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12728 9518 12756 10202
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12622 9072 12678 9081
rect 12622 9007 12678 9016
rect 12806 9072 12862 9081
rect 12806 9007 12862 9016
rect 12820 8566 12848 9007
rect 12912 8634 12940 11562
rect 13004 11354 13032 11716
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 8560 12860 8566
rect 12440 8492 12492 8498
rect 12544 8486 12664 8514
rect 12808 8502 12860 8508
rect 12440 8434 12492 8440
rect 12438 8392 12494 8401
rect 12494 8350 12572 8378
rect 12438 8327 12494 8336
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7993 12480 8230
rect 12438 7984 12494 7993
rect 12438 7919 12494 7928
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7546 12388 7754
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12452 6798 12480 7919
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6458 12480 6598
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12452 5817 12480 6258
rect 12544 6186 12572 8350
rect 12636 6866 12664 8486
rect 12820 7546 12848 8502
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 7410 12940 7890
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12806 6896 12862 6905
rect 12624 6860 12676 6866
rect 12806 6831 12862 6840
rect 12624 6802 12676 6808
rect 12820 6798 12848 6831
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12912 6225 12940 6258
rect 12898 6216 12954 6225
rect 12532 6180 12584 6186
rect 12898 6151 12954 6160
rect 12532 6122 12584 6128
rect 12544 5914 12572 6122
rect 12532 5908 12584 5914
rect 13004 5896 13032 11018
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13188 10538 13216 10678
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10305 13216 10474
rect 13174 10296 13230 10305
rect 13174 10231 13230 10240
rect 13280 10146 13308 11750
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13188 10118 13308 10146
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 9042 13124 9454
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13096 7732 13124 8978
rect 13188 8838 13216 10118
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13280 8634 13308 9454
rect 13372 9042 13400 11562
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13464 10146 13492 11290
rect 13556 10674 13584 12650
rect 13648 11354 13676 13806
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11898 13768 12174
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13820 11280 13872 11286
rect 13740 11240 13820 11268
rect 13740 10810 13768 11240
rect 13820 11222 13872 11228
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10266 13584 10610
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13464 10118 13676 10146
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13464 9110 13492 9998
rect 13648 9330 13676 10118
rect 13832 9994 13860 10542
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9586 13860 9930
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13726 9344 13782 9353
rect 13648 9302 13726 9330
rect 13726 9279 13782 9288
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8090 13400 8978
rect 13740 8974 13768 9279
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8634 13768 8910
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13450 7848 13506 7857
rect 13176 7744 13228 7750
rect 13096 7704 13176 7732
rect 13176 7686 13228 7692
rect 12584 5868 12664 5896
rect 13004 5868 13124 5896
rect 12532 5850 12584 5856
rect 12438 5808 12494 5817
rect 12438 5743 12440 5752
rect 12492 5743 12494 5752
rect 12440 5714 12492 5720
rect 12452 5574 12480 5714
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4321 12480 4422
rect 12438 4312 12494 4321
rect 12438 4247 12494 4256
rect 12544 3194 12572 4558
rect 12636 4457 12664 5868
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12820 5166 12848 5578
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12622 4448 12678 4457
rect 12622 4383 12678 4392
rect 12636 3738 12664 4383
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12728 4049 12756 4082
rect 12714 4040 12770 4049
rect 12714 3975 12770 3984
rect 12820 3738 12848 5102
rect 12912 5030 12940 5646
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 13004 4486 13032 5714
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12544 2990 12572 3130
rect 13004 3058 13032 4422
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 11428 604 11480 610
rect 11428 546 11480 552
rect 11532 480 11560 2518
rect 11980 2440 12032 2446
rect 11978 2408 11980 2417
rect 12032 2408 12034 2417
rect 11978 2343 12034 2352
rect 12162 2408 12218 2417
rect 12162 2343 12164 2352
rect 12216 2343 12218 2352
rect 12164 2314 12216 2320
rect 12348 604 12400 610
rect 12348 546 12400 552
rect 12360 480 12388 546
rect 13096 480 13124 5868
rect 13188 5302 13216 7686
rect 13266 5536 13322 5545
rect 13266 5471 13322 5480
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4729 13216 5034
rect 13174 4720 13230 4729
rect 13174 4655 13230 4664
rect 13176 4004 13228 4010
rect 13280 3992 13308 5471
rect 13228 3964 13308 3992
rect 13176 3946 13228 3952
rect 13266 3632 13322 3641
rect 13266 3567 13322 3576
rect 13280 2990 13308 3567
rect 13372 3369 13400 7822
rect 13450 7783 13506 7792
rect 13464 7546 13492 7783
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13464 6186 13492 6802
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 4826 13492 5510
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13358 3360 13414 3369
rect 13358 3295 13414 3304
rect 13268 2984 13320 2990
rect 13464 2961 13492 3946
rect 13556 3738 13584 8298
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13740 7274 13768 7375
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13832 7041 13860 7142
rect 13818 7032 13874 7041
rect 13818 6967 13874 6976
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6254 13676 6598
rect 13740 6322 13768 6734
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13740 6118 13768 6258
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5710 13768 6054
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13544 3732 13596 3738
rect 13820 3732 13872 3738
rect 13544 3674 13596 3680
rect 13648 3692 13820 3720
rect 13268 2926 13320 2932
rect 13450 2952 13506 2961
rect 13450 2887 13506 2896
rect 13464 2582 13492 2887
rect 13648 2650 13676 3692
rect 13820 3674 13872 3680
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13832 2922 13860 3538
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13832 2650 13860 2858
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13832 1465 13860 2246
rect 13818 1456 13874 1465
rect 13818 1391 13874 1400
rect 13924 480 13952 13806
rect 15382 13424 15438 13433
rect 14004 13388 14056 13394
rect 15382 13359 15384 13368
rect 14004 13330 14056 13336
rect 15436 13359 15438 13368
rect 15384 13330 15436 13336
rect 14016 13161 14044 13330
rect 14648 13184 14700 13190
rect 14002 13152 14058 13161
rect 14648 13126 14700 13132
rect 14002 13087 14058 13096
rect 14016 12986 14044 13087
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14016 11150 14044 12106
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14016 10198 14044 10406
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 14016 9722 14044 10134
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14016 8634 14044 9658
rect 14108 9489 14136 12718
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 12442 14228 12582
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14568 11082 14596 12786
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14188 9512 14240 9518
rect 14094 9480 14150 9489
rect 14188 9454 14240 9460
rect 14094 9415 14150 9424
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9110 14136 9318
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14200 8430 14228 9454
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 8430 14320 8774
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14200 7410 14228 8366
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 6390 14044 6598
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14200 5166 14228 7346
rect 14292 7342 14320 7686
rect 14660 7342 14688 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12986 15424 13330
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15396 11898 15424 12242
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14752 10266 14780 11086
rect 14844 10810 14872 11222
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14936 9178 14964 9454
rect 15304 9178 15332 10406
rect 15396 10198 15424 11834
rect 15764 10810 15792 12038
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15764 10470 15792 10746
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15750 10296 15806 10305
rect 15750 10231 15806 10240
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15396 9722 15424 10134
rect 15764 10062 15792 10231
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14936 8945 14964 9114
rect 14922 8936 14978 8945
rect 14922 8871 14978 8880
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14738 8528 14794 8537
rect 15580 8498 15608 9386
rect 15764 9178 15792 9998
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15948 8974 15976 14214
rect 16028 12776 16080 12782
rect 16026 12744 16028 12753
rect 16080 12744 16082 12753
rect 16026 12679 16082 12688
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 11914 16252 12582
rect 16040 11886 16252 11914
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 14738 8463 14794 8472
rect 15568 8492 15620 8498
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14292 6662 14320 7278
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4826 14228 5102
rect 14292 5001 14320 6598
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14476 5914 14504 6326
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14476 5574 14504 5850
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14278 4992 14334 5001
rect 14278 4927 14334 4936
rect 14554 4856 14610 4865
rect 14188 4820 14240 4826
rect 14554 4791 14610 4800
rect 14188 4762 14240 4768
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 3942 14044 4626
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14568 2990 14596 4791
rect 14660 4078 14688 7278
rect 14752 5817 14780 8463
rect 15568 8434 15620 8440
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14844 6934 14872 8366
rect 15580 8090 15608 8434
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 6928 14884 6934
rect 14832 6870 14884 6876
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6390 14872 6598
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 6384 14884 6390
rect 14830 6352 14832 6361
rect 14884 6352 14886 6361
rect 14830 6287 14886 6296
rect 14844 6261 14872 6287
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14738 5808 14794 5817
rect 14738 5743 14794 5752
rect 14752 5370 14780 5743
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14844 5166 14872 6122
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5914 14964 6054
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5273 15332 7822
rect 15764 7274 15792 8502
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15488 6089 15516 6802
rect 15660 6792 15712 6798
rect 15566 6760 15622 6769
rect 15660 6734 15712 6740
rect 15566 6695 15622 6704
rect 15474 6080 15530 6089
rect 15474 6015 15530 6024
rect 15488 5914 15516 6015
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15290 5264 15346 5273
rect 15290 5199 15346 5208
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14752 3194 14780 5034
rect 14844 4486 14872 5102
rect 15382 4584 15438 4593
rect 15382 4519 15384 4528
rect 15436 4519 15438 4528
rect 15384 4490 15436 4496
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4214 14872 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15382 4312 15438 4321
rect 15382 4247 15438 4256
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14108 2009 14136 2450
rect 14094 2000 14150 2009
rect 14094 1935 14150 1944
rect 14844 610 14872 3878
rect 14936 3670 14964 4014
rect 15396 3738 15424 4247
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15382 3224 15438 3233
rect 15382 3159 15438 3168
rect 15396 2990 15424 3159
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15200 2576 15252 2582
rect 15198 2544 15200 2553
rect 15252 2544 15254 2553
rect 15198 2479 15254 2488
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 2009 15332 2246
rect 15290 2000 15346 2009
rect 15290 1935 15346 1944
rect 15396 1193 15424 2450
rect 15382 1184 15438 1193
rect 15382 1119 15438 1128
rect 14740 604 14792 610
rect 14740 546 14792 552
rect 14832 604 14884 610
rect 14832 546 14884 552
rect 14752 480 14780 546
rect 15580 480 15608 6695
rect 15672 6322 15700 6734
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15856 5914 15884 6666
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16040 5234 16068 11886
rect 16316 11778 16344 15302
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 16578 13968 16634 13977
rect 16578 13903 16634 13912
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16224 11750 16344 11778
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 11218 16160 11562
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16224 6866 16252 11750
rect 16302 11656 16358 11665
rect 16302 11591 16304 11600
rect 16356 11591 16358 11600
rect 16304 11562 16356 11568
rect 16316 11286 16344 11562
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16408 10266 16436 13126
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16500 10577 16528 10678
rect 16486 10568 16542 10577
rect 16486 10503 16542 10512
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16408 9654 16436 10202
rect 16500 10198 16528 10503
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16316 7954 16344 8366
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16500 7410 16528 9998
rect 16592 9110 16620 13903
rect 16670 13832 16726 13841
rect 16670 13767 16726 13776
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16592 8634 16620 9046
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8022 16712 13767
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 23478 11656 23534 11665
rect 23478 11591 23534 11600
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 16960 10810 16988 11154
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16776 8566 16804 9114
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16868 8022 16896 10542
rect 18524 10538 18552 11154
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17512 9722 17540 10134
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17236 9110 17264 9454
rect 17512 9382 17540 9658
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8498 17264 9046
rect 17406 8936 17462 8945
rect 17406 8871 17462 8880
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17038 8256 17094 8265
rect 17038 8191 17094 8200
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16868 7886 16896 7958
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16868 7546 16896 7822
rect 17052 7818 17080 8191
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16224 6322 16252 6802
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16118 5808 16174 5817
rect 16118 5743 16120 5752
rect 16172 5743 16174 5752
rect 16120 5714 16172 5720
rect 16132 5370 16160 5714
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16408 4826 16436 6734
rect 16500 5846 16528 7142
rect 16854 6896 16910 6905
rect 16854 6831 16856 6840
rect 16908 6831 16910 6840
rect 16856 6802 16908 6808
rect 16578 6216 16634 6225
rect 16578 6151 16580 6160
rect 16632 6151 16634 6160
rect 16580 6122 16632 6128
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16500 5370 16528 5782
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15658 3768 15714 3777
rect 15658 3703 15660 3712
rect 15712 3703 15714 3712
rect 15660 3674 15712 3680
rect 15672 3058 15700 3674
rect 15764 3534 15792 3946
rect 15856 3942 15884 4626
rect 16408 4214 16436 4762
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15856 3641 15884 3878
rect 16500 3670 16528 5306
rect 16592 5098 16620 5850
rect 16868 5710 16896 6802
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16776 4826 16804 5170
rect 17052 5114 17080 7754
rect 17420 7546 17448 8871
rect 17512 7993 17540 9318
rect 17498 7984 17554 7993
rect 17498 7919 17554 7928
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17420 7274 17448 7482
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17420 7002 17448 7210
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17236 6390 17264 6734
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17144 5234 17172 6122
rect 17420 6118 17448 6598
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5846 17448 6054
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17052 5086 17172 5114
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17052 3738 17080 4558
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16488 3664 16540 3670
rect 15842 3632 15898 3641
rect 15842 3567 15898 3576
rect 16302 3632 16358 3641
rect 16488 3606 16540 3612
rect 16302 3567 16358 3576
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15764 3194 15792 3470
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 16316 480 16344 3567
rect 16500 3126 16528 3606
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16500 2922 16528 3062
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16684 2689 16712 3334
rect 16670 2680 16726 2689
rect 16670 2615 16726 2624
rect 16684 2582 16712 2615
rect 16672 2576 16724 2582
rect 17052 2553 17080 3674
rect 16672 2518 16724 2524
rect 17038 2544 17094 2553
rect 17038 2479 17094 2488
rect 17144 480 17172 5086
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17236 2582 17264 4558
rect 17512 3942 17540 4694
rect 17696 4622 17724 10474
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17788 9722 17816 10066
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 6458 17816 9658
rect 17972 9466 18000 9998
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9518 18184 9862
rect 17880 9450 18000 9466
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 17868 9444 18000 9450
rect 17920 9438 18000 9444
rect 17868 9386 17920 9392
rect 18156 9330 18184 9454
rect 18064 9302 18184 9330
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8634 17908 8910
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17972 8129 18000 8842
rect 18064 8514 18092 9302
rect 18064 8486 18184 8514
rect 17958 8120 18014 8129
rect 17958 8055 18014 8064
rect 17972 8022 18000 8055
rect 17960 8016 18012 8022
rect 18156 7970 18184 8486
rect 17960 7958 18012 7964
rect 18064 7942 18184 7970
rect 18064 7018 18092 7942
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18156 7410 18184 7822
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17880 6990 18092 7018
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 5914 17908 6990
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6186 18092 6598
rect 18144 6248 18196 6254
rect 18248 6225 18276 9318
rect 18340 9110 18368 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19076 9722 19104 10066
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18510 9344 18566 9353
rect 18510 9279 18566 9288
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18340 8634 18368 9046
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18420 8560 18472 8566
rect 18418 8528 18420 8537
rect 18472 8528 18474 8537
rect 18418 8463 18474 8472
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18340 7002 18368 7278
rect 18432 7206 18460 7958
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18432 6934 18460 7142
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18524 6780 18552 9279
rect 19076 9194 19104 9658
rect 20180 9654 20208 11018
rect 23492 10130 23520 11591
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 23662 10568 23718 10577
rect 23662 10503 23718 10512
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23492 9722 23520 10066
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 18984 9178 19104 9194
rect 19168 9178 19196 9454
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 18972 9172 19104 9178
rect 19024 9166 19104 9172
rect 19156 9172 19208 9178
rect 18972 9114 19024 9120
rect 19156 9114 19208 9120
rect 19168 8362 19196 9114
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19628 8498 19656 8910
rect 20364 8634 20392 9386
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19168 8090 19196 8298
rect 19352 8090 19380 8434
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19430 8120 19486 8129
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19340 8084 19392 8090
rect 19622 8112 19918 8132
rect 19430 8055 19432 8064
rect 19340 8026 19392 8032
rect 19484 8055 19486 8064
rect 19432 8026 19484 8032
rect 18694 7848 18750 7857
rect 18694 7783 18750 7792
rect 18602 7712 18658 7721
rect 18602 7647 18658 7656
rect 18432 6752 18552 6780
rect 18328 6384 18380 6390
rect 18326 6352 18328 6361
rect 18380 6352 18382 6361
rect 18432 6322 18460 6752
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18326 6287 18382 6296
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18432 6225 18460 6258
rect 18144 6190 18196 6196
rect 18234 6216 18290 6225
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 17960 6112 18012 6118
rect 18064 6089 18092 6122
rect 17960 6054 18012 6060
rect 18050 6080 18106 6089
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17776 5704 17828 5710
rect 17774 5672 17776 5681
rect 17828 5672 17830 5681
rect 17774 5607 17830 5616
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 3097 17356 3334
rect 17314 3088 17370 3097
rect 17314 3023 17316 3032
rect 17368 3023 17370 3032
rect 17316 2994 17368 3000
rect 17328 2963 17356 2994
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17512 2009 17540 3878
rect 17696 3738 17724 3946
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17498 2000 17554 2009
rect 17498 1935 17554 1944
rect 17972 480 18000 6054
rect 18050 6015 18106 6024
rect 18156 5914 18184 6190
rect 18234 6151 18290 6160
rect 18418 6216 18474 6225
rect 18418 6151 18474 6160
rect 18524 5914 18552 6394
rect 18616 6118 18644 7647
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18326 4992 18382 5001
rect 18064 2582 18092 4966
rect 18326 4927 18382 4936
rect 18340 4078 18368 4927
rect 18432 4826 18460 5646
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18156 3777 18184 3878
rect 18142 3768 18198 3777
rect 18142 3703 18198 3712
rect 18340 3670 18368 4014
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18234 3224 18290 3233
rect 18234 3159 18290 3168
rect 18248 2922 18276 3159
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18052 2576 18104 2582
rect 18512 2576 18564 2582
rect 18052 2518 18104 2524
rect 18510 2544 18512 2553
rect 18564 2544 18566 2553
rect 18510 2479 18566 2488
rect 18708 480 18736 7783
rect 19338 7440 19394 7449
rect 19444 7410 19472 8026
rect 19522 7576 19578 7585
rect 19522 7511 19578 7520
rect 19338 7375 19394 7384
rect 19432 7404 19484 7410
rect 19352 7177 19380 7375
rect 19432 7346 19484 7352
rect 19536 7290 19564 7511
rect 19444 7262 19564 7290
rect 19984 7268 20036 7274
rect 19338 7168 19394 7177
rect 19338 7103 19394 7112
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19076 6458 19104 6870
rect 19260 6458 19288 6938
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 18878 6216 18934 6225
rect 18878 6151 18934 6160
rect 18892 5302 18920 6151
rect 19076 5846 19104 6394
rect 19260 6254 19288 6394
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19076 5370 19104 5782
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 19076 4758 19104 5306
rect 19260 5098 19288 5510
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19064 4752 19116 4758
rect 18878 4720 18934 4729
rect 19064 4694 19116 4700
rect 18878 4655 18880 4664
rect 18932 4655 18934 4664
rect 18880 4626 18932 4632
rect 18786 4584 18842 4593
rect 18786 4519 18842 4528
rect 18800 3058 18828 4519
rect 18892 4214 18920 4626
rect 19076 4282 19104 4694
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 19076 3670 19104 4218
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19076 3369 19104 3606
rect 19062 3360 19118 3369
rect 19062 3295 19118 3304
rect 19076 3194 19104 3295
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18800 2446 18828 2994
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19444 626 19472 7262
rect 19984 7210 20036 7216
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19996 7002 20024 7210
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 19996 6905 20024 6938
rect 19982 6896 20038 6905
rect 19982 6831 20038 6840
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19904 6322 19932 6598
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19536 5370 19564 6190
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20088 5914 20116 6190
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19996 5234 20024 5510
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4214 20024 5034
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 20074 4176 20130 4185
rect 20074 4111 20076 4120
rect 20128 4111 20130 4120
rect 20076 4082 20128 4088
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20074 3904 20130 3913
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 3194 19564 3674
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19536 2854 19564 3130
rect 19628 3126 19656 3334
rect 19996 3194 20024 3878
rect 20074 3839 20130 3848
rect 20088 3738 20116 3839
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20350 3360 20406 3369
rect 20350 3295 20406 3304
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19628 2961 19656 3062
rect 19614 2952 19670 2961
rect 19614 2887 19670 2896
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19444 598 19564 626
rect 19536 480 19564 598
rect 20364 480 20392 3295
rect 20456 2650 20484 9590
rect 23676 9518 23704 10503
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20732 8090 20760 8434
rect 20824 8362 20852 8570
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20812 7880 20864 7886
rect 20718 7848 20774 7857
rect 20812 7822 20864 7828
rect 20718 7783 20774 7792
rect 20732 7546 20760 7783
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20732 6730 20760 7278
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20640 5370 20668 5714
rect 20732 5681 20760 6190
rect 20718 5672 20774 5681
rect 20718 5607 20774 5616
rect 20824 5545 20852 7822
rect 20916 6780 20944 8910
rect 21284 8566 21312 9454
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21560 8401 21588 9318
rect 22466 9072 22522 9081
rect 21916 9036 21968 9042
rect 22466 9007 22522 9016
rect 21916 8978 21968 8984
rect 21546 8392 21602 8401
rect 21456 8356 21508 8362
rect 21928 8362 21956 8978
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21546 8327 21602 8336
rect 21916 8356 21968 8362
rect 21456 8298 21508 8304
rect 21916 8298 21968 8304
rect 21086 8256 21142 8265
rect 21086 8191 21142 8200
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 21008 7002 21036 7890
rect 21100 7410 21128 8191
rect 21272 7744 21324 7750
rect 21178 7712 21234 7721
rect 21272 7686 21324 7692
rect 21178 7647 21234 7656
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21192 7274 21220 7647
rect 21284 7449 21312 7686
rect 21270 7440 21326 7449
rect 21270 7375 21326 7384
rect 21284 7342 21312 7375
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 20996 6792 21048 6798
rect 20916 6752 20996 6780
rect 20916 5914 20944 6752
rect 20996 6734 21048 6740
rect 21100 6458 21128 6870
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21086 5672 21142 5681
rect 21086 5607 21142 5616
rect 20810 5536 20866 5545
rect 20810 5471 20866 5480
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 21100 5234 21128 5607
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 4185 20852 4558
rect 20810 4176 20866 4185
rect 20810 4111 20866 4120
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20732 3738 20760 3946
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20916 3670 20944 4966
rect 21100 4842 21128 5170
rect 21008 4826 21128 4842
rect 20996 4820 21128 4826
rect 21048 4814 21128 4820
rect 20996 4762 21048 4768
rect 21192 4321 21220 6938
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21284 6254 21312 6598
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21178 4312 21234 4321
rect 21178 4247 21234 4256
rect 21362 4176 21418 4185
rect 20996 4140 21048 4146
rect 21362 4111 21418 4120
rect 20996 4082 21048 4088
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 21008 3602 21036 4082
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21008 2650 21036 3538
rect 21376 2922 21404 4111
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21468 2854 21496 8298
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21744 7313 21772 7346
rect 21730 7304 21786 7313
rect 21730 7239 21786 7248
rect 21914 7168 21970 7177
rect 21914 7103 21970 7112
rect 21640 6384 21692 6390
rect 21638 6352 21640 6361
rect 21692 6352 21694 6361
rect 21548 6316 21600 6322
rect 21638 6287 21694 6296
rect 21548 6258 21600 6264
rect 21560 6225 21588 6258
rect 21546 6216 21602 6225
rect 21546 6151 21602 6160
rect 21824 6112 21876 6118
rect 21730 6080 21786 6089
rect 21824 6054 21876 6060
rect 21730 6015 21786 6024
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21652 4282 21680 4694
rect 21744 4622 21772 6015
rect 21836 5778 21864 6054
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21928 5234 21956 7103
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21744 4146 21772 4558
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 21928 3738 21956 4966
rect 22020 4162 22048 8774
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22112 6798 22140 8366
rect 22374 7984 22430 7993
rect 22480 7954 22508 9007
rect 23938 8392 23994 8401
rect 23296 8356 23348 8362
rect 23938 8327 23994 8336
rect 23296 8298 23348 8304
rect 22374 7919 22430 7928
rect 22468 7948 22520 7954
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22204 6458 22232 7686
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22204 5914 22232 6394
rect 22388 6361 22416 7919
rect 22468 7890 22520 7896
rect 22480 7546 22508 7890
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22558 6896 22614 6905
rect 22558 6831 22560 6840
rect 22612 6831 22614 6840
rect 22560 6802 22612 6808
rect 22572 6458 22600 6802
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22374 6352 22430 6361
rect 22374 6287 22430 6296
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22388 5778 22416 6287
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22572 5817 22600 5850
rect 22558 5808 22614 5817
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22376 5772 22428 5778
rect 22558 5743 22614 5752
rect 22928 5772 22980 5778
rect 22376 5714 22428 5720
rect 22928 5714 22980 5720
rect 22112 5370 22140 5714
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22388 5302 22416 5714
rect 22940 5370 22968 5714
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22020 4146 22140 4162
rect 22020 4140 22152 4146
rect 22020 4134 22100 4140
rect 22100 4082 22152 4088
rect 22008 4004 22060 4010
rect 22204 3992 22232 4558
rect 22060 3964 22232 3992
rect 22008 3946 22060 3952
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22558 3768 22614 3777
rect 21916 3732 21968 3738
rect 22558 3703 22614 3712
rect 21916 3674 21968 3680
rect 22572 3602 22600 3703
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20548 2310 20576 2450
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 20548 1601 20576 2246
rect 20534 1592 20590 1601
rect 20534 1527 20590 1536
rect 21100 480 21128 2314
rect 21192 1873 21220 2382
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 21178 1864 21234 1873
rect 21178 1799 21234 1808
rect 21928 480 21956 2246
rect 22480 1329 22508 3470
rect 22572 3194 22600 3538
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22664 1986 22692 3878
rect 23308 3641 23336 8298
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23294 3632 23350 3641
rect 23294 3567 23350 3576
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23308 2145 23336 2858
rect 23400 2650 23428 7686
rect 23584 7410 23612 7890
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23492 6390 23520 7142
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23584 4593 23612 7346
rect 23952 6866 23980 8327
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5681 23704 6054
rect 23662 5672 23718 5681
rect 23662 5607 23718 5616
rect 23860 5114 23888 6598
rect 23952 6458 23980 6802
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 24044 5778 24072 9318
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 24044 5370 24072 5714
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24136 5166 24164 9862
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24688 7177 24716 7278
rect 24768 7200 24820 7206
rect 24674 7168 24730 7177
rect 24768 7142 24820 7148
rect 24674 7103 24730 7112
rect 24674 6760 24730 6769
rect 24674 6695 24730 6704
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6254 24716 6695
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24124 5160 24176 5166
rect 24030 5128 24086 5137
rect 23664 5092 23716 5098
rect 23860 5086 23980 5114
rect 23664 5034 23716 5040
rect 23570 4584 23626 4593
rect 23570 4519 23626 4528
rect 23676 4185 23704 5034
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 23662 4176 23718 4185
rect 23662 4111 23718 4120
rect 23570 4040 23626 4049
rect 23570 3975 23626 3984
rect 23664 4004 23716 4010
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23492 3233 23520 3878
rect 23478 3224 23534 3233
rect 23584 3194 23612 3975
rect 23664 3946 23716 3952
rect 23478 3159 23534 3168
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23584 2990 23612 3130
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23676 2802 23704 3946
rect 23860 3913 23888 4966
rect 23952 4078 23980 5086
rect 24124 5102 24176 5108
rect 24030 5063 24086 5072
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23940 3936 23992 3942
rect 23846 3904 23902 3913
rect 23940 3878 23992 3884
rect 23846 3839 23902 3848
rect 23492 2774 23704 2802
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23294 2136 23350 2145
rect 23294 2071 23350 2080
rect 22664 1958 22784 1986
rect 22466 1320 22522 1329
rect 22466 1255 22522 1264
rect 22756 480 22784 1958
rect 23492 480 23520 2774
rect 23952 2553 23980 3878
rect 24044 3738 24072 5063
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 24044 3194 24072 3538
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24044 3097 24072 3130
rect 24030 3088 24086 3097
rect 24030 3023 24086 3032
rect 23938 2544 23994 2553
rect 23848 2508 23900 2514
rect 23938 2479 23994 2488
rect 23848 2450 23900 2456
rect 23860 2417 23888 2450
rect 24032 2440 24084 2446
rect 23846 2408 23902 2417
rect 24032 2382 24084 2388
rect 23846 2343 23902 2352
rect 24044 2009 24072 2382
rect 24030 2000 24086 2009
rect 24030 1935 24086 1944
rect 24136 1737 24164 4422
rect 24228 4049 24256 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24214 4040 24270 4049
rect 24214 3975 24270 3984
rect 24688 3942 24716 4626
rect 24780 4078 24808 7142
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 24860 6384 24912 6390
rect 24858 6352 24860 6361
rect 24912 6352 24914 6361
rect 24858 6287 24914 6296
rect 25148 5778 25176 6598
rect 25516 6118 25544 6802
rect 25504 6112 25556 6118
rect 25502 6080 25504 6089
rect 25556 6080 25558 6089
rect 25502 6015 25558 6024
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 25148 5370 25176 5714
rect 25318 5672 25374 5681
rect 25318 5607 25320 5616
rect 25372 5607 25374 5616
rect 27526 5672 27582 5681
rect 27526 5607 27582 5616
rect 25320 5578 25372 5584
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 26700 5296 26752 5302
rect 26700 5238 26752 5244
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25870 4040 25926 4049
rect 25870 3975 25926 3984
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 24688 3505 24716 3878
rect 24674 3496 24730 3505
rect 24674 3431 24730 3440
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 3120 24268 3126
rect 24216 3062 24268 3068
rect 24122 1728 24178 1737
rect 24122 1663 24178 1672
rect 24228 1442 24256 3062
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24228 1414 24348 1442
rect 24320 480 24348 1414
rect 25148 480 25176 3878
rect 25226 3632 25282 3641
rect 25226 3567 25282 3576
rect 25240 2990 25268 3567
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25596 2440 25648 2446
rect 25594 2408 25596 2417
rect 25648 2408 25650 2417
rect 25594 2343 25650 2352
rect 25884 480 25912 3975
rect 26712 480 26740 5238
rect 27540 480 27568 5607
rect 1398 439 1454 448
rect 1950 0 2006 480
rect 2778 0 2834 480
rect 3514 0 3570 480
rect 4342 0 4398 480
rect 5170 0 5226 480
rect 5906 0 5962 480
rect 6734 0 6790 480
rect 7562 0 7618 480
rect 8298 0 8354 480
rect 9126 0 9182 480
rect 9954 0 10010 480
rect 10690 0 10746 480
rect 11518 0 11574 480
rect 12346 0 12402 480
rect 13082 0 13138 480
rect 13910 0 13966 480
rect 14738 0 14794 480
rect 15566 0 15622 480
rect 16302 0 16358 480
rect 17130 0 17186 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19522 0 19578 480
rect 20350 0 20406 480
rect 21086 0 21142 480
rect 21914 0 21970 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 24306 0 24362 480
rect 25134 0 25190 480
rect 25870 0 25926 480
rect 26698 0 26754 480
rect 27526 0 27582 480
<< via2 >>
rect 1950 27376 2006 27432
rect 1490 26288 1546 26344
rect 1398 25336 1454 25392
rect 1582 24248 1638 24304
rect 1490 23160 1546 23216
rect 1398 21936 1454 21992
rect 1490 21120 1546 21176
rect 1674 20748 1676 20768
rect 1676 20748 1728 20768
rect 1728 20748 1730 20768
rect 1674 20712 1730 20748
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1582 13912 1638 13968
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 1766 14320 1822 14376
rect 1766 13776 1822 13832
rect 1766 12280 1822 12336
rect 1674 11736 1730 11792
rect 1674 11464 1730 11520
rect 2226 15852 2228 15872
rect 2228 15852 2280 15872
rect 2280 15852 2282 15872
rect 2226 15816 2282 15852
rect 2134 15308 2136 15328
rect 2136 15308 2188 15328
rect 2188 15308 2190 15328
rect 2134 15272 2190 15308
rect 2134 13504 2190 13560
rect 2134 12416 2190 12472
rect 2042 11212 2098 11248
rect 2042 11192 2044 11212
rect 2044 11192 2096 11212
rect 2096 11192 2098 11212
rect 1582 9696 1638 9752
rect 1950 9560 2006 9616
rect 1858 8336 1914 8392
rect 1766 6840 1822 6896
rect 1582 6316 1638 6352
rect 1582 6296 1584 6316
rect 1584 6296 1636 6316
rect 1636 6296 1638 6316
rect 1858 5616 1914 5672
rect 1858 5228 1914 5264
rect 1858 5208 1860 5228
rect 1860 5208 1912 5228
rect 1912 5208 1914 5228
rect 2134 9288 2190 9344
rect 2318 9560 2374 9616
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 5538 20032 5594 20088
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 2594 19352 2650 19408
rect 2594 16088 2650 16144
rect 2502 9152 2558 9208
rect 2226 7384 2282 7440
rect 1858 3884 1860 3904
rect 1860 3884 1912 3904
rect 1912 3884 1914 3904
rect 1858 3848 1914 3884
rect 3054 13912 3110 13968
rect 2962 12824 3018 12880
rect 2870 11620 2926 11656
rect 2870 11600 2872 11620
rect 2872 11600 2924 11620
rect 2924 11600 2926 11620
rect 2778 10104 2834 10160
rect 2502 4664 2558 4720
rect 4066 19080 4122 19136
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 4066 17720 4122 17776
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 3698 14864 3754 14920
rect 3514 11872 3570 11928
rect 3514 10004 3516 10024
rect 3516 10004 3568 10024
rect 3568 10004 3570 10024
rect 3514 9968 3570 10004
rect 3790 14068 3846 14104
rect 3790 14048 3792 14068
rect 3792 14048 3844 14068
rect 3844 14048 3846 14068
rect 3698 13368 3754 13424
rect 3790 11056 3846 11112
rect 3698 10920 3754 10976
rect 3606 9560 3662 9616
rect 3054 7656 3110 7712
rect 3330 7248 3386 7304
rect 2686 6332 2688 6352
rect 2688 6332 2740 6352
rect 2740 6332 2742 6352
rect 2686 6296 2742 6332
rect 3054 4140 3110 4176
rect 3054 4120 3056 4140
rect 3056 4120 3108 4140
rect 3108 4120 3110 4140
rect 2502 3712 2558 3768
rect 2410 3576 2466 3632
rect 2042 3304 2098 3360
rect 1122 1128 1178 1184
rect 2134 3032 2190 3088
rect 2318 2624 2374 2680
rect 2686 2372 2742 2408
rect 2686 2352 2688 2372
rect 2688 2352 2740 2372
rect 2740 2352 2742 2372
rect 1950 1944 2006 2000
rect 1398 448 1454 504
rect 3974 13912 4030 13968
rect 3882 10784 3938 10840
rect 4250 13504 4306 13560
rect 3974 9152 4030 9208
rect 3974 8744 4030 8800
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4158 7792 4214 7848
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 3790 6568 3846 6624
rect 3974 6196 3976 6216
rect 3976 6196 4028 6216
rect 4028 6196 4030 6216
rect 3974 6160 4030 6196
rect 3422 992 3478 1048
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4986 10104 5042 10160
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5170 10548 5172 10568
rect 5172 10548 5224 10568
rect 5224 10548 5226 10568
rect 5170 10512 5226 10548
rect 5538 12280 5594 12336
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5722 11636 5724 11656
rect 5724 11636 5776 11656
rect 5776 11636 5778 11656
rect 5722 11600 5778 11636
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6090 9288 6146 9344
rect 5630 9152 5686 9208
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5538 7384 5594 7440
rect 4526 6024 4582 6080
rect 4250 4664 4306 4720
rect 4066 4528 4122 4584
rect 3974 2916 4030 2952
rect 3974 2896 3976 2916
rect 3976 2896 4028 2916
rect 4028 2896 4030 2916
rect 4250 3340 4252 3360
rect 4252 3340 4304 3360
rect 4304 3340 4306 3360
rect 4250 3304 4306 3340
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 10138 18264 10194 18320
rect 9494 16088 9550 16144
rect 6366 13776 6422 13832
rect 6918 11736 6974 11792
rect 7470 13812 7472 13832
rect 7472 13812 7524 13832
rect 7524 13812 7526 13832
rect 7470 13776 7526 13812
rect 7378 12416 7434 12472
rect 6734 11076 6790 11112
rect 6734 11056 6736 11076
rect 6736 11056 6788 11076
rect 6788 11056 6790 11076
rect 6734 10920 6790 10976
rect 5170 6840 5226 6896
rect 6182 6840 6238 6896
rect 4342 2760 4398 2816
rect 3882 2488 3938 2544
rect 4066 2488 4122 2544
rect 3882 1808 3938 1864
rect 4250 1672 4306 1728
rect 4158 1536 4214 1592
rect 3790 1264 3846 1320
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5906 6332 5908 6352
rect 5908 6332 5960 6352
rect 5960 6332 5962 6352
rect 5906 6296 5962 6332
rect 6274 6180 6330 6216
rect 6274 6160 6276 6180
rect 6276 6160 6328 6180
rect 6328 6160 6330 6180
rect 5538 5752 5594 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5262 4684 5318 4720
rect 5262 4664 5264 4684
rect 5264 4664 5316 4684
rect 5316 4664 5318 4684
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6458 8880 6514 8936
rect 6458 8336 6514 8392
rect 6090 3848 6146 3904
rect 5722 3712 5778 3768
rect 5538 3440 5594 3496
rect 5998 3440 6054 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5354 3032 5410 3088
rect 5814 2488 5870 2544
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7194 11464 7250 11520
rect 7378 10512 7434 10568
rect 6182 2896 6238 2952
rect 6274 2372 6330 2408
rect 6274 2352 6276 2372
rect 6276 2352 6328 2372
rect 6328 2352 6330 2372
rect 6182 2080 6238 2136
rect 7654 4256 7710 4312
rect 7930 7948 7986 7984
rect 7930 7928 7932 7948
rect 7932 7928 7984 7948
rect 7984 7928 7986 7948
rect 7838 5480 7894 5536
rect 7838 4392 7894 4448
rect 8666 13096 8722 13152
rect 8390 9560 8446 9616
rect 8206 1400 8262 1456
rect 8758 7284 8760 7304
rect 8760 7284 8812 7304
rect 8812 7284 8814 7304
rect 8758 7248 8814 7284
rect 8758 6060 8760 6080
rect 8760 6060 8812 6080
rect 8812 6060 8814 6080
rect 8758 6024 8814 6060
rect 8758 5108 8760 5128
rect 8760 5108 8812 5128
rect 8812 5108 8814 5128
rect 8758 5072 8814 5108
rect 8666 3712 8722 3768
rect 8574 3304 8630 3360
rect 8758 2080 8814 2136
rect 8666 1808 8722 1864
rect 8482 1536 8538 1592
rect 8758 1536 8814 1592
rect 8482 1264 8538 1320
rect 8482 992 8538 1048
rect 9126 7248 9182 7304
rect 9126 3848 9182 3904
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 11150 17740 11206 17776
rect 11150 17720 11152 17740
rect 11152 17720 11204 17740
rect 11204 17720 11206 17740
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9586 10920 9642 10976
rect 9586 9968 9642 10024
rect 9770 5616 9826 5672
rect 9586 5092 9642 5128
rect 9586 5072 9588 5092
rect 9588 5072 9640 5092
rect 9640 5072 9642 5092
rect 9862 4392 9918 4448
rect 9770 2352 9826 2408
rect 9678 2080 9734 2136
rect 10046 13776 10102 13832
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10690 13948 10692 13968
rect 10692 13948 10744 13968
rect 10744 13948 10746 13968
rect 10690 13912 10746 13948
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10230 12724 10232 12744
rect 10232 12724 10284 12744
rect 10284 12724 10286 12744
rect 10230 12688 10286 12724
rect 10598 12824 10654 12880
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10874 12416 10930 12472
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10414 11228 10416 11248
rect 10416 11228 10468 11248
rect 10468 11228 10470 11248
rect 10414 11192 10470 11228
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10506 10104 10562 10160
rect 10506 9424 10562 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10874 10124 10930 10160
rect 10874 10104 10876 10124
rect 10876 10104 10928 10124
rect 10928 10104 10930 10124
rect 11518 13776 11574 13832
rect 11334 10648 11390 10704
rect 10874 9424 10930 9480
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10782 8372 10784 8392
rect 10784 8372 10836 8392
rect 10836 8372 10838 8392
rect 10782 8336 10838 8372
rect 11058 8880 11114 8936
rect 11058 7812 11114 7848
rect 11058 7792 11060 7812
rect 11060 7792 11112 7812
rect 11112 7792 11114 7812
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10322 6704 10378 6760
rect 10874 6976 10930 7032
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10138 5616 10194 5672
rect 10230 5480 10286 5536
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10782 5752 10838 5808
rect 10782 4800 10838 4856
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10506 1672 10562 1728
rect 11058 7112 11114 7168
rect 10966 4548 11022 4584
rect 10966 4528 10968 4548
rect 10968 4528 11020 4548
rect 11020 4528 11022 4548
rect 10966 3440 11022 3496
rect 10966 3032 11022 3088
rect 11150 2896 11206 2952
rect 11886 10104 11942 10160
rect 12070 12688 12126 12744
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 15474 16632 15530 16688
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 15566 15952 15622 16008
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 12438 13096 12494 13152
rect 11702 4664 11758 4720
rect 11794 4392 11850 4448
rect 11702 3460 11758 3496
rect 11702 3440 11704 3460
rect 11704 3440 11756 3460
rect 11756 3440 11758 3460
rect 12530 9560 12586 9616
rect 12622 9016 12678 9072
rect 12806 9016 12862 9072
rect 12438 8336 12494 8392
rect 12438 7928 12494 7984
rect 12806 6840 12862 6896
rect 12898 6160 12954 6216
rect 13174 10240 13230 10296
rect 13726 9288 13782 9344
rect 12438 5772 12494 5808
rect 12438 5752 12440 5772
rect 12440 5752 12492 5772
rect 12492 5752 12494 5772
rect 12438 4256 12494 4312
rect 12622 4392 12678 4448
rect 12714 3984 12770 4040
rect 11978 2388 11980 2408
rect 11980 2388 12032 2408
rect 12032 2388 12034 2408
rect 11978 2352 12034 2388
rect 12162 2372 12218 2408
rect 12162 2352 12164 2372
rect 12164 2352 12216 2372
rect 12216 2352 12218 2372
rect 13266 5480 13322 5536
rect 13174 4664 13230 4720
rect 13266 3576 13322 3632
rect 13450 7792 13506 7848
rect 13358 3304 13414 3360
rect 13726 7384 13782 7440
rect 13818 6976 13874 7032
rect 13450 2896 13506 2952
rect 13818 1400 13874 1456
rect 15382 13388 15438 13424
rect 15382 13368 15384 13388
rect 15384 13368 15436 13388
rect 15436 13368 15438 13388
rect 14002 13096 14058 13152
rect 14094 9424 14150 9480
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15750 10240 15806 10296
rect 14922 8880 14978 8936
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14738 8472 14794 8528
rect 16026 12724 16028 12744
rect 16028 12724 16080 12744
rect 16080 12724 16082 12744
rect 16026 12688 16082 12724
rect 14278 4936 14334 4992
rect 14554 4800 14610 4856
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14830 6332 14832 6352
rect 14832 6332 14884 6352
rect 14884 6332 14886 6352
rect 14830 6296 14886 6332
rect 14738 5752 14794 5808
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15566 6704 15622 6760
rect 15474 6024 15530 6080
rect 15290 5208 15346 5264
rect 15382 4548 15438 4584
rect 15382 4528 15384 4548
rect 15384 4528 15436 4548
rect 15436 4528 15438 4548
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15382 4256 15438 4312
rect 14094 1944 14150 2000
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15382 3168 15438 3224
rect 15198 2524 15200 2544
rect 15200 2524 15252 2544
rect 15252 2524 15254 2544
rect 15198 2488 15254 2524
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15290 1944 15346 2000
rect 15382 1128 15438 1184
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 16578 13912 16634 13968
rect 16302 11620 16358 11656
rect 16302 11600 16304 11620
rect 16304 11600 16356 11620
rect 16356 11600 16358 11620
rect 16486 10512 16542 10568
rect 16670 13776 16726 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23478 11600 23534 11656
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 17406 8880 17462 8936
rect 17038 8200 17094 8256
rect 16118 5772 16174 5808
rect 16118 5752 16120 5772
rect 16120 5752 16172 5772
rect 16172 5752 16174 5772
rect 16854 6860 16910 6896
rect 16854 6840 16856 6860
rect 16856 6840 16908 6860
rect 16908 6840 16910 6860
rect 16578 6180 16634 6216
rect 16578 6160 16580 6180
rect 16580 6160 16632 6180
rect 16632 6160 16634 6180
rect 15658 3732 15714 3768
rect 15658 3712 15660 3732
rect 15660 3712 15712 3732
rect 15712 3712 15714 3732
rect 17498 7928 17554 7984
rect 15842 3576 15898 3632
rect 16302 3576 16358 3632
rect 16670 2624 16726 2680
rect 17038 2488 17094 2544
rect 17958 8064 18014 8120
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18510 9288 18566 9344
rect 18418 8508 18420 8528
rect 18420 8508 18472 8528
rect 18472 8508 18474 8528
rect 18418 8472 18474 8508
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23662 10512 23718 10568
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19430 8084 19486 8120
rect 19430 8064 19432 8084
rect 19432 8064 19484 8084
rect 19484 8064 19486 8084
rect 18694 7792 18750 7848
rect 18602 7656 18658 7712
rect 18326 6332 18328 6352
rect 18328 6332 18380 6352
rect 18380 6332 18382 6352
rect 18326 6296 18382 6332
rect 17774 5652 17776 5672
rect 17776 5652 17828 5672
rect 17828 5652 17830 5672
rect 17774 5616 17830 5652
rect 17314 3052 17370 3088
rect 17314 3032 17316 3052
rect 17316 3032 17368 3052
rect 17368 3032 17370 3052
rect 17498 1944 17554 2000
rect 18050 6024 18106 6080
rect 18234 6160 18290 6216
rect 18418 6160 18474 6216
rect 18326 4936 18382 4992
rect 18142 3712 18198 3768
rect 18234 3168 18290 3224
rect 18510 2524 18512 2544
rect 18512 2524 18564 2544
rect 18564 2524 18566 2544
rect 18510 2488 18566 2524
rect 19338 7384 19394 7440
rect 19522 7520 19578 7576
rect 19338 7112 19394 7168
rect 18878 6160 18934 6216
rect 18878 4684 18934 4720
rect 18878 4664 18880 4684
rect 18880 4664 18932 4684
rect 18932 4664 18934 4684
rect 18786 4528 18842 4584
rect 19062 3304 19118 3360
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19982 6840 20038 6896
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20074 4140 20130 4176
rect 20074 4120 20076 4140
rect 20076 4120 20128 4140
rect 20128 4120 20130 4140
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20074 3848 20130 3904
rect 20350 3304 20406 3360
rect 19614 2896 19670 2952
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20718 7792 20774 7848
rect 20718 5616 20774 5672
rect 22466 9016 22522 9072
rect 21546 8336 21602 8392
rect 21086 8200 21142 8256
rect 21178 7656 21234 7712
rect 21270 7384 21326 7440
rect 21086 5616 21142 5672
rect 20810 5480 20866 5536
rect 20810 4120 20866 4176
rect 21178 4256 21234 4312
rect 21362 4120 21418 4176
rect 21730 7248 21786 7304
rect 21914 7112 21970 7168
rect 21638 6332 21640 6352
rect 21640 6332 21692 6352
rect 21692 6332 21694 6352
rect 21638 6296 21694 6332
rect 21546 6160 21602 6216
rect 21730 6024 21786 6080
rect 22374 7928 22430 7984
rect 23938 8336 23994 8392
rect 22558 6860 22614 6896
rect 22558 6840 22560 6860
rect 22560 6840 22612 6860
rect 22612 6840 22614 6860
rect 22374 6296 22430 6352
rect 22558 5752 22614 5808
rect 22558 3712 22614 3768
rect 20534 1536 20590 1592
rect 21178 1808 21234 1864
rect 23294 3576 23350 3632
rect 23662 5616 23718 5672
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24674 7112 24730 7168
rect 24674 6704 24730 6760
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23570 4528 23626 4584
rect 23662 4120 23718 4176
rect 23570 3984 23626 4040
rect 23478 3168 23534 3224
rect 24030 5072 24086 5128
rect 23846 3848 23902 3904
rect 23294 2080 23350 2136
rect 22466 1264 22522 1320
rect 24030 3032 24086 3088
rect 23938 2488 23994 2544
rect 23846 2352 23902 2408
rect 24030 1944 24086 2000
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24214 3984 24270 4040
rect 24858 6332 24860 6352
rect 24860 6332 24912 6352
rect 24912 6332 24914 6352
rect 24858 6296 24914 6332
rect 25502 6060 25504 6080
rect 25504 6060 25556 6080
rect 25556 6060 25558 6080
rect 25502 6024 25558 6060
rect 25318 5636 25374 5672
rect 25318 5616 25320 5636
rect 25320 5616 25372 5636
rect 25372 5616 25374 5636
rect 27526 5616 27582 5672
rect 25870 3984 25926 4040
rect 24674 3440 24730 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 1672 24178 1728
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25226 3576 25282 3632
rect 25594 2388 25596 2408
rect 25596 2388 25648 2408
rect 25648 2388 25650 2408
rect 25594 2352 25650 2388
<< metal3 >>
rect 0 27434 480 27464
rect 1945 27434 2011 27437
rect 0 27432 2011 27434
rect 0 27376 1950 27432
rect 2006 27376 2011 27432
rect 0 27374 2011 27376
rect 0 27344 480 27374
rect 1945 27371 2011 27374
rect 0 26346 480 26376
rect 1485 26346 1551 26349
rect 0 26344 1551 26346
rect 0 26288 1490 26344
rect 1546 26288 1551 26344
rect 0 26286 1551 26288
rect 0 26256 480 26286
rect 1485 26283 1551 26286
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 480 25334
rect 1393 25331 1459 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24306 480 24336
rect 1577 24306 1643 24309
rect 0 24304 1643 24306
rect 0 24248 1582 24304
rect 1638 24248 1643 24304
rect 0 24246 1643 24248
rect 0 24216 480 24246
rect 1577 24243 1643 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23218 480 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 480 23158
rect 1485 23155 1551 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 22206 1410 22266
rect 0 22176 480 22206
rect 1350 21997 1410 22206
rect 1350 21992 1459 21997
rect 1350 21936 1398 21992
rect 1454 21936 1459 21992
rect 1350 21934 1459 21936
rect 1393 21931 1459 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10277 21248 10597 21249
rect 0 21178 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1485 21178 1551 21181
rect 0 21176 1551 21178
rect 0 21120 1490 21176
rect 1546 21120 1551 21176
rect 0 21118 1551 21120
rect 0 21088 480 21118
rect 1485 21115 1551 21118
rect 1669 20772 1735 20773
rect 1669 20768 1716 20772
rect 1780 20770 1786 20772
rect 1669 20712 1674 20768
rect 1669 20708 1716 20712
rect 1780 20710 1826 20770
rect 1780 20708 1786 20710
rect 1669 20707 1735 20708
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5533 20090 5599 20093
rect 0 20088 5599 20090
rect 0 20032 5538 20088
rect 5594 20032 5599 20088
rect 0 20030 5599 20032
rect 0 20000 480 20030
rect 5533 20027 5599 20030
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 2589 19412 2655 19413
rect 2589 19408 2636 19412
rect 2700 19410 2706 19412
rect 2589 19352 2594 19408
rect 2589 19348 2636 19352
rect 2700 19350 2746 19410
rect 2700 19348 2706 19350
rect 2589 19347 2655 19348
rect 0 19138 480 19168
rect 4061 19138 4127 19141
rect 0 19136 4127 19138
rect 0 19080 4066 19136
rect 4122 19080 4127 19136
rect 0 19078 4127 19080
rect 0 19048 480 19078
rect 4061 19075 4127 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 10133 18322 10199 18325
rect 1166 18320 10199 18322
rect 1166 18264 10138 18320
rect 10194 18264 10199 18320
rect 1166 18262 10199 18264
rect 0 18050 480 18080
rect 1166 18050 1226 18262
rect 10133 18259 10199 18262
rect 0 17990 1226 18050
rect 1485 18052 1551 18053
rect 1485 18048 1532 18052
rect 1596 18050 1602 18052
rect 1485 17992 1490 18048
rect 0 17960 480 17990
rect 1485 17988 1532 17992
rect 1596 17990 1642 18050
rect 1596 17988 1602 17990
rect 1485 17987 1551 17988
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 4061 17778 4127 17781
rect 11145 17778 11211 17781
rect 4061 17776 11211 17778
rect 4061 17720 4066 17776
rect 4122 17720 11150 17776
rect 11206 17720 11211 17776
rect 4061 17718 11211 17720
rect 4061 17715 4127 17718
rect 11145 17715 11211 17718
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17098 480 17128
rect 0 17038 674 17098
rect 0 17008 480 17038
rect 614 16690 674 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 15469 16690 15535 16693
rect 614 16688 15535 16690
rect 614 16632 15474 16688
rect 15530 16632 15535 16688
rect 614 16630 15535 16632
rect 15469 16627 15535 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2589 16146 2655 16149
rect 9489 16146 9555 16149
rect 2589 16144 9555 16146
rect 2589 16088 2594 16144
rect 2650 16088 9494 16144
rect 9550 16088 9555 16144
rect 2589 16086 9555 16088
rect 2589 16083 2655 16086
rect 9489 16083 9555 16086
rect 0 16010 480 16040
rect 15561 16010 15627 16013
rect 0 16008 15627 16010
rect 0 15952 15566 16008
rect 15622 15952 15627 16008
rect 0 15950 15627 15952
rect 0 15920 480 15950
rect 15561 15947 15627 15950
rect 2221 15876 2287 15877
rect 2221 15874 2268 15876
rect 2176 15872 2268 15874
rect 2176 15816 2226 15872
rect 2176 15814 2268 15816
rect 2221 15812 2268 15814
rect 2332 15812 2338 15876
rect 2221 15811 2287 15812
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 2129 15332 2195 15333
rect 2078 15330 2084 15332
rect 2038 15270 2084 15330
rect 2148 15328 2195 15332
rect 2190 15272 2195 15328
rect 2078 15268 2084 15270
rect 2148 15268 2195 15272
rect 2129 15267 2195 15268
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14922 480 14952
rect 3693 14922 3759 14925
rect 0 14920 3759 14922
rect 0 14864 3698 14920
rect 3754 14864 3759 14920
rect 0 14862 3759 14864
rect 0 14832 480 14862
rect 3693 14859 3759 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1761 14376 1827 14381
rect 1761 14320 1766 14376
rect 1822 14320 1827 14376
rect 1761 14315 1827 14320
rect 1764 14106 1824 14315
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 3785 14106 3851 14109
rect 1764 14104 3851 14106
rect 1764 14048 3790 14104
rect 3846 14048 3851 14104
rect 1764 14046 3851 14048
rect 3785 14043 3851 14046
rect 0 13970 480 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 480 13910
rect 1577 13907 1643 13910
rect 3049 13970 3115 13973
rect 3969 13970 4035 13973
rect 3049 13968 4035 13970
rect 3049 13912 3054 13968
rect 3110 13912 3974 13968
rect 4030 13912 4035 13968
rect 3049 13910 4035 13912
rect 3049 13907 3115 13910
rect 3969 13907 4035 13910
rect 10685 13970 10751 13973
rect 16573 13970 16639 13973
rect 10685 13968 16639 13970
rect 10685 13912 10690 13968
rect 10746 13912 16578 13968
rect 16634 13912 16639 13968
rect 10685 13910 16639 13912
rect 10685 13907 10751 13910
rect 16573 13907 16639 13910
rect 1761 13834 1827 13837
rect 6361 13834 6427 13837
rect 1761 13832 6427 13834
rect 1761 13776 1766 13832
rect 1822 13776 6366 13832
rect 6422 13776 6427 13832
rect 1761 13774 6427 13776
rect 1761 13771 1827 13774
rect 6361 13771 6427 13774
rect 7465 13834 7531 13837
rect 10041 13834 10107 13837
rect 7465 13832 10107 13834
rect 7465 13776 7470 13832
rect 7526 13776 10046 13832
rect 10102 13776 10107 13832
rect 7465 13774 10107 13776
rect 7465 13771 7531 13774
rect 10041 13771 10107 13774
rect 11513 13834 11579 13837
rect 16665 13834 16731 13837
rect 11513 13832 16731 13834
rect 11513 13776 11518 13832
rect 11574 13776 16670 13832
rect 16726 13776 16731 13832
rect 11513 13774 16731 13776
rect 11513 13771 11579 13774
rect 16665 13771 16731 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 2129 13562 2195 13565
rect 4245 13562 4311 13565
rect 2129 13560 4311 13562
rect 2129 13504 2134 13560
rect 2190 13504 4250 13560
rect 4306 13504 4311 13560
rect 2129 13502 4311 13504
rect 2129 13499 2195 13502
rect 4245 13499 4311 13502
rect 3693 13426 3759 13429
rect 15377 13426 15443 13429
rect 3693 13424 15443 13426
rect 3693 13368 3698 13424
rect 3754 13368 15382 13424
rect 15438 13368 15443 13424
rect 3693 13366 15443 13368
rect 3693 13363 3759 13366
rect 15377 13363 15443 13366
rect 8661 13154 8727 13157
rect 12433 13154 12499 13157
rect 13997 13154 14063 13157
rect 8661 13152 14063 13154
rect 8661 13096 8666 13152
rect 8722 13096 12438 13152
rect 12494 13096 14002 13152
rect 14058 13096 14063 13152
rect 8661 13094 14063 13096
rect 8661 13091 8727 13094
rect 12433 13091 12499 13094
rect 13997 13091 14063 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12882 480 12912
rect 2957 12882 3023 12885
rect 0 12880 3023 12882
rect 0 12824 2962 12880
rect 3018 12824 3023 12880
rect 0 12822 3023 12824
rect 0 12792 480 12822
rect 2957 12819 3023 12822
rect 10593 12882 10659 12885
rect 10593 12880 10794 12882
rect 10593 12824 10598 12880
rect 10654 12824 10794 12880
rect 10593 12822 10794 12824
rect 10593 12819 10659 12822
rect 9990 12684 9996 12748
rect 10060 12746 10066 12748
rect 10225 12746 10291 12749
rect 10060 12744 10291 12746
rect 10060 12688 10230 12744
rect 10286 12688 10291 12744
rect 10060 12686 10291 12688
rect 10060 12684 10066 12686
rect 10225 12683 10291 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 2129 12474 2195 12477
rect 7373 12474 7439 12477
rect 2129 12472 7439 12474
rect 2129 12416 2134 12472
rect 2190 12416 7378 12472
rect 7434 12416 7439 12472
rect 2129 12414 7439 12416
rect 10734 12474 10794 12822
rect 12065 12746 12131 12749
rect 16021 12746 16087 12749
rect 12065 12744 16087 12746
rect 12065 12688 12070 12744
rect 12126 12688 16026 12744
rect 16082 12688 16087 12744
rect 12065 12686 16087 12688
rect 12065 12683 12131 12686
rect 16021 12683 16087 12686
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 10869 12474 10935 12477
rect 10734 12472 10935 12474
rect 10734 12416 10874 12472
rect 10930 12416 10935 12472
rect 10734 12414 10935 12416
rect 2129 12411 2195 12414
rect 7373 12411 7439 12414
rect 10869 12411 10935 12414
rect 1761 12338 1827 12341
rect 5533 12338 5599 12341
rect 1761 12336 5599 12338
rect 1761 12280 1766 12336
rect 1822 12280 5538 12336
rect 5594 12280 5599 12336
rect 1761 12278 5599 12280
rect 1761 12275 1827 12278
rect 5533 12275 5599 12278
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 3509 11930 3575 11933
rect 1534 11928 3575 11930
rect 1534 11872 3514 11928
rect 3570 11872 3575 11928
rect 1534 11870 3575 11872
rect 0 11794 480 11824
rect 1534 11794 1594 11870
rect 3509 11867 3575 11870
rect 0 11734 1594 11794
rect 1669 11794 1735 11797
rect 6913 11794 6979 11797
rect 1669 11792 6979 11794
rect 1669 11736 1674 11792
rect 1730 11736 6918 11792
rect 6974 11736 6979 11792
rect 1669 11734 6979 11736
rect 0 11704 480 11734
rect 1669 11731 1735 11734
rect 6913 11731 6979 11734
rect 2865 11658 2931 11661
rect 5717 11658 5783 11661
rect 2865 11656 5783 11658
rect 2865 11600 2870 11656
rect 2926 11600 5722 11656
rect 5778 11600 5783 11656
rect 2865 11598 5783 11600
rect 2865 11595 2931 11598
rect 5717 11595 5783 11598
rect 16297 11658 16363 11661
rect 23473 11658 23539 11661
rect 16297 11656 23539 11658
rect 16297 11600 16302 11656
rect 16358 11600 23478 11656
rect 23534 11600 23539 11656
rect 16297 11598 23539 11600
rect 16297 11595 16363 11598
rect 23473 11595 23539 11598
rect 1669 11522 1735 11525
rect 7189 11522 7255 11525
rect 1669 11520 7255 11522
rect 1669 11464 1674 11520
rect 1730 11464 7194 11520
rect 7250 11464 7255 11520
rect 1669 11462 7255 11464
rect 1669 11459 1735 11462
rect 7189 11459 7255 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2037 11250 2103 11253
rect 10409 11250 10475 11253
rect 2037 11248 10475 11250
rect 2037 11192 2042 11248
rect 2098 11192 10414 11248
rect 10470 11192 10475 11248
rect 2037 11190 10475 11192
rect 2037 11187 2103 11190
rect 10409 11187 10475 11190
rect 3785 11114 3851 11117
rect 6729 11114 6795 11117
rect 3785 11112 6795 11114
rect 3785 11056 3790 11112
rect 3846 11056 6734 11112
rect 6790 11056 6795 11112
rect 3785 11054 6795 11056
rect 3785 11051 3851 11054
rect 6729 11051 6795 11054
rect 3693 10978 3759 10981
rect 6729 10978 6795 10981
rect 9581 10978 9647 10981
rect 3693 10976 4124 10978
rect 3693 10920 3698 10976
rect 3754 10920 4124 10976
rect 3693 10918 4124 10920
rect 3693 10915 3759 10918
rect 0 10842 480 10872
rect 3877 10842 3943 10845
rect 0 10840 3943 10842
rect 0 10784 3882 10840
rect 3938 10784 3943 10840
rect 0 10782 3943 10784
rect 0 10752 480 10782
rect 3877 10779 3943 10782
rect 4064 10706 4124 10918
rect 6729 10976 9647 10978
rect 6729 10920 6734 10976
rect 6790 10920 9586 10976
rect 9642 10920 9647 10976
rect 6729 10918 9647 10920
rect 6729 10915 6795 10918
rect 9581 10915 9647 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 11329 10706 11395 10709
rect 4064 10704 11395 10706
rect 4064 10648 11334 10704
rect 11390 10648 11395 10704
rect 4064 10646 11395 10648
rect 11329 10643 11395 10646
rect 5165 10570 5231 10573
rect 7373 10570 7439 10573
rect 5165 10568 7439 10570
rect 5165 10512 5170 10568
rect 5226 10512 7378 10568
rect 7434 10512 7439 10568
rect 5165 10510 7439 10512
rect 5165 10507 5231 10510
rect 7373 10507 7439 10510
rect 16481 10570 16547 10573
rect 23657 10570 23723 10573
rect 16481 10568 23723 10570
rect 16481 10512 16486 10568
rect 16542 10512 23662 10568
rect 23718 10512 23723 10568
rect 16481 10510 23723 10512
rect 16481 10507 16547 10510
rect 23657 10507 23723 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 13169 10298 13235 10301
rect 15745 10298 15811 10301
rect 13169 10296 15811 10298
rect 13169 10240 13174 10296
rect 13230 10240 15750 10296
rect 15806 10240 15811 10296
rect 13169 10238 15811 10240
rect 13169 10235 13235 10238
rect 15745 10235 15811 10238
rect 2773 10162 2839 10165
rect 4981 10162 5047 10165
rect 2773 10160 5047 10162
rect 2773 10104 2778 10160
rect 2834 10104 4986 10160
rect 5042 10104 5047 10160
rect 2773 10102 5047 10104
rect 2773 10099 2839 10102
rect 4981 10099 5047 10102
rect 9990 10100 9996 10164
rect 10060 10162 10066 10164
rect 10501 10162 10567 10165
rect 10060 10160 10567 10162
rect 10060 10104 10506 10160
rect 10562 10104 10567 10160
rect 10060 10102 10567 10104
rect 10060 10100 10066 10102
rect 10501 10099 10567 10102
rect 10869 10162 10935 10165
rect 11881 10162 11947 10165
rect 10869 10160 11947 10162
rect 10869 10104 10874 10160
rect 10930 10104 11886 10160
rect 11942 10104 11947 10160
rect 10869 10102 11947 10104
rect 10869 10099 10935 10102
rect 11881 10099 11947 10102
rect 3509 10026 3575 10029
rect 9581 10026 9647 10029
rect 3509 10024 9647 10026
rect 3509 9968 3514 10024
rect 3570 9968 9586 10024
rect 9642 9968 9647 10024
rect 3509 9966 9647 9968
rect 3509 9963 3575 9966
rect 9581 9963 9647 9966
rect 5610 9824 5930 9825
rect 0 9754 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 0 9664 480 9694
rect 1577 9691 1643 9694
rect 1945 9618 2011 9621
rect 2078 9618 2084 9620
rect 1945 9616 2084 9618
rect 1945 9560 1950 9616
rect 2006 9560 2084 9616
rect 1945 9558 2084 9560
rect 1945 9555 2011 9558
rect 2078 9556 2084 9558
rect 2148 9556 2154 9620
rect 2313 9618 2379 9621
rect 3601 9618 3667 9621
rect 2313 9616 3667 9618
rect 2313 9560 2318 9616
rect 2374 9560 3606 9616
rect 3662 9560 3667 9616
rect 2313 9558 3667 9560
rect 2313 9555 2379 9558
rect 3601 9555 3667 9558
rect 8385 9618 8451 9621
rect 12525 9618 12591 9621
rect 8385 9616 12591 9618
rect 8385 9560 8390 9616
rect 8446 9560 12530 9616
rect 12586 9560 12591 9616
rect 8385 9558 12591 9560
rect 8385 9555 8451 9558
rect 12525 9555 12591 9558
rect 10501 9482 10567 9485
rect 10726 9482 10732 9484
rect 10501 9480 10732 9482
rect 10501 9424 10506 9480
rect 10562 9424 10732 9480
rect 10501 9422 10732 9424
rect 10501 9419 10567 9422
rect 10726 9420 10732 9422
rect 10796 9420 10802 9484
rect 10869 9482 10935 9485
rect 14089 9482 14155 9485
rect 10869 9480 14155 9482
rect 10869 9424 10874 9480
rect 10930 9424 14094 9480
rect 14150 9424 14155 9480
rect 10869 9422 14155 9424
rect 10869 9419 10935 9422
rect 14089 9419 14155 9422
rect 2129 9346 2195 9349
rect 6085 9346 6151 9349
rect 2129 9344 6151 9346
rect 2129 9288 2134 9344
rect 2190 9288 6090 9344
rect 6146 9288 6151 9344
rect 2129 9286 6151 9288
rect 2129 9283 2195 9286
rect 6085 9283 6151 9286
rect 13721 9346 13787 9349
rect 18505 9346 18571 9349
rect 13721 9344 18571 9346
rect 13721 9288 13726 9344
rect 13782 9288 18510 9344
rect 18566 9288 18571 9344
rect 13721 9286 18571 9288
rect 13721 9283 13787 9286
rect 18505 9283 18571 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2497 9210 2563 9213
rect 3969 9210 4035 9213
rect 5625 9210 5691 9213
rect 2497 9208 5691 9210
rect 2497 9152 2502 9208
rect 2558 9152 3974 9208
rect 4030 9152 5630 9208
rect 5686 9152 5691 9208
rect 2497 9150 5691 9152
rect 2497 9147 2563 9150
rect 3969 9147 4035 9150
rect 5625 9147 5691 9150
rect 12617 9074 12683 9077
rect 12801 9074 12867 9077
rect 22461 9074 22527 9077
rect 12617 9072 22527 9074
rect 12617 9016 12622 9072
rect 12678 9016 12806 9072
rect 12862 9016 22466 9072
rect 22522 9016 22527 9072
rect 12617 9014 22527 9016
rect 12617 9011 12683 9014
rect 12801 9011 12867 9014
rect 22461 9011 22527 9014
rect 6453 8938 6519 8941
rect 11053 8938 11119 8941
rect 6453 8936 11119 8938
rect 6453 8880 6458 8936
rect 6514 8880 11058 8936
rect 11114 8880 11119 8936
rect 6453 8878 11119 8880
rect 6453 8875 6519 8878
rect 11053 8875 11119 8878
rect 14917 8938 14983 8941
rect 17401 8938 17467 8941
rect 14917 8936 17467 8938
rect 14917 8880 14922 8936
rect 14978 8880 17406 8936
rect 17462 8880 17467 8936
rect 14917 8878 17467 8880
rect 14917 8875 14983 8878
rect 17401 8875 17467 8878
rect 0 8802 480 8832
rect 3969 8802 4035 8805
rect 0 8800 4035 8802
rect 0 8744 3974 8800
rect 4030 8744 4035 8800
rect 0 8742 4035 8744
rect 0 8712 480 8742
rect 3969 8739 4035 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 14733 8530 14799 8533
rect 18413 8530 18479 8533
rect 14733 8528 18479 8530
rect 14733 8472 14738 8528
rect 14794 8472 18418 8528
rect 18474 8472 18479 8528
rect 14733 8470 18479 8472
rect 14733 8467 14799 8470
rect 18413 8467 18479 8470
rect 1853 8394 1919 8397
rect 6453 8394 6519 8397
rect 1853 8392 6519 8394
rect 1853 8336 1858 8392
rect 1914 8336 6458 8392
rect 6514 8336 6519 8392
rect 1853 8334 6519 8336
rect 1853 8331 1919 8334
rect 6453 8331 6519 8334
rect 10777 8394 10843 8397
rect 12433 8394 12499 8397
rect 21541 8394 21607 8397
rect 23933 8394 23999 8397
rect 10777 8392 12499 8394
rect 10777 8336 10782 8392
rect 10838 8336 12438 8392
rect 12494 8336 12499 8392
rect 10777 8334 12499 8336
rect 10777 8331 10843 8334
rect 12433 8331 12499 8334
rect 19382 8334 20178 8394
rect 17033 8258 17099 8261
rect 19382 8258 19442 8334
rect 17033 8256 19442 8258
rect 17033 8200 17038 8256
rect 17094 8200 19442 8256
rect 17033 8198 19442 8200
rect 20118 8258 20178 8334
rect 21541 8392 23999 8394
rect 21541 8336 21546 8392
rect 21602 8336 23938 8392
rect 23994 8336 23999 8392
rect 21541 8334 23999 8336
rect 21541 8331 21607 8334
rect 23933 8331 23999 8334
rect 21081 8258 21147 8261
rect 20118 8256 21147 8258
rect 20118 8200 21086 8256
rect 21142 8200 21147 8256
rect 20118 8198 21147 8200
rect 17033 8195 17099 8198
rect 21081 8195 21147 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 17953 8122 18019 8125
rect 19425 8122 19491 8125
rect 17953 8120 19491 8122
rect 17953 8064 17958 8120
rect 18014 8064 19430 8120
rect 19486 8064 19491 8120
rect 17953 8062 19491 8064
rect 17953 8059 18019 8062
rect 19425 8059 19491 8062
rect 7925 7986 7991 7989
rect 12433 7986 12499 7989
rect 7925 7984 12499 7986
rect 7925 7928 7930 7984
rect 7986 7928 12438 7984
rect 12494 7928 12499 7984
rect 7925 7926 12499 7928
rect 7925 7923 7991 7926
rect 12433 7923 12499 7926
rect 17493 7986 17559 7989
rect 22369 7986 22435 7989
rect 17493 7984 22435 7986
rect 17493 7928 17498 7984
rect 17554 7928 22374 7984
rect 22430 7928 22435 7984
rect 17493 7926 22435 7928
rect 17493 7923 17559 7926
rect 22369 7923 22435 7926
rect 4153 7850 4219 7853
rect 11053 7850 11119 7853
rect 4153 7848 11119 7850
rect 4153 7792 4158 7848
rect 4214 7792 11058 7848
rect 11114 7792 11119 7848
rect 4153 7790 11119 7792
rect 4153 7787 4219 7790
rect 11053 7787 11119 7790
rect 13445 7850 13511 7853
rect 18689 7850 18755 7853
rect 20713 7850 20779 7853
rect 13445 7848 20779 7850
rect 13445 7792 13450 7848
rect 13506 7792 18694 7848
rect 18750 7792 20718 7848
rect 20774 7792 20779 7848
rect 13445 7790 20779 7792
rect 13445 7787 13511 7790
rect 18689 7787 18755 7790
rect 20713 7787 20779 7790
rect 0 7714 480 7744
rect 3049 7714 3115 7717
rect 0 7712 3115 7714
rect 0 7656 3054 7712
rect 3110 7656 3115 7712
rect 0 7654 3115 7656
rect 0 7624 480 7654
rect 3049 7651 3115 7654
rect 18597 7714 18663 7717
rect 21173 7714 21239 7717
rect 18597 7712 21239 7714
rect 18597 7656 18602 7712
rect 18658 7656 21178 7712
rect 21234 7656 21239 7712
rect 18597 7654 21239 7656
rect 18597 7651 18663 7654
rect 21173 7651 21239 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 19517 7578 19583 7581
rect 15334 7576 19583 7578
rect 15334 7520 19522 7576
rect 19578 7520 19583 7576
rect 15334 7518 19583 7520
rect 2221 7442 2287 7445
rect 5533 7442 5599 7445
rect 2221 7440 5599 7442
rect 2221 7384 2226 7440
rect 2282 7384 5538 7440
rect 5594 7384 5599 7440
rect 2221 7382 5599 7384
rect 2221 7379 2287 7382
rect 5533 7379 5599 7382
rect 13721 7442 13787 7445
rect 15334 7442 15394 7518
rect 19517 7515 19583 7518
rect 13721 7440 15394 7442
rect 13721 7384 13726 7440
rect 13782 7384 15394 7440
rect 13721 7382 15394 7384
rect 19333 7442 19399 7445
rect 21265 7442 21331 7445
rect 19333 7440 21331 7442
rect 19333 7384 19338 7440
rect 19394 7384 21270 7440
rect 21326 7384 21331 7440
rect 19333 7382 21331 7384
rect 13721 7379 13787 7382
rect 19333 7379 19399 7382
rect 21265 7379 21331 7382
rect 3325 7306 3391 7309
rect 8753 7306 8819 7309
rect 3325 7304 8819 7306
rect 3325 7248 3330 7304
rect 3386 7248 8758 7304
rect 8814 7248 8819 7304
rect 3325 7246 8819 7248
rect 3325 7243 3391 7246
rect 8753 7243 8819 7246
rect 9121 7306 9187 7309
rect 21725 7306 21791 7309
rect 9121 7304 21791 7306
rect 9121 7248 9126 7304
rect 9182 7248 21730 7304
rect 21786 7248 21791 7304
rect 9121 7246 21791 7248
rect 9121 7243 9187 7246
rect 21725 7243 21791 7246
rect 11053 7170 11119 7173
rect 19333 7170 19399 7173
rect 11053 7168 19399 7170
rect 11053 7112 11058 7168
rect 11114 7112 19338 7168
rect 19394 7112 19399 7168
rect 11053 7110 19399 7112
rect 11053 7107 11119 7110
rect 19333 7107 19399 7110
rect 21909 7170 21975 7173
rect 24669 7170 24735 7173
rect 21909 7168 24735 7170
rect 21909 7112 21914 7168
rect 21970 7112 24674 7168
rect 24730 7112 24735 7168
rect 21909 7110 24735 7112
rect 21909 7107 21975 7110
rect 24669 7107 24735 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 10869 7034 10935 7037
rect 13813 7034 13879 7037
rect 10869 7032 13879 7034
rect 10869 6976 10874 7032
rect 10930 6976 13818 7032
rect 13874 6976 13879 7032
rect 10869 6974 13879 6976
rect 10869 6971 10935 6974
rect 13813 6971 13879 6974
rect 1761 6898 1827 6901
rect 4061 6898 4127 6901
rect 1761 6896 4127 6898
rect 1761 6840 1766 6896
rect 1822 6840 4066 6896
rect 4122 6840 4127 6896
rect 1761 6838 4127 6840
rect 1761 6835 1827 6838
rect 4061 6835 4127 6838
rect 5165 6898 5231 6901
rect 6177 6898 6243 6901
rect 5165 6896 6243 6898
rect 5165 6840 5170 6896
rect 5226 6840 6182 6896
rect 6238 6840 6243 6896
rect 5165 6838 6243 6840
rect 5165 6835 5231 6838
rect 6177 6835 6243 6838
rect 12801 6898 12867 6901
rect 16849 6898 16915 6901
rect 12801 6896 16915 6898
rect 12801 6840 12806 6896
rect 12862 6840 16854 6896
rect 16910 6840 16915 6896
rect 12801 6838 16915 6840
rect 12801 6835 12867 6838
rect 16849 6835 16915 6838
rect 19977 6898 20043 6901
rect 22553 6898 22619 6901
rect 19977 6896 22619 6898
rect 19977 6840 19982 6896
rect 20038 6840 22558 6896
rect 22614 6840 22619 6896
rect 19977 6838 22619 6840
rect 19977 6835 20043 6838
rect 22553 6835 22619 6838
rect 10317 6762 10383 6765
rect 10726 6762 10732 6764
rect 10317 6760 10732 6762
rect 10317 6704 10322 6760
rect 10378 6704 10732 6760
rect 10317 6702 10732 6704
rect 10317 6699 10383 6702
rect 10726 6700 10732 6702
rect 10796 6762 10802 6764
rect 15561 6762 15627 6765
rect 24669 6762 24735 6765
rect 10796 6760 24735 6762
rect 10796 6704 15566 6760
rect 15622 6704 24674 6760
rect 24730 6704 24735 6760
rect 10796 6702 24735 6704
rect 10796 6700 10802 6702
rect 15561 6699 15627 6702
rect 24669 6699 24735 6702
rect 0 6626 480 6656
rect 3785 6626 3851 6629
rect 0 6624 3851 6626
rect 0 6568 3790 6624
rect 3846 6568 3851 6624
rect 0 6566 3851 6568
rect 0 6536 480 6566
rect 3785 6563 3851 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 1577 6354 1643 6357
rect 1710 6354 1716 6356
rect 1577 6352 1716 6354
rect 1577 6296 1582 6352
rect 1638 6296 1716 6352
rect 1577 6294 1716 6296
rect 1577 6291 1643 6294
rect 1710 6292 1716 6294
rect 1780 6292 1786 6356
rect 2681 6354 2747 6357
rect 5901 6354 5967 6357
rect 2681 6352 5967 6354
rect 2681 6296 2686 6352
rect 2742 6296 5906 6352
rect 5962 6296 5967 6352
rect 2681 6294 5967 6296
rect 2681 6291 2747 6294
rect 5901 6291 5967 6294
rect 14825 6354 14891 6357
rect 18321 6354 18387 6357
rect 21633 6354 21699 6357
rect 14825 6352 21699 6354
rect 14825 6296 14830 6352
rect 14886 6296 18326 6352
rect 18382 6296 21638 6352
rect 21694 6296 21699 6352
rect 14825 6294 21699 6296
rect 14825 6291 14891 6294
rect 18321 6291 18387 6294
rect 21633 6291 21699 6294
rect 22369 6354 22435 6357
rect 24853 6354 24919 6357
rect 22369 6352 24919 6354
rect 22369 6296 22374 6352
rect 22430 6296 24858 6352
rect 24914 6296 24919 6352
rect 22369 6294 24919 6296
rect 22369 6291 22435 6294
rect 24853 6291 24919 6294
rect 3969 6218 4035 6221
rect 6269 6218 6335 6221
rect 12893 6218 12959 6221
rect 3969 6216 12959 6218
rect 3969 6160 3974 6216
rect 4030 6160 6274 6216
rect 6330 6160 12898 6216
rect 12954 6160 12959 6216
rect 3969 6158 12959 6160
rect 3969 6155 4035 6158
rect 6269 6155 6335 6158
rect 12893 6155 12959 6158
rect 16573 6218 16639 6221
rect 18229 6218 18295 6221
rect 16573 6216 18295 6218
rect 16573 6160 16578 6216
rect 16634 6160 18234 6216
rect 18290 6160 18295 6216
rect 16573 6158 18295 6160
rect 16573 6155 16639 6158
rect 18229 6155 18295 6158
rect 18413 6218 18479 6221
rect 18873 6218 18939 6221
rect 21541 6218 21607 6221
rect 18413 6216 21607 6218
rect 18413 6160 18418 6216
rect 18474 6160 18878 6216
rect 18934 6160 21546 6216
rect 21602 6160 21607 6216
rect 18413 6158 21607 6160
rect 18413 6155 18479 6158
rect 18873 6155 18939 6158
rect 21541 6155 21607 6158
rect 4521 6082 4587 6085
rect 8753 6082 8819 6085
rect 4521 6080 8819 6082
rect 4521 6024 4526 6080
rect 4582 6024 8758 6080
rect 8814 6024 8819 6080
rect 4521 6022 8819 6024
rect 4521 6019 4587 6022
rect 8753 6019 8819 6022
rect 15469 6082 15535 6085
rect 18045 6082 18111 6085
rect 15469 6080 18111 6082
rect 15469 6024 15474 6080
rect 15530 6024 18050 6080
rect 18106 6024 18111 6080
rect 15469 6022 18111 6024
rect 15469 6019 15535 6022
rect 18045 6019 18111 6022
rect 21725 6082 21791 6085
rect 25497 6082 25563 6085
rect 21725 6080 25563 6082
rect 21725 6024 21730 6080
rect 21786 6024 25502 6080
rect 25558 6024 25563 6080
rect 21725 6022 25563 6024
rect 21725 6019 21791 6022
rect 25497 6019 25563 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 5533 5810 5599 5813
rect 10777 5810 10843 5813
rect 5533 5808 10843 5810
rect 5533 5752 5538 5808
rect 5594 5752 10782 5808
rect 10838 5752 10843 5808
rect 5533 5750 10843 5752
rect 5533 5747 5599 5750
rect 10777 5747 10843 5750
rect 12433 5810 12499 5813
rect 14733 5810 14799 5813
rect 12433 5808 14799 5810
rect 12433 5752 12438 5808
rect 12494 5752 14738 5808
rect 14794 5752 14799 5808
rect 12433 5750 14799 5752
rect 12433 5747 12499 5750
rect 14733 5747 14799 5750
rect 16113 5810 16179 5813
rect 22553 5810 22619 5813
rect 16113 5808 22619 5810
rect 16113 5752 16118 5808
rect 16174 5752 22558 5808
rect 22614 5752 22619 5808
rect 16113 5750 22619 5752
rect 16113 5747 16179 5750
rect 22553 5747 22619 5750
rect 0 5674 480 5704
rect 1853 5674 1919 5677
rect 0 5672 1919 5674
rect 0 5616 1858 5672
rect 1914 5616 1919 5672
rect 0 5614 1919 5616
rect 0 5584 480 5614
rect 1853 5611 1919 5614
rect 9765 5674 9831 5677
rect 10133 5674 10199 5677
rect 17769 5674 17835 5677
rect 20713 5674 20779 5677
rect 9765 5672 10199 5674
rect 9765 5616 9770 5672
rect 9826 5616 10138 5672
rect 10194 5616 10199 5672
rect 9765 5614 10199 5616
rect 9765 5611 9831 5614
rect 10133 5611 10199 5614
rect 14782 5614 15394 5674
rect 7833 5538 7899 5541
rect 10225 5538 10291 5541
rect 7833 5536 10291 5538
rect 7833 5480 7838 5536
rect 7894 5480 10230 5536
rect 10286 5480 10291 5536
rect 7833 5478 10291 5480
rect 7833 5475 7899 5478
rect 10225 5475 10291 5478
rect 13261 5538 13327 5541
rect 14782 5538 14842 5614
rect 13261 5536 14842 5538
rect 13261 5480 13266 5536
rect 13322 5480 14842 5536
rect 13261 5478 14842 5480
rect 15334 5538 15394 5614
rect 17769 5672 20779 5674
rect 17769 5616 17774 5672
rect 17830 5616 20718 5672
rect 20774 5616 20779 5672
rect 17769 5614 20779 5616
rect 17769 5611 17835 5614
rect 20713 5611 20779 5614
rect 21081 5674 21147 5677
rect 23657 5674 23723 5677
rect 21081 5672 23723 5674
rect 21081 5616 21086 5672
rect 21142 5616 23662 5672
rect 23718 5616 23723 5672
rect 21081 5614 23723 5616
rect 21081 5611 21147 5614
rect 23657 5611 23723 5614
rect 25313 5674 25379 5677
rect 27521 5674 27587 5677
rect 25313 5672 27587 5674
rect 25313 5616 25318 5672
rect 25374 5616 27526 5672
rect 27582 5616 27587 5672
rect 25313 5614 27587 5616
rect 25313 5611 25379 5614
rect 27521 5611 27587 5614
rect 20805 5538 20871 5541
rect 15334 5536 20871 5538
rect 15334 5480 20810 5536
rect 20866 5480 20871 5536
rect 15334 5478 20871 5480
rect 13261 5475 13327 5478
rect 20805 5475 20871 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 1853 5266 1919 5269
rect 15285 5266 15351 5269
rect 1853 5264 15351 5266
rect 1853 5208 1858 5264
rect 1914 5208 15290 5264
rect 15346 5208 15351 5264
rect 1853 5206 15351 5208
rect 1853 5203 1919 5206
rect 15285 5203 15351 5206
rect 8753 5130 8819 5133
rect 9581 5130 9647 5133
rect 24025 5130 24091 5133
rect 8753 5128 24091 5130
rect 8753 5072 8758 5128
rect 8814 5072 9586 5128
rect 9642 5072 24030 5128
rect 24086 5072 24091 5128
rect 8753 5070 24091 5072
rect 8753 5067 8819 5070
rect 9581 5067 9647 5070
rect 24025 5067 24091 5070
rect 14273 4994 14339 4997
rect 18321 4994 18387 4997
rect 14273 4992 18387 4994
rect 14273 4936 14278 4992
rect 14334 4936 18326 4992
rect 18382 4936 18387 4992
rect 14273 4934 18387 4936
rect 14273 4931 14339 4934
rect 18321 4931 18387 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 10777 4858 10843 4861
rect 14549 4858 14615 4861
rect 10777 4856 14615 4858
rect 10777 4800 10782 4856
rect 10838 4800 14554 4856
rect 14610 4800 14615 4856
rect 10777 4798 14615 4800
rect 10777 4795 10843 4798
rect 14549 4795 14615 4798
rect 2497 4722 2563 4725
rect 4245 4722 4311 4725
rect 2497 4720 4311 4722
rect 2497 4664 2502 4720
rect 2558 4664 4250 4720
rect 4306 4664 4311 4720
rect 2497 4662 4311 4664
rect 2497 4659 2563 4662
rect 4245 4659 4311 4662
rect 5257 4722 5323 4725
rect 11697 4722 11763 4725
rect 5257 4720 11763 4722
rect 5257 4664 5262 4720
rect 5318 4664 11702 4720
rect 11758 4664 11763 4720
rect 5257 4662 11763 4664
rect 5257 4659 5323 4662
rect 11697 4659 11763 4662
rect 13169 4722 13235 4725
rect 18873 4722 18939 4725
rect 13169 4720 18939 4722
rect 13169 4664 13174 4720
rect 13230 4664 18878 4720
rect 18934 4664 18939 4720
rect 13169 4662 18939 4664
rect 13169 4659 13235 4662
rect 18873 4659 18939 4662
rect 0 4586 480 4616
rect 4061 4586 4127 4589
rect 10961 4586 11027 4589
rect 15377 4586 15443 4589
rect 0 4584 4127 4586
rect 0 4528 4066 4584
rect 4122 4528 4127 4584
rect 0 4526 4127 4528
rect 0 4496 480 4526
rect 4061 4523 4127 4526
rect 5398 4584 11027 4586
rect 5398 4528 10966 4584
rect 11022 4528 11027 4584
rect 5398 4526 11027 4528
rect 2262 4388 2268 4452
rect 2332 4450 2338 4452
rect 5398 4450 5458 4526
rect 10961 4523 11027 4526
rect 12942 4584 15443 4586
rect 12942 4528 15382 4584
rect 15438 4528 15443 4584
rect 12942 4526 15443 4528
rect 2332 4390 5458 4450
rect 7833 4450 7899 4453
rect 9857 4450 9923 4453
rect 7833 4448 9923 4450
rect 7833 4392 7838 4448
rect 7894 4392 9862 4448
rect 9918 4392 9923 4448
rect 7833 4390 9923 4392
rect 2332 4388 2338 4390
rect 7833 4387 7899 4390
rect 9857 4387 9923 4390
rect 11789 4450 11855 4453
rect 12617 4450 12683 4453
rect 12942 4450 13002 4526
rect 15377 4523 15443 4526
rect 18781 4586 18847 4589
rect 23565 4586 23631 4589
rect 18781 4584 23631 4586
rect 18781 4528 18786 4584
rect 18842 4528 23570 4584
rect 23626 4528 23631 4584
rect 18781 4526 23631 4528
rect 18781 4523 18847 4526
rect 23565 4523 23631 4526
rect 11789 4448 13002 4450
rect 11789 4392 11794 4448
rect 11850 4392 12622 4448
rect 12678 4392 13002 4448
rect 11789 4390 13002 4392
rect 11789 4387 11855 4390
rect 12617 4387 12683 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7649 4314 7715 4317
rect 12433 4314 12499 4317
rect 7649 4312 12499 4314
rect 7649 4256 7654 4312
rect 7710 4256 12438 4312
rect 12494 4256 12499 4312
rect 7649 4254 12499 4256
rect 7649 4251 7715 4254
rect 12433 4251 12499 4254
rect 15377 4314 15443 4317
rect 21173 4314 21239 4317
rect 15377 4312 21239 4314
rect 15377 4256 15382 4312
rect 15438 4256 21178 4312
rect 21234 4256 21239 4312
rect 15377 4254 21239 4256
rect 15377 4251 15443 4254
rect 21173 4251 21239 4254
rect 3049 4178 3115 4181
rect 20069 4178 20135 4181
rect 20805 4178 20871 4181
rect 3049 4176 20871 4178
rect 3049 4120 3054 4176
rect 3110 4120 20074 4176
rect 20130 4120 20810 4176
rect 20866 4120 20871 4176
rect 3049 4118 20871 4120
rect 3049 4115 3115 4118
rect 20069 4115 20135 4118
rect 20805 4115 20871 4118
rect 21357 4178 21423 4181
rect 23657 4178 23723 4181
rect 21357 4176 23723 4178
rect 21357 4120 21362 4176
rect 21418 4120 23662 4176
rect 23718 4120 23723 4176
rect 21357 4118 23723 4120
rect 21357 4115 21423 4118
rect 23657 4115 23723 4118
rect 1526 3980 1532 4044
rect 1596 4042 1602 4044
rect 12709 4042 12775 4045
rect 23565 4042 23631 4045
rect 1596 4040 12775 4042
rect 1596 3984 12714 4040
rect 12770 3984 12775 4040
rect 1596 3982 12775 3984
rect 1596 3980 1602 3982
rect 12709 3979 12775 3982
rect 14414 4040 23631 4042
rect 14414 3984 23570 4040
rect 23626 3984 23631 4040
rect 14414 3982 23631 3984
rect 1853 3906 1919 3909
rect 2262 3906 2268 3908
rect 1853 3904 2268 3906
rect 1853 3848 1858 3904
rect 1914 3848 2268 3904
rect 1853 3846 2268 3848
rect 1853 3843 1919 3846
rect 2262 3844 2268 3846
rect 2332 3844 2338 3908
rect 6085 3906 6151 3909
rect 9121 3906 9187 3909
rect 6085 3904 9187 3906
rect 6085 3848 6090 3904
rect 6146 3848 9126 3904
rect 9182 3848 9187 3904
rect 6085 3846 9187 3848
rect 6085 3843 6151 3846
rect 9121 3843 9187 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 2497 3770 2563 3773
rect 2630 3770 2636 3772
rect 2497 3768 2636 3770
rect 2497 3712 2502 3768
rect 2558 3712 2636 3768
rect 2497 3710 2636 3712
rect 2497 3707 2563 3710
rect 2630 3708 2636 3710
rect 2700 3708 2706 3772
rect 5717 3770 5783 3773
rect 6126 3770 6132 3772
rect 5582 3768 6132 3770
rect 5582 3712 5722 3768
rect 5778 3712 6132 3768
rect 5582 3710 6132 3712
rect 2405 3634 2471 3637
rect 5582 3634 5642 3710
rect 5717 3707 5783 3710
rect 6126 3708 6132 3710
rect 6196 3708 6202 3772
rect 8661 3770 8727 3773
rect 14414 3770 14474 3982
rect 23565 3979 23631 3982
rect 24209 4042 24275 4045
rect 25865 4042 25931 4045
rect 24209 4040 25931 4042
rect 24209 3984 24214 4040
rect 24270 3984 25870 4040
rect 25926 3984 25931 4040
rect 24209 3982 25931 3984
rect 24209 3979 24275 3982
rect 25865 3979 25931 3982
rect 20069 3906 20135 3909
rect 23841 3906 23907 3909
rect 20069 3904 23907 3906
rect 20069 3848 20074 3904
rect 20130 3848 23846 3904
rect 23902 3848 23907 3904
rect 20069 3846 23907 3848
rect 20069 3843 20135 3846
rect 23841 3843 23907 3846
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 8661 3768 10196 3770
rect 8661 3712 8666 3768
rect 8722 3712 10196 3768
rect 8661 3710 10196 3712
rect 8661 3707 8727 3710
rect 2405 3632 5642 3634
rect 2405 3576 2410 3632
rect 2466 3576 5642 3632
rect 2405 3574 5642 3576
rect 10136 3634 10196 3710
rect 10688 3710 14474 3770
rect 15653 3770 15719 3773
rect 18137 3770 18203 3773
rect 22553 3772 22619 3773
rect 15653 3768 18203 3770
rect 15653 3712 15658 3768
rect 15714 3712 18142 3768
rect 18198 3712 18203 3768
rect 15653 3710 18203 3712
rect 10688 3668 10748 3710
rect 15653 3707 15719 3710
rect 18137 3707 18203 3710
rect 22502 3708 22508 3772
rect 22572 3770 22619 3772
rect 22572 3768 22664 3770
rect 22614 3712 22664 3768
rect 22572 3710 22664 3712
rect 22572 3708 22619 3710
rect 22553 3707 22619 3708
rect 10550 3634 10748 3668
rect 10136 3608 10748 3634
rect 13261 3634 13327 3637
rect 15837 3634 15903 3637
rect 16297 3634 16363 3637
rect 13261 3632 16363 3634
rect 10136 3574 10610 3608
rect 13261 3576 13266 3632
rect 13322 3576 15842 3632
rect 15898 3576 16302 3632
rect 16358 3576 16363 3632
rect 13261 3574 16363 3576
rect 2405 3571 2471 3574
rect 13261 3571 13327 3574
rect 15837 3571 15903 3574
rect 16297 3571 16363 3574
rect 23289 3634 23355 3637
rect 25221 3634 25287 3637
rect 23289 3632 25287 3634
rect 23289 3576 23294 3632
rect 23350 3576 25226 3632
rect 25282 3576 25287 3632
rect 23289 3574 25287 3576
rect 23289 3571 23355 3574
rect 25221 3571 25287 3574
rect 0 3498 480 3528
rect 5533 3498 5599 3501
rect 0 3496 5599 3498
rect 0 3440 5538 3496
rect 5594 3440 5599 3496
rect 0 3438 5599 3440
rect 0 3408 480 3438
rect 5533 3435 5599 3438
rect 5993 3498 6059 3501
rect 10961 3498 11027 3501
rect 5993 3496 11027 3498
rect 5993 3440 5998 3496
rect 6054 3440 10966 3496
rect 11022 3440 11027 3496
rect 5993 3438 11027 3440
rect 5993 3435 6059 3438
rect 10961 3435 11027 3438
rect 11697 3498 11763 3501
rect 24669 3498 24735 3501
rect 11697 3496 24735 3498
rect 11697 3440 11702 3496
rect 11758 3440 24674 3496
rect 24730 3440 24735 3496
rect 11697 3438 24735 3440
rect 11697 3435 11763 3438
rect 24669 3435 24735 3438
rect 2037 3362 2103 3365
rect 4245 3362 4311 3365
rect 2037 3360 4311 3362
rect 2037 3304 2042 3360
rect 2098 3304 4250 3360
rect 4306 3304 4311 3360
rect 2037 3302 4311 3304
rect 2037 3299 2103 3302
rect 4245 3299 4311 3302
rect 8569 3362 8635 3365
rect 13353 3362 13419 3365
rect 8569 3360 13419 3362
rect 8569 3304 8574 3360
rect 8630 3304 13358 3360
rect 13414 3304 13419 3360
rect 8569 3302 13419 3304
rect 8569 3299 8635 3302
rect 13353 3299 13419 3302
rect 19057 3362 19123 3365
rect 20345 3362 20411 3365
rect 19057 3360 20411 3362
rect 19057 3304 19062 3360
rect 19118 3304 20350 3360
rect 20406 3304 20411 3360
rect 19057 3302 20411 3304
rect 19057 3299 19123 3302
rect 20345 3299 20411 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 15377 3226 15443 3229
rect 18229 3226 18295 3229
rect 23473 3226 23539 3229
rect 15377 3224 17602 3226
rect 15377 3168 15382 3224
rect 15438 3168 17602 3224
rect 15377 3166 17602 3168
rect 15377 3163 15443 3166
rect 2129 3090 2195 3093
rect 5349 3090 5415 3093
rect 2129 3088 5415 3090
rect 2129 3032 2134 3088
rect 2190 3032 5354 3088
rect 5410 3032 5415 3088
rect 2129 3030 5415 3032
rect 2129 3027 2195 3030
rect 5349 3027 5415 3030
rect 10961 3090 11027 3093
rect 17309 3090 17375 3093
rect 10961 3088 17375 3090
rect 10961 3032 10966 3088
rect 11022 3032 17314 3088
rect 17370 3032 17375 3088
rect 10961 3030 17375 3032
rect 17542 3090 17602 3166
rect 18229 3224 23539 3226
rect 18229 3168 18234 3224
rect 18290 3168 23478 3224
rect 23534 3168 23539 3224
rect 18229 3166 23539 3168
rect 18229 3163 18295 3166
rect 23473 3163 23539 3166
rect 24025 3090 24091 3093
rect 17542 3088 24091 3090
rect 17542 3032 24030 3088
rect 24086 3032 24091 3088
rect 17542 3030 24091 3032
rect 10961 3027 11027 3030
rect 17309 3027 17375 3030
rect 24025 3027 24091 3030
rect 3969 2954 4035 2957
rect 6177 2954 6243 2957
rect 11145 2954 11211 2957
rect 3969 2952 6243 2954
rect 3969 2896 3974 2952
rect 4030 2896 6182 2952
rect 6238 2896 6243 2952
rect 3969 2894 6243 2896
rect 3969 2891 4035 2894
rect 6177 2891 6243 2894
rect 9998 2952 11211 2954
rect 9998 2896 11150 2952
rect 11206 2896 11211 2952
rect 9998 2894 11211 2896
rect 4337 2818 4403 2821
rect 9998 2818 10058 2894
rect 11145 2891 11211 2894
rect 13445 2954 13511 2957
rect 19609 2954 19675 2957
rect 13445 2952 19675 2954
rect 13445 2896 13450 2952
rect 13506 2896 19614 2952
rect 19670 2896 19675 2952
rect 13445 2894 19675 2896
rect 13445 2891 13511 2894
rect 19609 2891 19675 2894
rect 4337 2816 10058 2818
rect 4337 2760 4342 2816
rect 4398 2760 10058 2816
rect 4337 2758 10058 2760
rect 4337 2755 4403 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2313 2682 2379 2685
rect 16665 2682 16731 2685
rect 2313 2680 7666 2682
rect 2313 2624 2318 2680
rect 2374 2624 7666 2680
rect 2313 2622 7666 2624
rect 2313 2619 2379 2622
rect 0 2546 480 2576
rect 3877 2546 3943 2549
rect 0 2544 3943 2546
rect 0 2488 3882 2544
rect 3938 2488 3943 2544
rect 0 2486 3943 2488
rect 0 2456 480 2486
rect 3877 2483 3943 2486
rect 4061 2546 4127 2549
rect 5809 2546 5875 2549
rect 4061 2544 5875 2546
rect 4061 2488 4066 2544
rect 4122 2488 5814 2544
rect 5870 2488 5875 2544
rect 4061 2486 5875 2488
rect 7606 2546 7666 2622
rect 16665 2680 17602 2682
rect 16665 2624 16670 2680
rect 16726 2624 17602 2680
rect 16665 2622 17602 2624
rect 16665 2619 16731 2622
rect 15193 2546 15259 2549
rect 7606 2544 15259 2546
rect 7606 2488 15198 2544
rect 15254 2488 15259 2544
rect 7606 2486 15259 2488
rect 4061 2483 4127 2486
rect 5809 2483 5875 2486
rect 15193 2483 15259 2486
rect 17033 2546 17099 2549
rect 17033 2544 17372 2546
rect 17033 2488 17038 2544
rect 17094 2488 17372 2544
rect 17033 2486 17372 2488
rect 17033 2483 17099 2486
rect 2681 2410 2747 2413
rect 6269 2410 6335 2413
rect 2681 2408 6335 2410
rect 2681 2352 2686 2408
rect 2742 2352 6274 2408
rect 6330 2352 6335 2408
rect 2681 2350 6335 2352
rect 2681 2347 2747 2350
rect 6269 2347 6335 2350
rect 9765 2410 9831 2413
rect 11973 2410 12039 2413
rect 9765 2408 12039 2410
rect 9765 2352 9770 2408
rect 9826 2352 11978 2408
rect 12034 2352 12039 2408
rect 9765 2350 12039 2352
rect 9765 2347 9831 2350
rect 11973 2347 12039 2350
rect 12157 2410 12223 2413
rect 12157 2408 17234 2410
rect 12157 2352 12162 2408
rect 12218 2352 17234 2408
rect 12157 2350 17234 2352
rect 12157 2347 12223 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 6177 2138 6243 2141
rect 8753 2138 8819 2141
rect 6177 2136 8819 2138
rect 6177 2080 6182 2136
rect 6238 2080 8758 2136
rect 8814 2080 8819 2136
rect 6177 2078 8819 2080
rect 6177 2075 6243 2078
rect 8753 2075 8819 2078
rect 9673 2138 9739 2141
rect 17174 2138 17234 2350
rect 17312 2274 17372 2486
rect 17542 2410 17602 2622
rect 18505 2546 18571 2549
rect 23933 2546 23999 2549
rect 18505 2544 23999 2546
rect 18505 2488 18510 2544
rect 18566 2488 23938 2544
rect 23994 2488 23999 2544
rect 18505 2486 23999 2488
rect 18505 2483 18571 2486
rect 23933 2483 23999 2486
rect 23841 2410 23907 2413
rect 25589 2410 25655 2413
rect 17542 2408 23907 2410
rect 17542 2352 23846 2408
rect 23902 2352 23907 2408
rect 17542 2350 23907 2352
rect 23841 2347 23907 2350
rect 23982 2408 25655 2410
rect 23982 2352 25594 2408
rect 25650 2352 25655 2408
rect 23982 2350 25655 2352
rect 23982 2274 24042 2350
rect 25589 2347 25655 2350
rect 17312 2214 24042 2274
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 23289 2138 23355 2141
rect 9673 2136 14842 2138
rect 9673 2080 9678 2136
rect 9734 2080 14842 2136
rect 9673 2078 14842 2080
rect 17174 2136 23355 2138
rect 17174 2080 23294 2136
rect 23350 2080 23355 2136
rect 17174 2078 23355 2080
rect 9673 2075 9739 2078
rect 1945 2002 2011 2005
rect 14089 2002 14155 2005
rect 1945 2000 14155 2002
rect 1945 1944 1950 2000
rect 2006 1944 14094 2000
rect 14150 1944 14155 2000
rect 1945 1942 14155 1944
rect 14782 2002 14842 2078
rect 23289 2075 23355 2078
rect 15285 2002 15351 2005
rect 14782 2000 15351 2002
rect 14782 1944 15290 2000
rect 15346 1944 15351 2000
rect 14782 1942 15351 1944
rect 1945 1939 2011 1942
rect 14089 1939 14155 1942
rect 15285 1939 15351 1942
rect 17493 2002 17559 2005
rect 24025 2002 24091 2005
rect 17493 2000 24091 2002
rect 17493 1944 17498 2000
rect 17554 1944 24030 2000
rect 24086 1944 24091 2000
rect 17493 1942 24091 1944
rect 17493 1939 17559 1942
rect 24025 1939 24091 1942
rect 3877 1866 3943 1869
rect 8661 1866 8727 1869
rect 21173 1866 21239 1869
rect 3877 1864 8727 1866
rect 3877 1808 3882 1864
rect 3938 1808 8666 1864
rect 8722 1808 8727 1864
rect 3877 1806 8727 1808
rect 3877 1803 3943 1806
rect 8661 1803 8727 1806
rect 8894 1864 21239 1866
rect 8894 1808 21178 1864
rect 21234 1808 21239 1864
rect 8894 1806 21239 1808
rect 4245 1730 4311 1733
rect 8894 1730 8954 1806
rect 21173 1803 21239 1806
rect 4245 1728 8954 1730
rect 4245 1672 4250 1728
rect 4306 1672 8954 1728
rect 4245 1670 8954 1672
rect 10501 1730 10567 1733
rect 24117 1730 24183 1733
rect 10501 1728 24183 1730
rect 10501 1672 10506 1728
rect 10562 1672 24122 1728
rect 24178 1672 24183 1728
rect 10501 1670 24183 1672
rect 4245 1667 4311 1670
rect 10501 1667 10567 1670
rect 24117 1667 24183 1670
rect 4153 1594 4219 1597
rect 8477 1594 8543 1597
rect 4153 1592 8543 1594
rect 4153 1536 4158 1592
rect 4214 1536 8482 1592
rect 8538 1536 8543 1592
rect 4153 1534 8543 1536
rect 4153 1531 4219 1534
rect 8477 1531 8543 1534
rect 8753 1594 8819 1597
rect 20529 1594 20595 1597
rect 8753 1592 20595 1594
rect 8753 1536 8758 1592
rect 8814 1536 20534 1592
rect 20590 1536 20595 1592
rect 8753 1534 20595 1536
rect 8753 1531 8819 1534
rect 20529 1531 20595 1534
rect 0 1458 480 1488
rect 8201 1458 8267 1461
rect 13813 1458 13879 1461
rect 0 1456 8267 1458
rect 0 1400 8206 1456
rect 8262 1400 8267 1456
rect 0 1398 8267 1400
rect 0 1368 480 1398
rect 8201 1395 8267 1398
rect 8342 1456 13879 1458
rect 8342 1400 13818 1456
rect 13874 1400 13879 1456
rect 8342 1398 13879 1400
rect 3785 1322 3851 1325
rect 8342 1322 8402 1398
rect 13813 1395 13879 1398
rect 3785 1320 8402 1322
rect 3785 1264 3790 1320
rect 3846 1264 8402 1320
rect 3785 1262 8402 1264
rect 8477 1322 8543 1325
rect 22461 1322 22527 1325
rect 8477 1320 22527 1322
rect 8477 1264 8482 1320
rect 8538 1264 22466 1320
rect 22522 1264 22527 1320
rect 8477 1262 22527 1264
rect 3785 1259 3851 1262
rect 8477 1259 8543 1262
rect 22461 1259 22527 1262
rect 1117 1186 1183 1189
rect 15377 1186 15443 1189
rect 1117 1184 15443 1186
rect 1117 1128 1122 1184
rect 1178 1128 15382 1184
rect 15438 1128 15443 1184
rect 1117 1126 15443 1128
rect 1117 1123 1183 1126
rect 15377 1123 15443 1126
rect 3417 1050 3483 1053
rect 8477 1050 8543 1053
rect 3417 1048 8543 1050
rect 3417 992 3422 1048
rect 3478 992 8482 1048
rect 8538 992 8543 1048
rect 3417 990 8543 992
rect 3417 987 3483 990
rect 8477 987 8543 990
rect 0 506 480 536
rect 1393 506 1459 509
rect 0 504 1459 506
rect 0 448 1398 504
rect 1454 448 1459 504
rect 0 446 1459 448
rect 0 416 480 446
rect 1393 443 1459 446
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 1716 20768 1780 20772
rect 1716 20712 1730 20768
rect 1730 20712 1780 20768
rect 1716 20708 1780 20712
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 2636 19408 2700 19412
rect 2636 19352 2650 19408
rect 2650 19352 2700 19408
rect 2636 19348 2700 19352
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 1532 18048 1596 18052
rect 1532 17992 1546 18048
rect 1546 17992 1596 18048
rect 1532 17988 1596 17992
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 2268 15872 2332 15876
rect 2268 15816 2282 15872
rect 2282 15816 2332 15872
rect 2268 15812 2332 15816
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 2084 15328 2148 15332
rect 2084 15272 2134 15328
rect 2134 15272 2148 15328
rect 2084 15268 2148 15272
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 9996 12684 10060 12748
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 9996 10100 10060 10164
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 2084 9556 2148 9620
rect 10732 9420 10796 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 10732 6700 10796 6764
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 1716 6292 1780 6356
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 2268 4388 2332 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 1532 3980 1596 4044
rect 2268 3844 2332 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 2636 3708 2700 3772
rect 6132 3708 6196 3772
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 22508 3768 22572 3772
rect 22508 3712 22558 3768
rect 22558 3712 22572 3768
rect 22508 3708 22572 3712
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 1715 20772 1781 20773
rect 1715 20708 1716 20772
rect 1780 20708 1781 20772
rect 1715 20707 1781 20708
rect 1531 18052 1597 18053
rect 1531 17988 1532 18052
rect 1596 17988 1597 18052
rect 1531 17987 1597 17988
rect 1534 4045 1594 17987
rect 1718 6357 1778 20707
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 2635 19412 2701 19413
rect 2635 19348 2636 19412
rect 2700 19348 2701 19412
rect 2635 19347 2701 19348
rect 2267 15876 2333 15877
rect 2267 15812 2268 15876
rect 2332 15812 2333 15876
rect 2267 15811 2333 15812
rect 2083 15332 2149 15333
rect 2083 15268 2084 15332
rect 2148 15268 2149 15332
rect 2083 15267 2149 15268
rect 2086 9621 2146 15267
rect 2083 9620 2149 9621
rect 2083 9556 2084 9620
rect 2148 9556 2149 9620
rect 2083 9555 2149 9556
rect 1715 6356 1781 6357
rect 1715 6292 1716 6356
rect 1780 6292 1781 6356
rect 1715 6291 1781 6292
rect 2270 4453 2330 15811
rect 2267 4452 2333 4453
rect 2267 4388 2268 4452
rect 2332 4388 2333 4452
rect 2267 4387 2333 4388
rect 1531 4044 1597 4045
rect 1531 3980 1532 4044
rect 1596 3980 1597 4044
rect 1531 3979 1597 3980
rect 2270 3909 2330 4387
rect 2267 3908 2333 3909
rect 2267 3844 2268 3908
rect 2332 3844 2333 3908
rect 2267 3843 2333 3844
rect 2638 3773 2698 19347
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9995 12748 10061 12749
rect 9995 12684 9996 12748
rect 10060 12684 10061 12748
rect 9995 12683 10061 12684
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 9998 10165 10058 12683
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9995 10164 10061 10165
rect 9995 10100 9996 10164
rect 10060 10100 10061 10164
rect 9995 10099 10061 10100
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 2635 3772 2701 3773
rect 2635 3708 2636 3772
rect 2700 3708 2701 3772
rect 2635 3707 2701 3708
rect 5610 3296 5931 4320
rect 10277 9280 10597 10304
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 10731 9484 10797 9485
rect 10731 9420 10732 9484
rect 10796 9420 10797 9484
rect 10731 9419 10797 9420
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10734 6765 10794 9419
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 10731 6764 10797 6765
rect 10731 6700 10732 6764
rect 10796 6700 10797 6764
rect 10731 6699 10797 6700
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 6046 3772 6282 3858
rect 6046 3708 6132 3772
rect 6132 3708 6196 3772
rect 6196 3708 6282 3772
rect 6046 3622 6282 3708
rect 22422 3772 22658 3858
rect 22422 3708 22508 3772
rect 22508 3708 22572 3772
rect 22572 3708 22658 3772
rect 22422 3622 22658 3708
<< metal5 >>
rect 6004 3858 22700 3900
rect 6004 3622 6046 3858
rect 6282 3622 22422 3858
rect 22658 3622 22700 3858
rect 6004 3580 22700 3622
use scs8hd_decap_3  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_8
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_41 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_45 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _232_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_48
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_54
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_53
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _207_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_109 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 682 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_140
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_196 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 774 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use scs8hd_conb_1  _208_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_80 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_116
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_124
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_170
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_174
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_9
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_83
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_87
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_100
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_104
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _105_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_221
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_225
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_237
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_9
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_21
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_25
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_47
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _143_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_151
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_204
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_81
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_85
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_161
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_165
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_18
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_22
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_63
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_119
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_136
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_198
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_207
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_248
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _106_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 314 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_253
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_265
timestamp 1586364061
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_273
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_267
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_14
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_53
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 590 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 314 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_264
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_20
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_24
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_nor3_4  _171_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 1234 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 406 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_228
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_248
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 24104 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_252
timestamp 1586364061
transform 1 0 24288 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_259
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_263
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_38
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_116
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_140
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_162
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_235
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 406 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 866 592
use scs8hd_decap_6  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_228
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 9752 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_103
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_157
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_161
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_229
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_241
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_38
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_35
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_50
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_61
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_65
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 1234 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 314 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_123
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_225
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_237
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_248
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_252
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_264
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_50
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_137
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 406 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_209
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_233
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_6  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_110
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 406 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_53
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 1050 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_76
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_26
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 406 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_181
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_54
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_82
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 4324 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_38
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_42
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_122
timestamp 1586364061
transform 1 0 12328 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_134
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_160
timestamp 1586364061
transform 1 0 15824 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_172
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_184
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_155
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_17
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 4508 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_57
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_99
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_103
timestamp 1586364061
transform 1 0 10580 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_127
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_139
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_160
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_172
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_184
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_196
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_208
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_9
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 590 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_43
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_25_50
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_18
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_106
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_17
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_29
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_136
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 590 592
use scs8hd_decap_6  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_60
timestamp 1586364061
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_55
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_6
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_10
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_46
timestamp 1586364061
transform 1 0 5336 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_6
timestamp 1586364061
transform 1 0 1656 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_10
timestamp 1586364061
transform 1 0 2024 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_46
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_14
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_50
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 15566 0 15622 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 16302 0 16358 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 17130 0 17186 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 17958 0 18014 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 18694 0 18750 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 19522 0 19578 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 386 0 442 480 6 bottom_left_grid_pin_13_
port 6 nsew default input
rlabel metal2 s 12346 0 12402 480 6 bottom_right_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 13082 0 13138 480 6 bottom_right_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 13910 0 13966 480 6 bottom_right_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 8298 0 8354 480 6 bottom_right_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 9126 0 9182 480 6 bottom_right_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 9954 0 10010 480 6 bottom_right_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 10690 0 10746 480 6 bottom_right_grid_pin_7_
port 13 nsew default input
rlabel metal2 s 11518 0 11574 480 6 bottom_right_grid_pin_9_
port 14 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal2 s 2778 0 2834 480 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 25134 0 25190 480 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 25870 0 25926 480 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal2 s 26698 0 26754 480 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 data_in
port 51 nsew default input
rlabel metal2 s 14738 0 14794 480 6 enable
port 52 nsew default input
rlabel metal3 s 0 416 480 536 6 left_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 0 26256 480 26376 6 left_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 0 27344 480 27464 6 left_top_grid_pin_15_
port 56 nsew default input
rlabel metal3 s 0 20000 480 20120 6 left_top_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 0 21088 480 21208 6 left_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 22176 480 22296 6 left_top_grid_pin_5_
port 59 nsew default input
rlabel metal3 s 0 23128 480 23248 6 left_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< properties >>
string FIXED_BBOX 0 0 27587 27464
<< end >>
