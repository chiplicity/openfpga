* NGSPICE file created from grid_clb.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfbbp_1 abstract view
.subckt scs8hd_dfbbp_1 CLK D Q QN RESETB SETB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_16 abstract view
.subckt scs8hd_clkbuf_16 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_1 abstract view
.subckt scs8hd_clkbuf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt grid_clb address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] address[7] address[8] address[9] bottom_width_0_height_0__pin_10_ bottom_width_0_height_0__pin_14_
+ bottom_width_0_height_0__pin_2_ bottom_width_0_height_0__pin_6_ clk data_in enable
+ left_width_0_height_0__pin_11_ left_width_0_height_0__pin_3_ left_width_0_height_0__pin_7_
+ reset right_width_0_height_0__pin_13_ right_width_0_height_0__pin_1_ right_width_0_height_0__pin_5_
+ right_width_0_height_0__pin_9_ set top_width_0_height_0__pin_0_ top_width_0_height_0__pin_12_
+ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_8_ vpwr vgnd
XFILLER_79_391 vgnd vpwr scs8hd_decap_12
XFILLER_36_19 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_54_225 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_461 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_77_328 vgnd vpwr scs8hd_decap_12
XFILLER_77_306 vgnd vpwr scs8hd_decap_12
XFILLER_77_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_SLEEPB _518_/Y vgnd vpwr scs8hd_diode_2
XFILLER_73_501 vgnd vpwr scs8hd_decap_12
XFILLER_45_214 vpwr vgnd scs8hd_fill_2
XFILLER_26_41 vgnd vpwr scs8hd_decap_8
XFILLER_33_409 vgnd vpwr scs8hd_decap_4
X_501_ _523_/A _499_/B _501_/Y vgnd vpwr scs8hd_nor2_4
X_432_ _454_/A _429_/X _432_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_442 vpwr vgnd scs8hd_fill_2
X_363_ _328_/X _360_/X _363_/Y vgnd vpwr scs8hd_nor2_4
X_294_ _294_/A _294_/X vgnd vpwr scs8hd_buf_1
XFILLER_42_84 vgnd vpwr scs8hd_decap_6
XFILLER_5_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_328 vpwr vgnd scs8hd_fill_2
XFILLER_76_394 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_269 vgnd vpwr scs8hd_decap_6
XFILLER_44_291 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__304__A _301_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_55_501 vgnd vpwr scs8hd_decap_12
XFILLER_67_383 vpwr vgnd scs8hd_fill_2
XANTENNA__396__D _471_/D vgnd vpwr scs8hd_diode_2
XFILLER_82_342 vgnd vpwr scs8hd_decap_12
XFILLER_70_515 vgnd vpwr scs8hd_fill_1
XFILLER_63_39 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_206 vgnd vpwr scs8hd_decap_8
XFILLER_82_397 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_324 vgnd vpwr scs8hd_decap_12
XFILLER_77_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _546_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_51 vpwr vgnd scs8hd_fill_2
XFILLER_73_353 vpwr vgnd scs8hd_fill_2
XFILLER_73_342 vpwr vgnd scs8hd_fill_2
XFILLER_18_236 vgnd vpwr scs8hd_fill_1
XFILLER_73_397 vpwr vgnd scs8hd_fill_2
X_415_ _509_/A _454_/A vgnd vpwr scs8hd_buf_1
XFILLER_53_50 vgnd vpwr scs8hd_decap_4
X_346_ address[8] _383_/B _320_/C _471_/D _346_/X vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _642_/HI ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_277_ _277_/A _590_/A _277_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_78_80 vgnd vpwr scs8hd_decap_12
XFILLER_68_169 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_501 vgnd vpwr scs8hd_decap_12
XFILLER_49_394 vpwr vgnd scs8hd_fill_2
XFILLER_64_364 vgnd vpwr scs8hd_decap_3
XFILLER_52_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _571_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_401 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_59_103 vpwr vgnd scs8hd_fill_2
XFILLER_59_114 vpwr vgnd scs8hd_fill_2
XFILLER_74_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_27 vgnd vpwr scs8hd_decap_4
XFILLER_67_180 vgnd vpwr scs8hd_decap_3
XFILLER_55_386 vpwr vgnd scs8hd_fill_2
XPHY_702 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_SLEEPB _492_/Y vgnd vpwr scs8hd_diode_2
XPHY_735 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_724 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_713 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_768 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_757 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_746 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_423 vgnd vpwr scs8hd_decap_4
XPHY_779 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_489 vgnd vpwr scs8hd_decap_12
XFILLER_23_75 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ _512_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_78_434 vgnd vpwr scs8hd_decap_12
XANTENNA__598__B _581_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_501 vgnd vpwr scs8hd_decap_12
XFILLER_61_301 vpwr vgnd scs8hd_fill_2
XFILLER_34_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ _469_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_71 vgnd vpwr scs8hd_decap_12
XFILLER_61_345 vpwr vgnd scs8hd_fill_2
XFILLER_61_367 vpwr vgnd scs8hd_fill_2
XFILLER_61_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_329_ _328_/X _322_/X _329_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ _426_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_478 vgnd vpwr scs8hd_decap_8
XANTENNA__301__B _597_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_489 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_301 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_253 vgnd vpwr scs8hd_decap_4
XFILLER_20_264 vgnd vpwr scs8hd_decap_8
XFILLER_69_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_SLEEPB _459_/Y vgnd vpwr scs8hd_diode_2
XFILLER_75_426 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_331 vpwr vgnd scs8hd_fill_2
XFILLER_28_342 vpwr vgnd scs8hd_fill_2
XFILLER_55_150 vgnd vpwr scs8hd_decap_4
XFILLER_16_504 vgnd vpwr scs8hd_decap_12
XFILLER_43_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q
+ _487_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y _624_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_41 vgnd vpwr scs8hd_decap_3
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_378 vpwr vgnd scs8hd_fill_2
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_587 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_576 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_565 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_598 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _617_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q
+ _444_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_452 vgnd vpwr scs8hd_decap_12
XFILLER_59_60 vgnd vpwr scs8hd_fill_1
XANTENNA__402__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_106 vpwr vgnd scs8hd_fill_2
XFILLER_66_448 vpwr vgnd scs8hd_fill_2
XFILLER_19_397 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ _392_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_61_131 vpwr vgnd scs8hd_fill_2
XFILLER_34_345 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ _338_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__312__A _274_/B vgnd vpwr scs8hd_diode_2
XFILLER_57_404 vgnd vpwr scs8hd_decap_3
XFILLER_29_106 vgnd vpwr scs8hd_decap_3
XFILLER_69_297 vpwr vgnd scs8hd_fill_2
XFILLER_57_437 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_470 vgnd vpwr scs8hd_decap_12
XFILLER_25_301 vpwr vgnd scs8hd_fill_2
XFILLER_25_323 vgnd vpwr scs8hd_decap_4
XFILLER_25_367 vgnd vpwr scs8hd_decap_4
XFILLER_80_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_SLEEPB _426_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_164 vgnd vpwr scs8hd_decap_8
XFILLER_71_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_337 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _577_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_466 vgnd vpwr scs8hd_decap_12
XFILLER_48_404 vgnd vpwr scs8hd_fill_1
XFILLER_29_85 vpwr vgnd scs8hd_fill_2
XFILLER_48_437 vgnd vpwr scs8hd_decap_4
XFILLER_48_459 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _285_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_470 vgnd vpwr scs8hd_decap_12
X_594_ _594_/A _594_/B _594_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_73 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _627_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_389 vpwr vgnd scs8hd_fill_2
XFILLER_43_175 vpwr vgnd scs8hd_fill_2
XFILLER_45_84 vpwr vgnd scs8hd_fill_2
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_197 vgnd vpwr scs8hd_decap_4
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_3_293 vgnd vpwr scs8hd_decap_12
XFILLER_66_234 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XFILLER_62_462 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__307__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_SLEEPB _379_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_201 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_57_234 vpwr vgnd scs8hd_fill_2
XFILLER_57_212 vpwr vgnd scs8hd_fill_2
XFILLER_17_109 vpwr vgnd scs8hd_fill_2
XFILLER_72_215 vgnd vpwr scs8hd_decap_12
XFILLER_82_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_31 vpwr vgnd scs8hd_fill_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_407 vpwr vgnd scs8hd_fill_2
XFILLER_36_418 vgnd vpwr scs8hd_decap_8
XFILLER_48_267 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_SLEEPB _513_/Y vgnd vpwr scs8hd_diode_2
X_646_ _646_/HI _646_/LO vgnd vpwr scs8hd_conb_1
XFILLER_63_248 vpwr vgnd scs8hd_fill_2
XFILLER_16_164 vgnd vpwr scs8hd_decap_8
X_577_ _274_/B _574_/X _577_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_292 vpwr vgnd scs8hd_fill_2
XFILLER_72_93 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_385 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_3
XFILLER_39_267 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_54_215 vgnd vpwr scs8hd_decap_4
XFILLER_27_418 vpwr vgnd scs8hd_fill_2
XFILLER_35_473 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vgnd vpwr scs8hd_decap_3
XFILLER_22_167 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_27 vgnd vpwr scs8hd_decap_12
XFILLER_77_318 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__500__A _522_/A vgnd vpwr scs8hd_diode_2
XFILLER_73_513 vgnd vpwr scs8hd_decap_3
XFILLER_18_418 vgnd vpwr scs8hd_fill_1
X_500_ _522_/A _499_/B _500_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_440 vgnd vpwr scs8hd_decap_12
X_431_ _442_/A _429_/X _431_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_64 vgnd vpwr scs8hd_fill_1
XFILLER_53_292 vgnd vpwr scs8hd_decap_8
X_362_ _325_/X _360_/X _362_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_134 vpwr vgnd scs8hd_fill_2
XFILLER_9_127 vpwr vgnd scs8hd_fill_2
X_293_ _278_/X _260_/B _294_/A vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_SLEEPB _480_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__410__A _409_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_248 vgnd vpwr scs8hd_decap_6
X_629_ _629_/A _629_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__304__B _304_/B vgnd vpwr scs8hd_diode_2
XANTENNA__320__A address[8] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_362 vpwr vgnd scs8hd_fill_2
XFILLER_55_513 vgnd vpwr scs8hd_decap_3
XFILLER_82_354 vgnd vpwr scs8hd_decap_12
XFILLER_27_237 vgnd vpwr scs8hd_decap_4
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_137 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_159 vgnd vpwr scs8hd_decap_12
XFILLER_58_340 vpwr vgnd scs8hd_fill_2
XFILLER_37_96 vpwr vgnd scs8hd_fill_2
X_414_ _442_/A _422_/B _414_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_443 vgnd vpwr scs8hd_fill_1
XFILLER_41_240 vpwr vgnd scs8hd_fill_2
X_345_ _515_/D _471_/D vgnd vpwr scs8hd_buf_1
XFILLER_41_262 vgnd vpwr scs8hd_decap_4
XFILLER_41_273 vpwr vgnd scs8hd_fill_2
X_276_ _276_/A _590_/A vgnd vpwr scs8hd_buf_1
XANTENNA__405__A _340_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _312_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_513 vgnd vpwr scs8hd_decap_3
XFILLER_64_343 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_398 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__315__A address[9] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _551_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_70_302 vgnd vpwr scs8hd_fill_1
XFILLER_15_207 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_736 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_725 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_714 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_703 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_769 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_758 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_747 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_32 vpwr vgnd scs8hd_fill_2
XFILLER_7_428 vgnd vpwr scs8hd_decap_12
XFILLER_23_65 vpwr vgnd scs8hd_fill_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_78_446 vgnd vpwr scs8hd_decap_12
XFILLER_65_118 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_513 vgnd vpwr scs8hd_decap_3
XFILLER_73_184 vgnd vpwr scs8hd_decap_12
XFILLER_46_398 vgnd vpwr scs8hd_decap_4
XFILLER_64_83 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_284 vpwr vgnd scs8hd_fill_2
XFILLER_80_93 vgnd vpwr scs8hd_decap_12
X_328_ _509_/A _328_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_259_ _259_/A _239_/A _286_/B _260_/B vgnd vpwr scs8hd_or3_4
XFILLER_6_483 vgnd vpwr scs8hd_decap_12
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_424 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_332 vpwr vgnd scs8hd_fill_2
XFILLER_64_140 vpwr vgnd scs8hd_fill_2
XFILLER_20_210 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_287 vgnd vpwr scs8hd_decap_12
XFILLER_69_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y _615_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_118 vpwr vgnd scs8hd_fill_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _244_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_54 vgnd vpwr scs8hd_decap_6
XFILLER_28_376 vpwr vgnd scs8hd_fill_2
XFILLER_28_387 vpwr vgnd scs8hd_fill_2
XFILLER_28_398 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_70_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_357 vpwr vgnd scs8hd_fill_2
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _624_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_577 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_566 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_599 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_588 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
XFILLER_11_298 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _644_/HI ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_464 vgnd vpwr scs8hd_decap_12
XANTENNA__402__B _404_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_276 vgnd vpwr scs8hd_decap_12
XFILLER_19_343 vpwr vgnd scs8hd_fill_2
XFILLER_46_140 vpwr vgnd scs8hd_fill_2
XFILLER_74_471 vgnd vpwr scs8hd_decap_12
XFILLER_19_376 vgnd vpwr scs8hd_decap_4
XFILLER_34_313 vpwr vgnd scs8hd_fill_2
XFILLER_34_324 vpwr vgnd scs8hd_fill_2
XFILLER_46_184 vgnd vpwr scs8hd_fill_1
XFILLER_34_357 vgnd vpwr scs8hd_decap_8
XFILLER_61_176 vgnd vpwr scs8hd_decap_3
XFILLER_61_165 vgnd vpwr scs8hd_decap_4
XANTENNA__312__B _309_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_57_449 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_482 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_346 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_154 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XANTENNA__503__A _425_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_SLEEPB _388_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_478 vgnd vpwr scs8hd_decap_12
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_416 vgnd vpwr scs8hd_decap_6
XFILLER_63_419 vpwr vgnd scs8hd_fill_2
XFILLER_56_482 vgnd vpwr scs8hd_decap_12
XFILLER_16_324 vgnd vpwr scs8hd_decap_12
XFILLER_45_30 vpwr vgnd scs8hd_fill_2
XFILLER_71_441 vgnd vpwr scs8hd_fill_1
X_593_ _593_/A _594_/B _593_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_346 vgnd vpwr scs8hd_decap_3
XFILLER_43_132 vgnd vpwr scs8hd_decap_3
XFILLER_16_379 vgnd vpwr scs8hd_fill_1
XFILLER_31_316 vpwr vgnd scs8hd_fill_2
XFILLER_43_154 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y _633_/A vgnd vpwr scs8hd_inv_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_327 vpwr vgnd scs8hd_fill_2
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_95 vpwr vgnd scs8hd_fill_2
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__413__A _413_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_66_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_416 vpwr vgnd scs8hd_fill_2
XFILLER_66_224 vpwr vgnd scs8hd_fill_2
XFILLER_19_140 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XFILLER_34_121 vgnd vpwr scs8hd_decap_8
XFILLER_62_474 vgnd vpwr scs8hd_decap_12
XFILLER_34_165 vgnd vpwr scs8hd_decap_8
XFILLER_34_187 vpwr vgnd scs8hd_fill_2
XFILLER_30_382 vpwr vgnd scs8hd_fill_2
XANTENNA__323__A _314_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_72_249 vpwr vgnd scs8hd_fill_2
XFILLER_53_441 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_SLEEPB _349_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_40_102 vgnd vpwr scs8hd_decap_4
XFILLER_40_113 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _641_/HI ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_382 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _285_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _563_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_54 vgnd vpwr scs8hd_fill_1
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_48_224 vgnd vpwr scs8hd_decap_3
XFILLER_48_257 vgnd vpwr scs8hd_fill_1
XFILLER_63_216 vgnd vpwr scs8hd_fill_1
XFILLER_48_279 vgnd vpwr scs8hd_decap_4
X_645_ _645_/HI _645_/LO vgnd vpwr scs8hd_conb_1
XFILLER_56_290 vgnd vpwr scs8hd_decap_8
XFILLER_16_154 vgnd vpwr scs8hd_fill_1
X_576_ _270_/B _574_/X _576_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__408__A address[6] vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_decap_3
XFILLER_12_382 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_249 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__318__A enable vgnd vpwr scs8hd_diode_2
XFILLER_35_485 vgnd vpwr scs8hd_decap_3
XFILLER_10_308 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _577_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_157 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_2_507 vgnd vpwr scs8hd_decap_8
XFILLER_77_39 vgnd vpwr scs8hd_decap_12
XANTENNA__500__B _499_/B vgnd vpwr scs8hd_diode_2
XFILLER_45_205 vgnd vpwr scs8hd_decap_4
XFILLER_26_452 vgnd vpwr scs8hd_decap_6
X_430_ _441_/A _429_/X _430_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_271 vpwr vgnd scs8hd_fill_2
X_361_ _314_/X _360_/X _361_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__228__A _578_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_179 vgnd vpwr scs8hd_decap_4
XFILLER_13_168 vgnd vpwr scs8hd_fill_1
X_292_ _277_/A _594_/A _292_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_190 vpwr vgnd scs8hd_fill_2
XFILLER_42_64 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_367 vgnd vpwr scs8hd_decap_12
XFILLER_68_308 vgnd vpwr scs8hd_fill_1
XFILLER_76_330 vgnd vpwr scs8hd_decap_6
XFILLER_36_205 vgnd vpwr scs8hd_fill_1
X_628_ _628_/A _628_/Y vgnd vpwr scs8hd_inv_8
X_559_ _585_/A _561_/B _559_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_73_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_183 vpwr vgnd scs8hd_fill_2
XANTENNA__601__A _575_/A vgnd vpwr scs8hd_diode_2
XANTENNA__320__B _383_/B vgnd vpwr scs8hd_diode_2
XFILLER_67_341 vpwr vgnd scs8hd_fill_2
XFILLER_82_311 vgnd vpwr scs8hd_decap_12
XFILLER_27_227 vgnd vpwr scs8hd_decap_3
XFILLER_27_249 vgnd vpwr scs8hd_decap_3
XFILLER_82_366 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _592_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_271 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_285 vgnd vpwr scs8hd_decap_8
XFILLER_50_263 vpwr vgnd scs8hd_fill_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_127 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_337 vgnd vpwr scs8hd_decap_12
XANTENNA__511__A _522_/A vgnd vpwr scs8hd_diode_2
XANTENNA__230__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_20 vpwr vgnd scs8hd_fill_2
XFILLER_73_322 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_75 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_413_ _413_/A _442_/A vgnd vpwr scs8hd_buf_1
XFILLER_26_271 vpwr vgnd scs8hd_fill_2
XFILLER_41_230 vpwr vgnd scs8hd_fill_2
XFILLER_53_96 vpwr vgnd scs8hd_fill_2
X_344_ _395_/A _344_/B _344_/Y vgnd vpwr scs8hd_nor2_4
X_275_ _242_/A _302_/B _276_/A vgnd vpwr scs8hd_or2_4
XANTENNA__405__B _405_/B vgnd vpwr scs8hd_diode_2
XANTENNA__421__A _523_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_93 vgnd vpwr scs8hd_decap_12
XFILLER_68_105 vgnd vpwr scs8hd_decap_8
XFILLER_49_352 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _583_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_447 vgnd vpwr scs8hd_decap_8
XFILLER_32_285 vpwr vgnd scs8hd_fill_2
XANTENNA__331__A _510_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_149 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_300 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_344 vgnd vpwr scs8hd_decap_3
XFILLER_70_325 vpwr vgnd scs8hd_fill_2
XFILLER_15_219 vpwr vgnd scs8hd_fill_2
XPHY_726 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_715 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_704 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_759 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_748 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_737 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_252 vpwr vgnd scs8hd_fill_2
XFILLER_23_274 vpwr vgnd scs8hd_fill_2
XFILLER_23_55 vpwr vgnd scs8hd_fill_2
XANTENNA__506__A _505_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XANTENNA__241__A _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_48_85 vgnd vpwr scs8hd_fill_1
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_325 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_46_388 vgnd vpwr scs8hd_decap_8
XFILLER_73_196 vgnd vpwr scs8hd_decap_12
XFILLER_61_358 vpwr vgnd scs8hd_fill_2
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XANTENNA__416__A _454_/A vgnd vpwr scs8hd_diode_2
X_327_ _327_/A _509_/A vgnd vpwr scs8hd_buf_1
X_258_ address[2] _259_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_495 vgnd vpwr scs8hd_decap_12
XFILLER_69_436 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _566_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _596_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_160 vgnd vpwr scs8hd_decap_4
XFILLER_64_152 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_185 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_369 vpwr vgnd scs8hd_fill_2
XFILLER_52_347 vgnd vpwr scs8hd_decap_3
XFILLER_60_380 vpwr vgnd scs8hd_fill_2
XANTENNA__326__A _325_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_299 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_75_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_6
XFILLER_28_322 vpwr vgnd scs8hd_fill_2
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
XFILLER_43_314 vpwr vgnd scs8hd_fill_2
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_336 vpwr vgnd scs8hd_fill_2
XFILLER_70_166 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_54 vgnd vpwr scs8hd_decap_8
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_578 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_211 vgnd vpwr scs8hd_fill_1
XFILLER_11_200 vpwr vgnd scs8hd_fill_2
XFILLER_34_65 vpwr vgnd scs8hd_fill_2
XANTENNA__236__A _249_/A vgnd vpwr scs8hd_diode_2
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_567 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_589 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_204 vgnd vpwr scs8hd_decap_12
XFILLER_50_64 vgnd vpwr scs8hd_decap_4
XFILLER_50_97 vgnd vpwr scs8hd_decap_6
XFILLER_59_62 vpwr vgnd scs8hd_fill_2
XFILLER_59_51 vgnd vpwr scs8hd_decap_3
XFILLER_3_476 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_66_428 vgnd vpwr scs8hd_decap_8
XFILLER_78_288 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_322 vgnd vpwr scs8hd_decap_3
XFILLER_74_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_152 vgnd vpwr scs8hd_fill_1
XFILLER_46_163 vgnd vpwr scs8hd_decap_6
XFILLER_61_144 vpwr vgnd scs8hd_fill_2
XFILLER_46_196 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_42_391 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_233 vpwr vgnd scs8hd_fill_2
XFILLER_69_222 vpwr vgnd scs8hd_fill_2
XFILLER_69_277 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _603_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_163 vgnd vpwr scs8hd_decap_6
XFILLER_52_122 vpwr vgnd scs8hd_fill_2
XFILLER_25_358 vpwr vgnd scs8hd_fill_2
XFILLER_40_328 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__503__B _495_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_435 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_43 vpwr vgnd scs8hd_fill_2
XFILLER_75_236 vgnd vpwr scs8hd_decap_3
XFILLER_75_258 vpwr vgnd scs8hd_fill_2
XFILLER_56_450 vpwr vgnd scs8hd_fill_2
X_592_ _592_/A _594_/B _592_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_303 vpwr vgnd scs8hd_fill_2
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_43_100 vpwr vgnd scs8hd_fill_2
XFILLER_56_494 vgnd vpwr scs8hd_decap_12
XFILLER_31_306 vgnd vpwr scs8hd_fill_1
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_30 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_SLEEPB _341_/Y vgnd vpwr scs8hd_diode_2
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _540_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_428 vgnd vpwr scs8hd_decap_3
XFILLER_54_409 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_144 vpwr vgnd scs8hd_fill_2
XFILLER_62_486 vgnd vpwr scs8hd_decap_12
XFILLER_22_328 vpwr vgnd scs8hd_fill_2
XANTENNA__604__A _604_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__323__B _322_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _561_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_269 vpwr vgnd scs8hd_fill_2
XFILLER_57_258 vgnd vpwr scs8hd_decap_6
XFILLER_65_291 vpwr vgnd scs8hd_fill_2
XFILLER_53_431 vpwr vgnd scs8hd_fill_2
XFILLER_13_317 vpwr vgnd scs8hd_fill_2
XFILLER_25_199 vpwr vgnd scs8hd_fill_2
XFILLER_40_147 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__514__A _425_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_88 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_56_41 vpwr vgnd scs8hd_fill_2
X_644_ _644_/HI _644_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_461 vpwr vgnd scs8hd_fill_2
X_575_ _575_/A _574_/X _575_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_161 vgnd vpwr scs8hd_decap_3
XPHY_150 vgnd vpwr scs8hd_decap_3
XFILLER_31_136 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__424__A _447_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q
+ _463_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_501 vgnd vpwr scs8hd_decap_12
XFILLER_39_225 vgnd vpwr scs8hd_decap_6
XFILLER_39_236 vpwr vgnd scs8hd_fill_2
XFILLER_82_515 vgnd vpwr scs8hd_fill_1
XFILLER_54_206 vgnd vpwr scs8hd_decap_8
XFILLER_47_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_SLEEPB _446_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q
+ _414_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__318__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__334__A _522_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q
+ _363_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_409 vgnd vpwr scs8hd_fill_1
XFILLER_26_11 vgnd vpwr scs8hd_decap_3
XFILLER_38_291 vgnd vpwr scs8hd_fill_1
XANTENNA__509__A _509_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_261 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_26_88 vgnd vpwr scs8hd_fill_1
X_360_ _367_/B _360_/X vgnd vpwr scs8hd_buf_1
XFILLER_41_412 vpwr vgnd scs8hd_fill_2
XFILLER_41_423 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vpwr vgnd scs8hd_fill_2
XFILLER_41_456 vgnd vpwr scs8hd_decap_3
XFILLER_41_467 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_41_478 vpwr vgnd scs8hd_fill_2
XFILLER_41_489 vgnd vpwr scs8hd_decap_12
XFILLER_42_43 vgnd vpwr scs8hd_decap_4
X_291_ _291_/A _594_/A vgnd vpwr scs8hd_buf_1
XFILLER_42_54 vgnd vpwr scs8hd_decap_4
XANTENNA__244__A _257_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _558_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_379 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_67_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_49_501 vgnd vpwr scs8hd_decap_12
XFILLER_67_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_627_ _627_/A _627_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__419__A _522_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_464 vpwr vgnd scs8hd_fill_2
XFILLER_44_250 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_475 vpwr vgnd scs8hd_fill_2
X_558_ _584_/A _561_/B _558_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_434 vpwr vgnd scs8hd_fill_2
X_489_ _522_/A _490_/B _489_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_191 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_195 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _608_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_309 vpwr vgnd scs8hd_fill_2
XANTENNA__601__B _600_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_SLEEPB _404_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__320__C _320_/C vgnd vpwr scs8hd_diode_2
XFILLER_67_320 vpwr vgnd scs8hd_fill_2
XFILLER_27_206 vpwr vgnd scs8hd_fill_2
XFILLER_82_323 vgnd vpwr scs8hd_decap_12
XANTENNA__329__A _328_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_401 vpwr vgnd scs8hd_fill_2
XFILLER_23_423 vpwr vgnd scs8hd_fill_2
XFILLER_35_283 vpwr vgnd scs8hd_fill_2
XFILLER_23_456 vpwr vgnd scs8hd_fill_2
XFILLER_23_489 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__511__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_349 vgnd vpwr scs8hd_decap_12
XFILLER_73_301 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_37_32 vpwr vgnd scs8hd_fill_2
XFILLER_73_334 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_65 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
X_412_ _441_/A _422_/B _412_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_423 vgnd vpwr scs8hd_fill_1
XFILLER_14_412 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_31 vgnd vpwr scs8hd_fill_1
XFILLER_53_75 vpwr vgnd scs8hd_fill_2
X_343_ _425_/A _395_/A vgnd vpwr scs8hd_buf_1
X_274_ _259_/A _274_/B _302_/B vgnd vpwr scs8hd_or2_4
XFILLER_41_286 vpwr vgnd scs8hd_fill_2
XFILLER_41_297 vpwr vgnd scs8hd_fill_2
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_68_139 vgnd vpwr scs8hd_fill_1
XFILLER_49_342 vpwr vgnd scs8hd_fill_2
XFILLER_49_364 vpwr vgnd scs8hd_fill_2
XFILLER_64_356 vgnd vpwr scs8hd_decap_8
XFILLER_52_507 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_261 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_SLEEPB _366_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_437 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _312_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__612__A _612_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_128 vpwr vgnd scs8hd_fill_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_67_150 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_515 vgnd vpwr scs8hd_fill_1
XFILLER_67_172 vgnd vpwr scs8hd_decap_8
XFILLER_67_161 vpwr vgnd scs8hd_fill_2
XFILLER_55_323 vpwr vgnd scs8hd_fill_2
XFILLER_55_367 vgnd vpwr scs8hd_decap_4
XFILLER_70_359 vgnd vpwr scs8hd_decap_8
XFILLER_70_348 vpwr vgnd scs8hd_fill_2
XPHY_727 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_716 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_705 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_749 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_738 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_242 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_23 vgnd vpwr scs8hd_decap_3
XFILLER_23_297 vpwr vgnd scs8hd_fill_2
XFILLER_23_78 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_SLEEPB _500_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__522__A _522_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__241__B _241_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_459 vgnd vpwr scs8hd_decap_12
XFILLER_48_42 vgnd vpwr scs8hd_decap_4
XFILLER_58_183 vgnd vpwr scs8hd_decap_4
XFILLER_58_194 vgnd vpwr scs8hd_fill_1
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__416__B _422_/B vgnd vpwr scs8hd_diode_2
X_326_ _325_/X _322_/X _326_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_257_ _257_/A _585_/A _257_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__432__A _454_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_404 vgnd vpwr scs8hd_decap_3
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_326 vgnd vpwr scs8hd_decap_8
XFILLER_37_378 vpwr vgnd scs8hd_fill_2
XFILLER_37_389 vpwr vgnd scs8hd_fill_2
XFILLER_52_337 vgnd vpwr scs8hd_fill_1
XANTENNA__607__A _607_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _640_/HI ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_60_392 vgnd vpwr scs8hd_fill_1
XANTENNA__326__B _322_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__342__A _302_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ _524_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_301 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_SLEEPB _467_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_175 vpwr vgnd scs8hd_fill_2
XFILLER_70_178 vgnd vpwr scs8hd_decap_12
XANTENNA__517__A _517_/A vgnd vpwr scs8hd_diode_2
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_381 vpwr vgnd scs8hd_fill_2
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_568 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ _481_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_579 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_216 vgnd vpwr scs8hd_decap_12
XFILLER_50_43 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_50_87 vgnd vpwr scs8hd_decap_4
XANTENNA__252__A _282_/C vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y _621_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_75_62 vgnd vpwr scs8hd_decap_12
XFILLER_75_51 vgnd vpwr scs8hd_decap_8
XFILLER_74_495 vgnd vpwr scs8hd_decap_12
XFILLER_61_123 vgnd vpwr scs8hd_fill_1
XFILLER_34_337 vpwr vgnd scs8hd_fill_2
XANTENNA__427__A _409_/A vgnd vpwr scs8hd_diode_2
X_309_ _308_/X _309_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _541_/Y vgnd vpwr scs8hd_diode_2
XFILLER_69_256 vpwr vgnd scs8hd_fill_2
XFILLER_57_418 vgnd vpwr scs8hd_decap_3
XFILLER_65_451 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_80_410 vgnd vpwr scs8hd_decap_12
XFILLER_65_462 vpwr vgnd scs8hd_fill_2
XFILLER_25_315 vpwr vgnd scs8hd_fill_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
XFILLER_37_197 vgnd vpwr scs8hd_decap_6
XANTENNA__337__A _523_/A vgnd vpwr scs8hd_diode_2
XFILLER_52_189 vgnd vpwr scs8hd_decap_4
XFILLER_40_318 vgnd vpwr scs8hd_fill_1
XFILLER_33_392 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q
+ _499_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_SLEEPB _434_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ _456_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_447 vgnd vpwr scs8hd_decap_12
XFILLER_29_66 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_462 vpwr vgnd scs8hd_fill_2
X_591_ _591_/A _594_/B _591_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_123 vpwr vgnd scs8hd_fill_2
XFILLER_45_54 vgnd vpwr scs8hd_decap_4
XFILLER_71_454 vpwr vgnd scs8hd_fill_2
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__247__A _247_/A vgnd vpwr scs8hd_diode_2
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_392 vgnd vpwr scs8hd_decap_3
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ _404_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_61_75 vpwr vgnd scs8hd_fill_2
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _531_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ _355_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_66_248 vpwr vgnd scs8hd_fill_2
XFILLER_47_451 vpwr vgnd scs8hd_fill_2
XFILLER_47_462 vpwr vgnd scs8hd_fill_2
XFILLER_62_421 vgnd vpwr scs8hd_decap_8
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_498 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_351 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__620__A _620_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _533_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_421 vpwr vgnd scs8hd_fill_2
XFILLER_53_410 vpwr vgnd scs8hd_fill_2
XFILLER_80_251 vgnd vpwr scs8hd_decap_12
XFILLER_53_465 vpwr vgnd scs8hd_fill_2
XFILLER_53_454 vpwr vgnd scs8hd_fill_2
XFILLER_25_134 vgnd vpwr scs8hd_decap_3
XFILLER_53_487 vgnd vpwr scs8hd_fill_1
XFILLER_25_189 vgnd vpwr scs8hd_decap_3
XFILLER_21_362 vpwr vgnd scs8hd_fill_2
XFILLER_21_395 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__514__B _505_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XANTENNA__530__A _582_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_64 vgnd vpwr scs8hd_decap_4
X_643_ _643_/HI _643_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_574_ _573_/X _574_/X vgnd vpwr scs8hd_buf_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y _616_/A vgnd vpwr scs8hd_buf_1
XFILLER_71_273 vpwr vgnd scs8hd_fill_2
XPHY_151 vgnd vpwr scs8hd_decap_3
XPHY_140 vgnd vpwr scs8hd_decap_3
XPHY_162 vgnd vpwr scs8hd_decap_3
XFILLER_8_300 vgnd vpwr scs8hd_decap_12
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_SLEEPB _521_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__424__B _411_/A vgnd vpwr scs8hd_diode_2
XANTENNA__440__A _448_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_513 vgnd vpwr scs8hd_decap_3
XFILLER_39_204 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_229 vgnd vpwr scs8hd_decap_4
XFILLER_47_270 vgnd vpwr scs8hd_decap_4
XFILLER_35_443 vpwr vgnd scs8hd_fill_2
XFILLER_50_457 vgnd vpwr scs8hd_fill_1
XFILLER_50_468 vgnd vpwr scs8hd_decap_12
XANTENNA__615__A _615_/A vgnd vpwr scs8hd_diode_2
XANTENNA__350__A _325_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_45_218 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_23 vgnd vpwr scs8hd_decap_8
XFILLER_38_281 vpwr vgnd scs8hd_fill_2
XANTENNA__509__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_67 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_13_126 vpwr vgnd scs8hd_fill_2
X_290_ _278_/X _330_/A _291_/A vgnd vpwr scs8hd_or2_4
XFILLER_41_446 vgnd vpwr scs8hd_decap_4
XANTENNA__525__A _425_/A vgnd vpwr scs8hd_diode_2
XANTENNA__244__B _582_/A vgnd vpwr scs8hd_diode_2
XANTENNA__260__A _242_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_49_513 vgnd vpwr scs8hd_decap_3
XFILLER_76_343 vgnd vpwr scs8hd_decap_6
XFILLER_76_321 vgnd vpwr scs8hd_decap_3
XFILLER_67_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_398 vgnd vpwr scs8hd_decap_12
XFILLER_36_229 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_626_ _626_/A _626_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_432 vpwr vgnd scs8hd_fill_2
XFILLER_44_240 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_487 vgnd vpwr scs8hd_fill_1
XFILLER_32_424 vgnd vpwr scs8hd_decap_4
X_557_ _583_/A _561_/B _557_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_457 vgnd vpwr scs8hd_fill_1
XFILLER_44_295 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_488_ _510_/A _490_/B _488_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__435__A _457_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__320__D _409_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_335 vgnd vpwr scs8hd_decap_6
XFILLER_67_398 vgnd vpwr scs8hd_decap_4
XANTENNA__329__B _322_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_240 vpwr vgnd scs8hd_fill_2
XANTENNA__345__A _515_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_321 vpwr vgnd scs8hd_fill_2
XFILLER_58_365 vgnd vpwr scs8hd_decap_12
XFILLER_58_354 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_37_55 vpwr vgnd scs8hd_fill_2
XFILLER_73_357 vpwr vgnd scs8hd_fill_2
XFILLER_37_88 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
X_411_ _411_/A _422_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _619_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_251 vgnd vpwr scs8hd_fill_1
XFILLER_53_54 vgnd vpwr scs8hd_fill_1
XFILLER_53_43 vpwr vgnd scs8hd_fill_2
XFILLER_14_446 vgnd vpwr scs8hd_decap_12
XFILLER_14_435 vpwr vgnd scs8hd_fill_2
X_342_ _302_/B _425_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_254 vpwr vgnd scs8hd_fill_2
X_273_ _277_/A _589_/A _273_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__255__A _242_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_490 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_321 vgnd vpwr scs8hd_decap_4
XFILLER_49_398 vpwr vgnd scs8hd_fill_2
X_609_ _609_/A _609_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_284 vpwr vgnd scs8hd_fill_2
XFILLER_32_232 vgnd vpwr scs8hd_decap_3
XFILLER_20_405 vgnd vpwr scs8hd_decap_12
XFILLER_32_254 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vpwr vgnd scs8hd_fill_2
XFILLER_32_298 vpwr vgnd scs8hd_fill_2
XFILLER_59_118 vpwr vgnd scs8hd_fill_2
XFILLER_59_107 vpwr vgnd scs8hd_fill_2
XFILLER_67_184 vgnd vpwr scs8hd_decap_12
XFILLER_82_187 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_717 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_706 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_739 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_728 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_287 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__522__B _523_/B vgnd vpwr scs8hd_diode_2
XANTENNA__241__C _286_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_3
XFILLER_58_140 vgnd vpwr scs8hd_decap_12
XFILLER_73_110 vgnd vpwr scs8hd_decap_12
XFILLER_46_324 vgnd vpwr scs8hd_decap_12
XFILLER_46_346 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_decap_3
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
X_325_ _413_/A _325_/X vgnd vpwr scs8hd_buf_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _585_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ _492_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_256_ _255_/X _585_/A vgnd vpwr scs8hd_buf_1
XANTENNA__432__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_69_416 vpwr vgnd scs8hd_fill_2
XFILLER_69_449 vpwr vgnd scs8hd_fill_2
XFILLER_37_302 vgnd vpwr scs8hd_fill_1
XFILLER_49_184 vpwr vgnd scs8hd_fill_2
XFILLER_49_195 vpwr vgnd scs8hd_fill_2
XFILLER_64_154 vpwr vgnd scs8hd_fill_2
XFILLER_52_305 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__623__A _623_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_132 vpwr vgnd scs8hd_fill_2
XFILLER_28_335 vgnd vpwr scs8hd_fill_1
XFILLER_28_346 vgnd vpwr scs8hd_decap_4
XFILLER_55_198 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_89 vgnd vpwr scs8hd_decap_3
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_569 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XFILLER_11_235 vgnd vpwr scs8hd_decap_8
XFILLER_7_228 vgnd vpwr scs8hd_decap_12
XANTENNA__533__A _585_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_77 vpwr vgnd scs8hd_fill_2
XANTENNA__252__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_78_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_86 vpwr vgnd scs8hd_fill_2
XFILLER_59_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_302 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_75_74 vgnd vpwr scs8hd_decap_12
XFILLER_46_187 vpwr vgnd scs8hd_fill_2
XANTENNA__427__B _382_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_382 vpwr vgnd scs8hd_fill_2
X_308_ _599_/A _231_/X _308_/X vgnd vpwr scs8hd_or2_4
XANTENNA__443__A _454_/A vgnd vpwr scs8hd_diode_2
X_239_ _239_/A _241_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _295_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_4
XFILLER_37_110 vpwr vgnd scs8hd_fill_2
XFILLER_80_422 vgnd vpwr scs8hd_decap_12
XFILLER_25_338 vpwr vgnd scs8hd_fill_2
XANTENNA__618__A _618_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_308 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_360 vgnd vpwr scs8hd_decap_6
XFILLER_33_371 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__353__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_36 vgnd vpwr scs8hd_fill_1
XFILLER_20_58 vgnd vpwr scs8hd_decap_3
XFILLER_0_404 vgnd vpwr scs8hd_decap_12
XFILLER_0_459 vgnd vpwr scs8hd_decap_6
XFILLER_29_89 vpwr vgnd scs8hd_fill_2
X_590_ _590_/A _594_/B _590_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_28_165 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__528__A _527_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_176 vpwr vgnd scs8hd_fill_2
XFILLER_71_444 vgnd vpwr scs8hd_fill_1
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_45_77 vpwr vgnd scs8hd_fill_2
XFILLER_45_88 vgnd vpwr scs8hd_decap_4
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _633_/Y vgnd vpwr scs8hd_diode_2
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_54 vgnd vpwr scs8hd_decap_4
XFILLER_8_515 vgnd vpwr scs8hd_fill_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__263__A _259_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_290 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vpwr vgnd scs8hd_fill_2
XFILLER_81_208 vgnd vpwr scs8hd_decap_12
XANTENNA__438__A _385_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_157 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_382 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_clkbuf_0_clk_A clk vgnd vpwr scs8hd_diode_2
XFILLER_30_363 vpwr vgnd scs8hd_fill_2
XFILLER_30_396 vgnd vpwr scs8hd_fill_1
XFILLER_57_216 vpwr vgnd scs8hd_fill_2
XFILLER_57_205 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_57_238 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_400 vgnd vpwr scs8hd_decap_3
XANTENNA__348__A _356_/B vgnd vpwr scs8hd_diode_2
XFILLER_80_263 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_46 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__530__B _529_/X vgnd vpwr scs8hd_diode_2
XFILLER_63_219 vpwr vgnd scs8hd_fill_2
X_642_ _642_/HI _642_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XFILLER_29_485 vgnd vpwr scs8hd_decap_3
XANTENNA__258__A address[2] vgnd vpwr scs8hd_diode_2
X_573_ _599_/A _552_/X _573_/X vgnd vpwr scs8hd_or2_4
XFILLER_71_252 vgnd vpwr scs8hd_decap_4
XFILLER_31_105 vpwr vgnd scs8hd_fill_2
XPHY_152 vgnd vpwr scs8hd_decap_3
XFILLER_71_296 vgnd vpwr scs8hd_decap_6
XPHY_141 vgnd vpwr scs8hd_decap_3
XPHY_130 vgnd vpwr scs8hd_decap_3
XFILLER_24_190 vpwr vgnd scs8hd_fill_2
XFILLER_31_149 vpwr vgnd scs8hd_fill_2
XPHY_163 vgnd vpwr scs8hd_decap_3
XFILLER_8_312 vgnd vpwr scs8hd_decap_12
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_396 vgnd vpwr scs8hd_fill_1
XFILLER_12_374 vpwr vgnd scs8hd_fill_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_330 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_477 vgnd vpwr scs8hd_decap_8
XFILLER_62_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_447 vpwr vgnd scs8hd_fill_2
XFILLER_50_436 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_193 vgnd vpwr scs8hd_decap_4
XANTENNA__631__A _631_/A vgnd vpwr scs8hd_diode_2
XANTENNA__350__B _348_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_12 vgnd vpwr scs8hd_decap_8
XFILLER_42_23 vgnd vpwr scs8hd_decap_8
XANTENNA__525__B _517_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_78 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__541__A _593_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__260__B _260_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_300 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_86 vgnd vpwr scs8hd_decap_12
XFILLER_36_208 vgnd vpwr scs8hd_decap_6
XFILLER_29_271 vpwr vgnd scs8hd_fill_2
X_625_ _625_/A _625_/Y vgnd vpwr scs8hd_inv_8
X_556_ _582_/A _561_/B _556_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_263 vgnd vpwr scs8hd_decap_12
XFILLER_32_469 vgnd vpwr scs8hd_decap_8
X_487_ _509_/A _490_/B _487_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__435__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_171 vgnd vpwr scs8hd_decap_3
XFILLER_40_491 vgnd vpwr scs8hd_decap_12
XANTENNA__451__A _451_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__626__A _626_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_296 vpwr vgnd scs8hd_fill_2
XFILLER_50_244 vpwr vgnd scs8hd_fill_2
XFILLER_23_469 vpwr vgnd scs8hd_fill_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__361__A _314_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_333 vgnd vpwr scs8hd_decap_3
XFILLER_58_311 vgnd vpwr scs8hd_decap_6
XFILLER_58_344 vpwr vgnd scs8hd_fill_2
XFILLER_58_377 vgnd vpwr scs8hd_decap_3
XFILLER_37_45 vgnd vpwr scs8hd_decap_4
X_410_ _409_/X _411_/A vgnd vpwr scs8hd_buf_1
XFILLER_81_391 vgnd vpwr scs8hd_decap_12
X_341_ _340_/X _344_/B _341_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__536__A _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_285 vgnd vpwr scs8hd_decap_3
XFILLER_26_296 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_272_ _271_/X _589_/A vgnd vpwr scs8hd_buf_1
XANTENNA__255__B _330_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA__271__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_141 vgnd vpwr scs8hd_decap_12
XFILLER_49_377 vgnd vpwr scs8hd_decap_3
XFILLER_64_369 vgnd vpwr scs8hd_decap_4
X_608_ _608_/A _608_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__446__A _457_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_274 vpwr vgnd scs8hd_fill_2
XFILLER_32_200 vpwr vgnd scs8hd_fill_2
X_539_ _591_/A _542_/B _539_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_244 vgnd vpwr scs8hd_decap_8
XFILLER_20_417 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_440 vgnd vpwr scs8hd_decap_12
XFILLER_71_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_67_130 vgnd vpwr scs8hd_decap_4
XFILLER_67_196 vgnd vpwr scs8hd_decap_12
XFILLER_55_358 vpwr vgnd scs8hd_fill_2
XFILLER_70_306 vpwr vgnd scs8hd_fill_2
XFILLER_82_199 vgnd vpwr scs8hd_decap_12
XPHY_718 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_707 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_200 vpwr vgnd scs8hd_fill_2
XANTENNA__356__A _395_/A vgnd vpwr scs8hd_diode_2
XPHY_729 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_428 vgnd vpwr scs8hd_decap_12
XFILLER_23_47 vpwr vgnd scs8hd_fill_2
XFILLER_23_69 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _625_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_66 vgnd vpwr scs8hd_decap_8
XFILLER_58_152 vgnd vpwr scs8hd_fill_1
XFILLER_48_77 vpwr vgnd scs8hd_fill_2
XFILLER_48_88 vgnd vpwr scs8hd_decap_4
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_61_317 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_328 vpwr vgnd scs8hd_fill_2
XFILLER_54_391 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__266__A _257_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_288 vgnd vpwr scs8hd_decap_4
XFILLER_14_266 vpwr vgnd scs8hd_fill_2
X_324_ _324_/A _413_/A vgnd vpwr scs8hd_buf_1
X_255_ _242_/A _330_/A _255_/X vgnd vpwr scs8hd_or2_4
XFILLER_6_410 vgnd vpwr scs8hd_decap_12
XFILLER_10_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _257_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_69_428 vgnd vpwr scs8hd_fill_1
XFILLER_49_152 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_347 vpwr vgnd scs8hd_fill_2
XFILLER_37_358 vpwr vgnd scs8hd_fill_2
XFILLER_64_144 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_225 vgnd vpwr scs8hd_decap_12
XFILLER_9_281 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_306 vgnd vpwr scs8hd_decap_8
XFILLER_34_46 vgnd vpwr scs8hd_decap_4
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_214 vpwr vgnd scs8hd_fill_2
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_394 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__533__B _529_/X vgnd vpwr scs8hd_diode_2
XFILLER_59_32 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_409 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_347 vgnd vpwr scs8hd_decap_6
XFILLER_46_133 vgnd vpwr scs8hd_decap_4
XFILLER_75_86 vgnd vpwr scs8hd_decap_12
XFILLER_19_358 vpwr vgnd scs8hd_fill_2
XFILLER_46_144 vgnd vpwr scs8hd_decap_8
XFILLER_61_114 vpwr vgnd scs8hd_fill_2
XFILLER_27_380 vpwr vgnd scs8hd_fill_2
XFILLER_34_317 vpwr vgnd scs8hd_fill_2
XFILLER_34_328 vpwr vgnd scs8hd_fill_2
XFILLER_46_199 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__427__C _409_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_SLEEPB _391_/Y vgnd vpwr scs8hd_diode_2
X_307_ address[4] _599_/A vgnd vpwr scs8hd_inv_8
XANTENNA__443__B _445_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_280 vgnd vpwr scs8hd_decap_12
X_238_ address[1] _239_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_100 vgnd vpwr scs8hd_decap_3
XFILLER_37_144 vpwr vgnd scs8hd_fill_2
XFILLER_37_155 vpwr vgnd scs8hd_fill_2
XFILLER_80_434 vgnd vpwr scs8hd_decap_12
XFILLER_21_501 vgnd vpwr scs8hd_decap_12
XFILLER_33_383 vpwr vgnd scs8hd_fill_2
XANTENNA__634__A _634_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__353__B _348_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_416 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XFILLER_75_228 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_144 vpwr vgnd scs8hd_fill_2
XFILLER_71_423 vpwr vgnd scs8hd_fill_2
XFILLER_71_401 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_114 vpwr vgnd scs8hd_fill_2
XFILLER_45_23 vgnd vpwr scs8hd_fill_1
XFILLER_45_45 vgnd vpwr scs8hd_decap_3
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XFILLER_71_489 vgnd vpwr scs8hd_decap_12
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_180 vgnd vpwr scs8hd_fill_1
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__544__A _596_/A vgnd vpwr scs8hd_diode_2
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_99 vgnd vpwr scs8hd_decap_4
XANTENNA__263__B _241_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_501 vgnd vpwr scs8hd_decap_12
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _301_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_SLEEPB _352_/Y vgnd vpwr scs8hd_diode_2
XFILLER_66_228 vgnd vpwr scs8hd_decap_6
XFILLER_47_431 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_144 vgnd vpwr scs8hd_decap_3
XFILLER_62_401 vgnd vpwr scs8hd_decap_8
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XANTENNA__438__B _471_/B vgnd vpwr scs8hd_diode_2
XFILLER_47_486 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _566_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__454__A _454_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_386 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__629__A _629_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_272 vpwr vgnd scs8hd_fill_2
XFILLER_25_103 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_SLEEPB _487_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_445 vpwr vgnd scs8hd_fill_2
XFILLER_25_158 vgnd vpwr scs8hd_decap_12
XFILLER_53_489 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_180 vgnd vpwr scs8hd_fill_1
XFILLER_40_128 vpwr vgnd scs8hd_fill_2
XANTENNA__364__A _391_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_515 vgnd vpwr scs8hd_fill_1
XFILLER_48_206 vgnd vpwr scs8hd_decap_8
X_641_ _641_/HI _641_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__539__A _591_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_283 vpwr vgnd scs8hd_fill_2
X_572_ _304_/B _562_/A _572_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_242 vpwr vgnd scs8hd_fill_2
XFILLER_71_220 vgnd vpwr scs8hd_decap_4
XFILLER_72_32 vgnd vpwr scs8hd_decap_12
XPHY_142 vgnd vpwr scs8hd_decap_3
XPHY_131 vgnd vpwr scs8hd_decap_3
XPHY_120 vgnd vpwr scs8hd_decap_3
XFILLER_24_180 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_decap_3
XPHY_153 vgnd vpwr scs8hd_decap_3
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__274__A _259_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_364 vgnd vpwr scs8hd_fill_1
XFILLER_8_324 vgnd vpwr scs8hd_decap_12
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_79_342 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA__449__A _385_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_401 vgnd vpwr scs8hd_decap_3
XFILLER_35_423 vpwr vgnd scs8hd_fill_2
XFILLER_62_231 vgnd vpwr scs8hd_decap_4
XFILLER_35_456 vgnd vpwr scs8hd_decap_3
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_489 vgnd vpwr scs8hd_decap_12
XFILLER_62_297 vpwr vgnd scs8hd_fill_2
XFILLER_22_128 vgnd vpwr scs8hd_decap_8
XFILLER_30_183 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_SLEEPB _454_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_504 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__359__A _358_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_220 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _248_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_53_275 vpwr vgnd scs8hd_fill_2
XFILLER_26_58 vgnd vpwr scs8hd_decap_6
XFILLER_41_404 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _597_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q
+ _518_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__541__B _542_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_312 vgnd vpwr scs8hd_decap_6
XFILLER_67_98 vgnd vpwr scs8hd_decap_4
XANTENNA__269__A _268_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q
+ _475_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_624_ _624_/A _624_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_445 vpwr vgnd scs8hd_fill_2
XFILLER_17_423 vpwr vgnd scs8hd_fill_2
XFILLER_29_283 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_489 vgnd vpwr scs8hd_decap_12
X_555_ _562_/A _561_/B vgnd vpwr scs8hd_buf_1
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
X_486_ _413_/A _490_/B _486_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_459 vgnd vpwr scs8hd_fill_1
XFILLER_12_161 vgnd vpwr scs8hd_decap_8
XFILLER_12_183 vgnd vpwr scs8hd_decap_8
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q
+ _432_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_187 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_301 vpwr vgnd scs8hd_fill_2
XFILLER_67_367 vgnd vpwr scs8hd_decap_3
XFILLER_67_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q
+ _375_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_82_304 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_SLEEPB _416_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_212 vpwr vgnd scs8hd_fill_2
XFILLER_23_437 vpwr vgnd scs8hd_fill_2
XFILLER_23_448 vpwr vgnd scs8hd_fill_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_50_267 vgnd vpwr scs8hd_decap_6
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XANTENNA__361__B _360_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _586_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_24 vpwr vgnd scs8hd_fill_2
XFILLER_73_326 vpwr vgnd scs8hd_fill_2
XFILLER_73_304 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_389 vgnd vpwr scs8hd_decap_8
XFILLER_37_79 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_34 vpwr vgnd scs8hd_fill_2
X_340_ _423_/A _340_/X vgnd vpwr scs8hd_buf_1
XFILLER_14_459 vgnd vpwr scs8hd_decap_12
XFILLER_41_234 vgnd vpwr scs8hd_decap_4
X_271_ _242_/A _271_/B _271_/X vgnd vpwr scs8hd_or2_4
XANTENNA__552__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__271__B _271_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_330 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_356 vpwr vgnd scs8hd_fill_2
XFILLER_49_367 vgnd vpwr scs8hd_fill_1
XFILLER_64_337 vgnd vpwr scs8hd_decap_4
X_607_ _607_/A _607_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__446__B _445_/B vgnd vpwr scs8hd_diode_2
XFILLER_60_510 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_17_297 vpwr vgnd scs8hd_fill_2
X_538_ _590_/A _542_/B _538_/Y vgnd vpwr scs8hd_nor2_4
X_469_ _447_/A _462_/A _469_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_429 vpwr vgnd scs8hd_fill_2
XFILLER_32_267 vpwr vgnd scs8hd_fill_2
XFILLER_9_452 vgnd vpwr scs8hd_decap_12
XANTENNA__462__A _462_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q
+ _349_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_SLEEPB _374_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_55_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_507 vgnd vpwr scs8hd_decap_8
XFILLER_82_156 vgnd vpwr scs8hd_decap_12
XFILLER_70_329 vgnd vpwr scs8hd_decap_4
XPHY_708 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _571_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_719 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_234 vpwr vgnd scs8hd_fill_2
XFILLER_23_256 vgnd vpwr scs8hd_decap_3
XANTENNA__356__B _356_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_8
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XANTENNA__372__A _314_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_SLEEPB _508_/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XANTENNA__547__A _599_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__266__B _587_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_323_ _314_/X _322_/X _323_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
X_254_ _286_/A _274_/B _330_/A vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__282__A _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
XFILLER_10_495 vgnd vpwr scs8hd_decap_12
XFILLER_6_422 vgnd vpwr scs8hd_decap_12
XFILLER_77_440 vgnd vpwr scs8hd_decap_12
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_37_315 vpwr vgnd scs8hd_fill_2
XFILLER_49_175 vpwr vgnd scs8hd_fill_2
XANTENNA__457__A _457_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_64_189 vgnd vpwr scs8hd_decap_4
XFILLER_60_351 vgnd vpwr scs8hd_decap_3
XFILLER_60_395 vpwr vgnd scs8hd_fill_2
XFILLER_60_384 vgnd vpwr scs8hd_decap_8
XFILLER_20_215 vgnd vpwr scs8hd_fill_1
XFILLER_20_237 vgnd vpwr scs8hd_decap_3
XFILLER_9_293 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_68_462 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_28_326 vgnd vpwr scs8hd_decap_3
XFILLER_28_337 vpwr vgnd scs8hd_fill_2
XFILLER_55_167 vpwr vgnd scs8hd_fill_2
XFILLER_55_156 vpwr vgnd scs8hd_fill_2
XANTENNA__367__A _340_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_359 vgnd vpwr scs8hd_decap_8
XFILLER_36_370 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_362 vpwr vgnd scs8hd_fill_2
XFILLER_34_69 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_403 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_SLEEPB _475_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_462 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_75_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__277__A _277_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_148 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_42_340 vgnd vpwr scs8hd_decap_4
XANTENNA__427__D _471_/D vgnd vpwr scs8hd_diode_2
X_306_ _305_/X _575_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_270 vgnd vpwr scs8hd_fill_1
X_237_ address[2] _286_/A vgnd vpwr scs8hd_inv_8
XFILLER_10_292 vgnd vpwr scs8hd_decap_12
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_226 vpwr vgnd scs8hd_fill_2
XFILLER_69_248 vpwr vgnd scs8hd_fill_2
XFILLER_69_237 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _545_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_281 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_80_446 vgnd vpwr scs8hd_decap_12
XFILLER_52_126 vgnd vpwr scs8hd_decap_6
XFILLER_21_513 vgnd vpwr scs8hd_decap_3
XFILLER_33_340 vgnd vpwr scs8hd_decap_4
XFILLER_60_181 vgnd vpwr scs8hd_decap_3
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_428 vgnd vpwr scs8hd_decap_6
XFILLER_29_47 vgnd vpwr scs8hd_decap_3
XFILLER_56_454 vpwr vgnd scs8hd_fill_2
XFILLER_28_134 vgnd vpwr scs8hd_fill_1
XFILLER_16_307 vpwr vgnd scs8hd_fill_2
XFILLER_43_104 vpwr vgnd scs8hd_fill_2
XFILLER_43_137 vgnd vpwr scs8hd_decap_4
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_351 vgnd vpwr scs8hd_decap_8
XFILLER_24_362 vgnd vpwr scs8hd_decap_4
XFILLER_61_34 vpwr vgnd scs8hd_fill_2
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_373 vgnd vpwr scs8hd_decap_8
XFILLER_24_384 vpwr vgnd scs8hd_fill_2
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__544__B _528_/X vgnd vpwr scs8hd_diode_2
XANTENNA__263__C _282_/C vgnd vpwr scs8hd_diode_2
XANTENNA__560__A _586_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_513 vgnd vpwr scs8hd_decap_3
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_421 vgnd vpwr scs8hd_decap_3
XANTENNA__438__C _409_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_104 vgnd vpwr scs8hd_decap_8
XFILLER_62_457 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_148 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_362 vpwr vgnd scs8hd_fill_2
XFILLER_15_351 vpwr vgnd scs8hd_fill_2
XFILLER_42_170 vgnd vpwr scs8hd_decap_8
XFILLER_42_181 vgnd vpwr scs8hd_decap_3
XANTENNA__454__B _456_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__470__A _448_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ _511_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_229 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ _468_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_65_262 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_295 vgnd vpwr scs8hd_decap_8
XFILLER_53_435 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_80_276 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__364__B _360_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_343 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ _424_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__380__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_23 vpwr vgnd scs8hd_fill_2
XFILLER_48_229 vgnd vpwr scs8hd_decap_3
X_640_ _640_/HI _640_/LO vgnd vpwr scs8hd_conb_1
XFILLER_56_45 vpwr vgnd scs8hd_fill_2
XANTENNA__539__B _542_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_443 vgnd vpwr scs8hd_fill_1
XFILLER_56_251 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ _368_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_465 vgnd vpwr scs8hd_decap_12
X_571_ _597_/A _562_/A _571_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_413 vpwr vgnd scs8hd_fill_2
XFILLER_71_232 vpwr vgnd scs8hd_fill_2
XFILLER_16_137 vpwr vgnd scs8hd_fill_2
XFILLER_72_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__555__A _562_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_44_468 vgnd vpwr scs8hd_decap_12
XPHY_143 vgnd vpwr scs8hd_decap_3
XPHY_132 vgnd vpwr scs8hd_decap_3
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_165 vgnd vpwr scs8hd_decap_3
XPHY_154 vgnd vpwr scs8hd_decap_3
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__274__B _274_/B vgnd vpwr scs8hd_diode_2
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__290__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_92 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_354 vgnd vpwr scs8hd_decap_12
XANTENNA__449__B _471_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q
+ _486_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_284 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__465__A _454_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_118 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _561_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_192 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q
+ _443_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_391 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_0_0_clk/X ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _616_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_424 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q
+ _391_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_265 vgnd vpwr scs8hd_decap_4
XFILLER_53_243 vgnd vpwr scs8hd_fill_1
XFILLER_26_468 vgnd vpwr scs8hd_decap_8
XFILLER_26_479 vgnd vpwr scs8hd_decap_12
XANTENNA__375__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_162 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_306 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ _335_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_623_ _623_/A _623_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XFILLER_17_479 vgnd vpwr scs8hd_decap_8
XFILLER_17_468 vpwr vgnd scs8hd_fill_2
X_554_ _553_/X _562_/A vgnd vpwr scs8hd_buf_1
XANTENNA__285__A _277_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_438 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_276 vgnd vpwr scs8hd_decap_4
X_485_ _407_/A _490_/B _485_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_449 vgnd vpwr scs8hd_decap_8
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XFILLER_8_144 vgnd vpwr scs8hd_decap_8
XFILLER_8_133 vpwr vgnd scs8hd_fill_2
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_4_361 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_184 vgnd vpwr scs8hd_decap_12
XFILLER_67_324 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _576_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_379 vpwr vgnd scs8hd_fill_2
XFILLER_35_221 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_405 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_35_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_460 vpwr vgnd scs8hd_fill_2
XFILLER_73_349 vpwr vgnd scs8hd_fill_2
XFILLER_73_338 vpwr vgnd scs8hd_fill_2
XFILLER_37_69 vgnd vpwr scs8hd_decap_4
XFILLER_26_254 vgnd vpwr scs8hd_fill_1
XFILLER_41_213 vpwr vgnd scs8hd_fill_2
XFILLER_53_79 vpwr vgnd scs8hd_fill_2
XFILLER_53_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_270_ _259_/A _270_/B _271_/B vgnd vpwr scs8hd_or2_4
XANTENNA__552__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_342 vgnd vpwr scs8hd_decap_12
XFILLER_49_302 vgnd vpwr scs8hd_decap_3
XFILLER_49_313 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_346 vgnd vpwr scs8hd_decap_6
XFILLER_76_154 vgnd vpwr scs8hd_decap_12
XFILLER_64_305 vgnd vpwr scs8hd_fill_1
XFILLER_57_390 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y _608_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
X_606_ _606_/A _606_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_537_ _589_/A _542_/B _537_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_224 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_SLEEPB _503_/Y vgnd vpwr scs8hd_diode_2
X_468_ _457_/A _467_/B _468_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
X_399_ _314_/X _404_/B _399_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_464 vgnd vpwr scs8hd_decap_12
XFILLER_40_290 vpwr vgnd scs8hd_fill_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_55_327 vpwr vgnd scs8hd_fill_2
XFILLER_82_168 vgnd vpwr scs8hd_decap_12
XPHY_709 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_63_382 vpwr vgnd scs8hd_fill_2
XANTENNA__372__B _376_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_290 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_132 vgnd vpwr scs8hd_fill_1
XFILLER_58_110 vgnd vpwr scs8hd_fill_1
XFILLER_58_154 vgnd vpwr scs8hd_decap_3
XFILLER_73_135 vgnd vpwr scs8hd_decap_12
XFILLER_58_187 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__547__B _526_/X vgnd vpwr scs8hd_diode_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
XFILLER_54_371 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_89 vgnd vpwr scs8hd_decap_3
X_322_ _344_/B _322_/X vgnd vpwr scs8hd_buf_1
XFILLER_80_44 vgnd vpwr scs8hd_decap_12
XANTENNA__563__A _589_/A vgnd vpwr scs8hd_diode_2
X_253_ _253_/A _274_/B vgnd vpwr scs8hd_buf_1
XANTENNA__282__B _241_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_434 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_SLEEPB _470_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_110 vpwr vgnd scs8hd_fill_2
XFILLER_49_132 vgnd vpwr scs8hd_decap_4
XFILLER_77_452 vgnd vpwr scs8hd_decap_12
XFILLER_64_102 vgnd vpwr scs8hd_decap_3
XANTENNA__457__B _456_/B vgnd vpwr scs8hd_diode_2
XFILLER_64_168 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_190 vgnd vpwr scs8hd_decap_12
XFILLER_60_363 vgnd vpwr scs8hd_decap_8
XANTENNA__473__A _481_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_249 vpwr vgnd scs8hd_fill_2
XFILLER_68_474 vgnd vpwr scs8hd_decap_12
XFILLER_28_305 vgnd vpwr scs8hd_fill_1
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA__367__B _367_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_105 vgnd vpwr scs8hd_decap_12
XFILLER_55_179 vpwr vgnd scs8hd_fill_2
XFILLER_43_319 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _544_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
XANTENNA__383__A address[8] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_47 vgnd vpwr scs8hd_decap_4
XFILLER_50_25 vgnd vpwr scs8hd_decap_4
XFILLER_3_415 vgnd vpwr scs8hd_decap_12
XFILLER_78_227 vgnd vpwr scs8hd_decap_12
XFILLER_59_56 vpwr vgnd scs8hd_fill_2
XFILLER_59_474 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_327 vgnd vpwr scs8hd_decap_3
XANTENNA__558__A _584_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_102 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _626_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__277__B _590_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_371 vpwr vgnd scs8hd_fill_2
XFILLER_61_127 vpwr vgnd scs8hd_fill_2
XFILLER_27_393 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
X_305_ _282_/C _241_/B _305_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_SLEEPB _437_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__293__A _278_/X vgnd vpwr scs8hd_diode_2
X_236_ _249_/A _242_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_69_216 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__468__A _457_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_293 vgnd vpwr scs8hd_decap_12
XFILLER_65_466 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_319 vpwr vgnd scs8hd_fill_2
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XFILLER_18_382 vgnd vpwr scs8hd_decap_4
XFILLER_18_393 vgnd vpwr scs8hd_decap_4
XFILLER_33_396 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_208 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _311_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__378__A _340_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XFILLER_56_466 vpwr vgnd scs8hd_fill_2
XFILLER_56_444 vgnd vpwr scs8hd_fill_1
XFILLER_28_124 vpwr vgnd scs8hd_fill_2
XFILLER_71_414 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_71_458 vgnd vpwr scs8hd_decap_12
XFILLER_45_58 vgnd vpwr scs8hd_fill_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_190 vpwr vgnd scs8hd_fill_2
XFILLER_51_171 vgnd vpwr scs8hd_fill_1
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_507 vgnd vpwr scs8hd_decap_8
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_79 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__560__B _561_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_260 vgnd vpwr scs8hd_decap_6
XANTENNA__288__A _288_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_455 vpwr vgnd scs8hd_fill_2
XFILLER_74_252 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XANTENNA__438__D _409_/D vgnd vpwr scs8hd_diode_2
XFILLER_47_466 vgnd vpwr scs8hd_decap_12
XFILLER_74_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_138 vgnd vpwr scs8hd_decap_4
XFILLER_15_330 vpwr vgnd scs8hd_fill_2
XFILLER_15_396 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_322 vgnd vpwr scs8hd_decap_3
XFILLER_35_91 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__470__B _462_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_65_241 vgnd vpwr scs8hd_fill_1
XFILLER_38_444 vgnd vpwr scs8hd_decap_12
XFILLER_53_425 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_SLEEPB _524_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_469 vgnd vpwr scs8hd_decap_12
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_80_288 vgnd vpwr scs8hd_decap_12
XFILLER_61_480 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_160 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_3
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_399 vpwr vgnd scs8hd_fill_2
XFILLER_31_27 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_400 vgnd vpwr scs8hd_decap_4
XFILLER_56_68 vgnd vpwr scs8hd_fill_1
XFILLER_29_477 vgnd vpwr scs8hd_decap_8
X_570_ _596_/A _562_/A _570_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_127 vgnd vpwr scs8hd_fill_1
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_72_56 vgnd vpwr scs8hd_decap_12
XFILLER_71_277 vpwr vgnd scs8hd_fill_2
XPHY_133 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_155 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_decap_3
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_388 vgnd vpwr scs8hd_decap_8
XFILLER_8_337 vgnd vpwr scs8hd_decap_12
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__571__A _597_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XANTENNA__290__B _330_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _591_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_208 vpwr vgnd scs8hd_fill_2
XFILLER_82_509 vgnd vpwr scs8hd_decap_6
XANTENNA__449__C _409_/C vgnd vpwr scs8hd_diode_2
XFILLER_47_241 vgnd vpwr scs8hd_decap_3
XFILLER_47_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_406 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__465__B _467_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
Xclkbuf_0_clk clk clkbuf_0_clk/X vgnd vpwr scs8hd_clkbuf_16
XANTENNA__481__A _448_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_285 vgnd vpwr scs8hd_decap_6
XFILLER_53_288 vpwr vgnd scs8hd_fill_2
XANTENNA__375__B _376_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_428 vgnd vpwr scs8hd_decap_3
XFILLER_21_130 vpwr vgnd scs8hd_fill_2
XFILLER_34_491 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__391__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_318 vgnd vpwr scs8hd_decap_12
XFILLER_1_513 vgnd vpwr scs8hd_decap_3
XFILLER_76_358 vgnd vpwr scs8hd_decap_12
X_622_ _622_/A _622_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_403 vgnd vpwr scs8hd_decap_4
XANTENNA__566__A _592_/A vgnd vpwr scs8hd_diode_2
X_553_ address[4] _552_/X _553_/X vgnd vpwr scs8hd_or2_4
XANTENNA__285__B _592_/A vgnd vpwr scs8hd_diode_2
X_484_ _491_/B _490_/B vgnd vpwr scs8hd_buf_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_373 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_79_196 vgnd vpwr scs8hd_decap_12
XFILLER_67_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _617_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _617_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__476__A _454_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_211 vgnd vpwr scs8hd_decap_4
XFILLER_50_203 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_225 vgnd vpwr scs8hd_decap_8
XFILLER_16_480 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_325 vgnd vpwr scs8hd_decap_8
XFILLER_73_306 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_233 vgnd vpwr scs8hd_fill_1
XANTENNA__386__A _385_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_417 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_266 vgnd vpwr scs8hd_decap_3
XFILLER_14_439 vgnd vpwr scs8hd_decap_4
XFILLER_41_258 vpwr vgnd scs8hd_fill_2
XFILLER_41_269 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_SLEEPB _326_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__552__C _578_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_78_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_354 vgnd vpwr scs8hd_decap_12
XFILLER_76_166 vgnd vpwr scs8hd_decap_12
XFILLER_64_317 vgnd vpwr scs8hd_decap_8
XFILLER_64_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
X_605_ _605_/A _605_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__296__A _282_/C vgnd vpwr scs8hd_diode_2
X_536_ _528_/X _542_/B vgnd vpwr scs8hd_buf_1
X_467_ _456_/A _467_/B _467_/Y vgnd vpwr scs8hd_nor2_4
X_398_ _405_/B _404_/B vgnd vpwr scs8hd_buf_1
XFILLER_9_476 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _281_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_306 vgnd vpwr scs8hd_decap_4
XFILLER_82_125 vgnd vpwr scs8hd_decap_12
XFILLER_48_391 vgnd vpwr scs8hd_decap_6
XFILLER_51_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_23_225 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_28 vpwr vgnd scs8hd_fill_2
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _635_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_122 vgnd vpwr scs8hd_decap_4
XFILLER_58_166 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_380 vpwr vgnd scs8hd_fill_2
XFILLER_73_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_54_383 vgnd vpwr scs8hd_decap_8
X_321_ _320_/X _344_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__563__B _568_/B vgnd vpwr scs8hd_diode_2
X_252_ _282_/C address[1] _253_/A vgnd vpwr scs8hd_or2_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__282__C _282_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_446 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_9 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_77_464 vgnd vpwr scs8hd_decap_12
XFILLER_37_328 vpwr vgnd scs8hd_fill_2
XFILLER_49_199 vgnd vpwr scs8hd_decap_3
XFILLER_64_158 vgnd vpwr scs8hd_fill_1
XFILLER_64_136 vpwr vgnd scs8hd_fill_2
XFILLER_33_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_SLEEPB _441_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_383 vpwr vgnd scs8hd_fill_2
X_519_ _413_/A _523_/B _519_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_206 vpwr vgnd scs8hd_fill_2
XFILLER_13_291 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_486 vgnd vpwr scs8hd_decap_12
XFILLER_55_114 vpwr vgnd scs8hd_fill_2
XFILLER_55_136 vgnd vpwr scs8hd_decap_3
XFILLER_70_117 vgnd vpwr scs8hd_decap_12
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _304_/Y vgnd vpwr scs8hd_diode_2
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__383__B _383_/B vgnd vpwr scs8hd_diode_2
XFILLER_50_15 vgnd vpwr scs8hd_decap_8
XFILLER_78_239 vgnd vpwr scs8hd_decap_12
XFILLER_59_431 vpwr vgnd scs8hd_fill_2
XFILLER_59_486 vpwr vgnd scs8hd_fill_2
XFILLER_19_306 vgnd vpwr scs8hd_decap_3
XFILLER_19_339 vpwr vgnd scs8hd_fill_2
XANTENNA__558__B _561_/B vgnd vpwr scs8hd_diode_2
XFILLER_74_456 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _591_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_501 vgnd vpwr scs8hd_decap_12
XFILLER_42_320 vpwr vgnd scs8hd_fill_2
XANTENNA__574__A _573_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_504 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__293__B _260_/B vgnd vpwr scs8hd_diode_2
X_304_ _301_/A _304_/B _304_/Y vgnd vpwr scs8hd_nor2_4
X_235_ address[3] _249_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_SLEEPB _399_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_7 vgnd vpwr scs8hd_fill_1
XFILLER_2_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_423 vgnd vpwr scs8hd_decap_4
XANTENNA__468__B _467_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_114 vpwr vgnd scs8hd_fill_2
XFILLER_65_434 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_489 vgnd vpwr scs8hd_decap_12
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_169 vgnd vpwr scs8hd_fill_1
XFILLER_80_459 vgnd vpwr scs8hd_decap_12
XANTENNA__484__A _491_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_38 vgnd vpwr scs8hd_decap_3
XFILLER_56_401 vgnd vpwr scs8hd_decap_8
XANTENNA__378__B _378_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_114 vgnd vpwr scs8hd_fill_1
XFILLER_45_15 vgnd vpwr scs8hd_decap_8
XFILLER_45_26 vpwr vgnd scs8hd_fill_2
XFILLER_71_437 vgnd vpwr scs8hd_decap_4
XFILLER_43_128 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__394__A _340_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_515 vgnd vpwr scs8hd_fill_1
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_58 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__569__A _294_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_47_412 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_74_242 vgnd vpwr scs8hd_fill_1
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
XFILLER_47_478 vgnd vpwr scs8hd_decap_8
XFILLER_47_489 vgnd vpwr scs8hd_decap_12
XFILLER_27_191 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_SLEEPB _361_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_194 vgnd vpwr scs8hd_decap_3
XFILLER_30_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__479__A _457_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_412 vgnd vpwr scs8hd_decap_4
XFILLER_65_231 vgnd vpwr scs8hd_decap_4
XFILLER_25_139 vpwr vgnd scs8hd_fill_2
XFILLER_18_180 vgnd vpwr scs8hd_fill_1
XFILLER_21_301 vpwr vgnd scs8hd_fill_2
XFILLER_21_323 vpwr vgnd scs8hd_fill_2
XFILLER_21_356 vgnd vpwr scs8hd_decap_4
XFILLER_21_378 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _565_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_507 vgnd vpwr scs8hd_decap_8
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XANTENNA__389__A _325_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_29_423 vpwr vgnd scs8hd_fill_2
XFILLER_29_456 vgnd vpwr scs8hd_decap_3
XFILLER_29_489 vgnd vpwr scs8hd_decap_12
XFILLER_16_106 vgnd vpwr scs8hd_decap_4
XFILLER_44_426 vgnd vpwr scs8hd_decap_12
XFILLER_72_68 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_decap_3
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XFILLER_31_109 vgnd vpwr scs8hd_decap_3
XPHY_156 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_decap_3
XFILLER_12_345 vpwr vgnd scs8hd_fill_2
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_194 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_378 vpwr vgnd scs8hd_fill_2
XFILLER_12_356 vgnd vpwr scs8hd_decap_8
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_349 vgnd vpwr scs8hd_decap_12
XANTENNA__571__B _562_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_367 vgnd vpwr scs8hd_decap_12
XANTENNA__299__A _286_/B vgnd vpwr scs8hd_diode_2
XANTENNA__449__D _471_/D vgnd vpwr scs8hd_diode_2
XFILLER_47_253 vpwr vgnd scs8hd_fill_2
XFILLER_62_201 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_47_297 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_62_289 vgnd vpwr scs8hd_decap_8
XFILLER_62_90 vpwr vgnd scs8hd_fill_2
XPHY_690 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__481__B _481_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_245 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA__391__B _387_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_337 vgnd vpwr scs8hd_decap_4
XFILLER_76_326 vpwr vgnd scs8hd_fill_2
X_621_ _621_/A _621_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_29_297 vpwr vgnd scs8hd_fill_2
XFILLER_44_223 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_552_ _380_/A address[7] _578_/C _515_/D _552_/X vgnd vpwr scs8hd_or4_4
XANTENNA__566__B _568_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_407 vgnd vpwr scs8hd_decap_8
X_483_ _482_/X _491_/B vgnd vpwr scs8hd_buf_1
XANTENNA__582__A _582_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_385 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_75_370 vpwr vgnd scs8hd_fill_2
XANTENNA__476__B _476_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_50_215 vgnd vpwr scs8hd_fill_1
XFILLER_23_418 vgnd vpwr scs8hd_decap_3
XFILLER_50_248 vpwr vgnd scs8hd_fill_2
XFILLER_16_492 vgnd vpwr scs8hd_decap_12
XANTENNA__492__A _425_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _539_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_348 vgnd vpwr scs8hd_decap_3
XFILLER_26_201 vpwr vgnd scs8hd_fill_2
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_407 vgnd vpwr scs8hd_decap_3
XFILLER_41_226 vpwr vgnd scs8hd_fill_2
XFILLER_22_462 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__552__D _515_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _560_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _639_/HI ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__577__A _274_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_178 vgnd vpwr scs8hd_decap_12
XFILLER_57_370 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_3
X_604_ _604_/A _604_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__296__B _241_/B vgnd vpwr scs8hd_diode_2
XFILLER_72_362 vgnd vpwr scs8hd_decap_4
XFILLER_17_278 vgnd vpwr scs8hd_decap_4
X_535_ _587_/A _529_/X _535_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_82 vgnd vpwr scs8hd_fill_1
XFILLER_32_204 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_466_ _466_/A _467_/B _466_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_451 vgnd vpwr scs8hd_decap_12
X_397_ _396_/X _405_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_134 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__487__A _509_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_137 vgnd vpwr scs8hd_decap_12
XFILLER_51_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_215 vgnd vpwr scs8hd_decap_8
XFILLER_23_248 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_15 vpwr vgnd scs8hd_fill_2
XANTENNA__397__A _396_/X vgnd vpwr scs8hd_diode_2
XFILLER_46_318 vgnd vpwr scs8hd_decap_4
XFILLER_73_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q
+ _412_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_226 vgnd vpwr scs8hd_decap_12
X_320_ address[8] _383_/B _320_/C _409_/D _320_/X vgnd vpwr scs8hd_or4_4
X_251_ _257_/A _584_/A _251_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_410 vgnd vpwr scs8hd_decap_12
XFILLER_80_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q
+ _362_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XFILLER_49_156 vpwr vgnd scs8hd_fill_2
XFILLER_77_476 vgnd vpwr scs8hd_decap_12
XFILLER_33_513 vgnd vpwr scs8hd_decap_3
XFILLER_45_362 vpwr vgnd scs8hd_fill_2
XFILLER_54_80 vgnd vpwr scs8hd_fill_1
X_518_ _407_/A _523_/B _518_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_398 vgnd vpwr scs8hd_decap_3
X_449_ _385_/A _471_/B _409_/C _471_/D _450_/A vgnd vpwr scs8hd_or4_4
XFILLER_9_241 vgnd vpwr scs8hd_decap_3
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_432 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_498 vgnd vpwr scs8hd_decap_12
XFILLER_55_104 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_318 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_SLEEPB _394_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_373 vgnd vpwr scs8hd_decap_4
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_343 vpwr vgnd scs8hd_fill_2
XFILLER_51_332 vgnd vpwr scs8hd_decap_4
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_207 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_428 vgnd vpwr scs8hd_decap_12
XFILLER_59_47 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_69 vgnd vpwr scs8hd_decap_4
XFILLER_59_443 vgnd vpwr scs8hd_decap_4
XFILLER_74_424 vgnd vpwr scs8hd_decap_12
XFILLER_19_318 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XFILLER_82_490 vgnd vpwr scs8hd_decap_6
XFILLER_61_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_303_ _302_/X _304_/B vgnd vpwr scs8hd_buf_1
XFILLER_42_376 vgnd vpwr scs8hd_decap_4
XFILLER_42_387 vpwr vgnd scs8hd_fill_2
XFILLER_42_398 vpwr vgnd scs8hd_fill_2
X_234_ _301_/A _257_/A vgnd vpwr scs8hd_buf_1
XANTENNA__590__A _590_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_273 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_288 vgnd vpwr scs8hd_decap_12
XFILLER_40_93 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_483 vgnd vpwr scs8hd_decap_12
XFILLER_37_148 vgnd vpwr scs8hd_decap_4
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XFILLER_37_159 vpwr vgnd scs8hd_fill_2
XFILLER_52_118 vpwr vgnd scs8hd_fill_2
XFILLER_18_373 vgnd vpwr scs8hd_decap_6
XFILLER_33_332 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_33_387 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_SLEEPB _355_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_240 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _569_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_148 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_118 vpwr vgnd scs8hd_fill_2
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__394__B _387_/A vgnd vpwr scs8hd_diode_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_184 vgnd vpwr scs8hd_decap_3
XFILLER_24_398 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_SLEEPB _490_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__569__B _562_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_273 vpwr vgnd scs8hd_fill_2
XFILLER_19_72 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_435 vgnd vpwr scs8hd_decap_4
XFILLER_74_265 vpwr vgnd scs8hd_fill_2
XFILLER_62_449 vgnd vpwr scs8hd_decap_6
XFILLER_62_438 vgnd vpwr scs8hd_decap_8
XANTENNA__585__A _585_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_376 vgnd vpwr scs8hd_decap_4
XFILLER_35_71 vgnd vpwr scs8hd_decap_3
XFILLER_30_346 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_81 vpwr vgnd scs8hd_fill_2
XANTENNA__479__B _476_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_468 vgnd vpwr scs8hd_decap_8
XFILLER_38_479 vgnd vpwr scs8hd_decap_12
XFILLER_80_202 vgnd vpwr scs8hd_decap_12
XFILLER_65_287 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_25_107 vpwr vgnd scs8hd_fill_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XANTENNA__495__A _495_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__389__B _387_/X vgnd vpwr scs8hd_diode_2
XFILLER_56_15 vgnd vpwr scs8hd_decap_8
XFILLER_29_446 vgnd vpwr scs8hd_fill_1
XFILLER_56_232 vgnd vpwr scs8hd_decap_8
XFILLER_71_224 vgnd vpwr scs8hd_fill_1
XFILLER_44_438 vgnd vpwr scs8hd_fill_1
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XFILLER_52_471 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_157 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_decap_3
XPHY_135 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_SLEEPB _457_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_335 vgnd vpwr scs8hd_fill_1
XFILLER_12_313 vgnd vpwr scs8hd_decap_12
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ _523_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__299__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_79_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_213 vgnd vpwr scs8hd_fill_1
XFILLER_62_246 vpwr vgnd scs8hd_fill_2
XFILLER_50_419 vgnd vpwr scs8hd_decap_6
XFILLER_15_140 vgnd vpwr scs8hd_decap_6
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_43_460 vpwr vgnd scs8hd_fill_2
XFILLER_43_471 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ _480_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_680 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_132 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_3
XPHY_691 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_187 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ _437_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_427 vpwr vgnd scs8hd_fill_2
XFILLER_38_276 vpwr vgnd scs8hd_fill_2
XFILLER_53_235 vpwr vgnd scs8hd_fill_2
XFILLER_53_224 vpwr vgnd scs8hd_fill_2
XFILLER_41_408 vpwr vgnd scs8hd_fill_2
XFILLER_41_419 vpwr vgnd scs8hd_fill_2
XFILLER_21_110 vgnd vpwr scs8hd_decap_8
XFILLER_21_121 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_39 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_SLEEPB _422_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_221 vpwr vgnd scs8hd_fill_2
X_620_ _620_/A _620_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_232 vpwr vgnd scs8hd_fill_2
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
X_551_ _274_/B _548_/X _551_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_449 vgnd vpwr scs8hd_decap_4
X_482_ _385_/A _382_/X _515_/C _482_/D _482_/X vgnd vpwr scs8hd_or4_4
XANTENNA__582__B _587_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q
+ _498_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _277_/Y vgnd vpwr scs8hd_diode_2
XFILLER_79_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q
+ _455_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_91 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ _403_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__492__B _491_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _530_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ _354_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_28 vpwr vgnd scs8hd_fill_2
XFILLER_81_330 vgnd vpwr scs8hd_decap_12
XFILLER_66_393 vgnd vpwr scs8hd_decap_4
XFILLER_26_224 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_SLEEPB _377_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_78_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_338 vpwr vgnd scs8hd_fill_2
XANTENNA__577__B _574_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_603_ _274_/B _600_/X _603_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_235 vpwr vgnd scs8hd_fill_2
XFILLER_17_224 vgnd vpwr scs8hd_decap_8
XFILLER_17_213 vpwr vgnd scs8hd_fill_2
XFILLER_27_72 vpwr vgnd scs8hd_fill_2
XANTENNA__296__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_72_341 vgnd vpwr scs8hd_fill_1
XFILLER_17_257 vpwr vgnd scs8hd_fill_2
X_534_ _586_/A _529_/X _534_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_396 vgnd vpwr scs8hd_fill_1
XFILLER_72_385 vgnd vpwr scs8hd_fill_1
X_465_ _454_/A _467_/B _465_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__593__A _593_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_463 vgnd vpwr scs8hd_decap_12
X_396_ _385_/A _382_/X _409_/C _471_/D _396_/X vgnd vpwr scs8hd_or4_4
XFILLER_43_71 vpwr vgnd scs8hd_fill_2
XFILLER_43_82 vpwr vgnd scs8hd_fill_2
XFILLER_9_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_SLEEPB _511_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_67_102 vgnd vpwr scs8hd_fill_1
XFILLER_67_157 vpwr vgnd scs8hd_fill_2
XFILLER_67_146 vpwr vgnd scs8hd_fill_2
XANTENNA__487__B _490_/B vgnd vpwr scs8hd_diode_2
XFILLER_67_168 vpwr vgnd scs8hd_fill_2
XFILLER_82_149 vgnd vpwr scs8hd_decap_6
XFILLER_63_352 vpwr vgnd scs8hd_fill_2
XFILLER_63_341 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_238 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_102 vgnd vpwr scs8hd_decap_8
XFILLER_48_38 vpwr vgnd scs8hd_fill_2
XFILLER_48_49 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_330 vgnd vpwr scs8hd_fill_1
XFILLER_39_393 vgnd vpwr scs8hd_decap_4
XFILLER_54_352 vpwr vgnd scs8hd_fill_2
XFILLER_54_341 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_171 vgnd vpwr scs8hd_decap_12
XFILLER_54_396 vgnd vpwr scs8hd_fill_1
XFILLER_14_249 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_250_ _249_/X _584_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_422 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_459 vgnd vpwr scs8hd_decap_12
XANTENNA__588__A _581_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_352 vpwr vgnd scs8hd_fill_2
XFILLER_60_322 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_517_ _517_/A _523_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_SLEEPB _478_/Y vgnd vpwr scs8hd_diode_2
X_448_ _448_/A _448_/B _448_/Y vgnd vpwr scs8hd_nor2_4
X_379_ _395_/A _378_/B _379_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_70_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y _630_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__498__A _509_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_308 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_503 vgnd vpwr scs8hd_decap_12
XFILLER_36_341 vgnd vpwr scs8hd_decap_3
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_377 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_8
XFILLER_59_422 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_74_436 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_54_160 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_182 vpwr vgnd scs8hd_fill_2
XFILLER_42_333 vgnd vpwr scs8hd_decap_3
X_302_ _278_/X _302_/B _302_/X vgnd vpwr scs8hd_or2_4
XFILLER_24_73 vgnd vpwr scs8hd_decap_3
X_233_ _233_/A _301_/A vgnd vpwr scs8hd_buf_1
XANTENNA__590__B _594_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_208 vgnd vpwr scs8hd_decap_8
XFILLER_2_495 vgnd vpwr scs8hd_decap_12
XFILLER_65_414 vgnd vpwr scs8hd_decap_3
XFILLER_65_403 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_344 vgnd vpwr scs8hd_fill_1
XFILLER_45_193 vpwr vgnd scs8hd_fill_2
XFILLER_60_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _618_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_274 vgnd vpwr scs8hd_fill_1
XFILLER_68_285 vpwr vgnd scs8hd_fill_2
XFILLER_56_436 vgnd vpwr scs8hd_decap_8
XFILLER_43_108 vgnd vpwr scs8hd_decap_3
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_366 vgnd vpwr scs8hd_fill_1
XFILLER_24_388 vpwr vgnd scs8hd_fill_2
XFILLER_61_49 vgnd vpwr scs8hd_decap_3
XFILLER_51_196 vpwr vgnd scs8hd_fill_2
XFILLER_51_174 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _549_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_241 vgnd vpwr scs8hd_fill_1
XFILLER_19_51 vgnd vpwr scs8hd_decap_4
XFILLER_19_62 vgnd vpwr scs8hd_fill_1
XANTENNA__585__B _587_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_303 vgnd vpwr scs8hd_decap_3
XPHY_840 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_314 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_65_266 vgnd vpwr scs8hd_decap_4
XFILLER_53_406 vpwr vgnd scs8hd_fill_2
XFILLER_53_417 vpwr vgnd scs8hd_fill_2
XFILLER_33_130 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _584_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ _491_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ _448_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_222 vgnd vpwr scs8hd_fill_1
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_56_49 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_16_119 vgnd vpwr scs8hd_decap_8
XFILLER_72_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_258 vpwr vgnd scs8hd_fill_2
XFILLER_71_236 vgnd vpwr scs8hd_decap_4
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XFILLER_52_450 vgnd vpwr scs8hd_decap_8
XPHY_103 vgnd vpwr scs8hd_decap_3
XFILLER_24_141 vpwr vgnd scs8hd_fill_2
XPHY_158 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_decap_3
XPHY_136 vgnd vpwr scs8hd_decap_3
XFILLER_52_483 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y _619_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__299__C address[3] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__596__A _596_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_233 vpwr vgnd scs8hd_fill_2
XFILLER_35_406 vpwr vgnd scs8hd_fill_2
XFILLER_47_266 vpwr vgnd scs8hd_fill_2
XFILLER_35_439 vpwr vgnd scs8hd_fill_2
XFILLER_15_130 vgnd vpwr scs8hd_fill_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_70_280 vgnd vpwr scs8hd_fill_1
XFILLER_15_196 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XPHY_670 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_692 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_681 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_166 vgnd vpwr scs8hd_decap_6
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_38_222 vgnd vpwr scs8hd_decap_4
XFILLER_81_501 vgnd vpwr scs8hd_decap_12
XFILLER_19_480 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_69_380 vpwr vgnd scs8hd_fill_2
XFILLER_67_59 vpwr vgnd scs8hd_fill_2
XFILLER_29_200 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_428 vpwr vgnd scs8hd_fill_2
X_550_ _270_/B _548_/X _550_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_203 vpwr vgnd scs8hd_fill_2
X_481_ _448_/A _481_/B _481_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_442 vgnd vpwr scs8hd_decap_4
XFILLER_4_398 vgnd vpwr scs8hd_decap_12
XFILLER_67_306 vgnd vpwr scs8hd_decap_3
XFILLER_75_350 vpwr vgnd scs8hd_fill_2
XFILLER_63_501 vgnd vpwr scs8hd_decap_12
XFILLER_35_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_206 vgnd vpwr scs8hd_decap_4
XFILLER_35_258 vpwr vgnd scs8hd_fill_2
XFILLER_31_464 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_192 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _632_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_317 vgnd vpwr scs8hd_fill_1
XFILLER_66_372 vgnd vpwr scs8hd_decap_6
XFILLER_26_236 vpwr vgnd scs8hd_fill_2
XFILLER_81_342 vgnd vpwr scs8hd_decap_12
XFILLER_26_247 vgnd vpwr scs8hd_decap_4
XFILLER_26_258 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_39 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XFILLER_49_317 vpwr vgnd scs8hd_fill_2
XFILLER_57_361 vgnd vpwr scs8hd_fill_1
X_602_ _270_/B _600_/X _602_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_501 vgnd vpwr scs8hd_decap_12
XFILLER_57_394 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_62 vgnd vpwr scs8hd_fill_1
XANTENNA__296__D _259_/A vgnd vpwr scs8hd_diode_2
X_533_ _585_/A _529_/X _533_/Y vgnd vpwr scs8hd_nor2_4
X_464_ _442_/A _467_/B _464_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__593__B _594_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_475 vgnd vpwr scs8hd_decap_12
X_395_ _395_/A _387_/A _395_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_272 vgnd vpwr scs8hd_decap_3
XFILLER_40_283 vgnd vpwr scs8hd_decap_4
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_80 vgnd vpwr scs8hd_decap_12
XFILLER_67_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_82_106 vgnd vpwr scs8hd_decap_12
XFILLER_63_386 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_283 vpwr vgnd scs8hd_fill_2
XFILLER_31_294 vpwr vgnd scs8hd_fill_2
XFILLER_58_136 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _575_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_501 vgnd vpwr scs8hd_decap_12
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_54_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_8
XFILLER_42_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_261 vpwr vgnd scs8hd_fill_2
XFILLER_10_434 vgnd vpwr scs8hd_decap_12
XFILLER_22_283 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_6
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_114 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_136 vgnd vpwr scs8hd_fill_1
XFILLER_77_489 vgnd vpwr scs8hd_decap_12
XFILLER_37_309 vgnd vpwr scs8hd_decap_4
XFILLER_57_180 vgnd vpwr scs8hd_decap_3
XFILLER_45_331 vpwr vgnd scs8hd_fill_2
X_516_ _516_/A _517_/A vgnd vpwr scs8hd_buf_1
XFILLER_60_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_447_ _447_/A _448_/B _447_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_210 vgnd vpwr scs8hd_decap_4
X_378_ _340_/X _378_/B _378_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XANTENNA__498__B _499_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_515 vgnd vpwr scs8hd_fill_1
XFILLER_36_364 vgnd vpwr scs8hd_decap_6
XFILLER_51_367 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_401 vpwr vgnd scs8hd_fill_2
XFILLER_75_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_489 vgnd vpwr scs8hd_decap_12
XFILLER_75_59 vpwr vgnd scs8hd_fill_2
XFILLER_74_448 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_459 vgnd vpwr scs8hd_decap_12
XFILLER_42_312 vgnd vpwr scs8hd_decap_8
XFILLER_27_397 vpwr vgnd scs8hd_fill_2
XFILLER_24_41 vpwr vgnd scs8hd_fill_2
X_301_ _301_/A _597_/A _301_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_85 vgnd vpwr scs8hd_decap_4
X_232_ address[4] _231_/X _233_/A vgnd vpwr scs8hd_or2_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_40_62 vpwr vgnd scs8hd_fill_2
XFILLER_40_73 vpwr vgnd scs8hd_fill_2
XFILLER_40_84 vgnd vpwr scs8hd_decap_3
XANTENNA__599__A _599_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_220 vgnd vpwr scs8hd_decap_12
XFILLER_49_71 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_301 vpwr vgnd scs8hd_fill_2
XFILLER_60_164 vgnd vpwr scs8hd_decap_8
XFILLER_33_356 vpwr vgnd scs8hd_fill_2
XFILLER_33_367 vpwr vgnd scs8hd_fill_2
XFILLER_60_186 vpwr vgnd scs8hd_fill_2
XFILLER_60_175 vgnd vpwr scs8hd_decap_4
XANTENNA__302__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_68_264 vpwr vgnd scs8hd_fill_2
XFILLER_68_253 vgnd vpwr scs8hd_decap_8
XFILLER_28_106 vgnd vpwr scs8hd_decap_8
XFILLER_28_128 vgnd vpwr scs8hd_decap_6
XFILLER_71_418 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_194 vgnd vpwr scs8hd_decap_4
XFILLER_51_153 vpwr vgnd scs8hd_fill_2
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_507 vgnd vpwr scs8hd_decap_8
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_220 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_404 vpwr vgnd scs8hd_fill_2
XFILLER_59_297 vpwr vgnd scs8hd_fill_2
XFILLER_59_286 vpwr vgnd scs8hd_fill_2
XFILLER_19_41 vgnd vpwr scs8hd_decap_4
XFILLER_19_106 vpwr vgnd scs8hd_fill_2
XFILLER_47_426 vgnd vpwr scs8hd_fill_1
XFILLER_74_256 vgnd vpwr scs8hd_decap_6
XFILLER_74_234 vgnd vpwr scs8hd_decap_8
XFILLER_74_289 vgnd vpwr scs8hd_decap_12
XFILLER_15_334 vpwr vgnd scs8hd_fill_2
XFILLER_42_131 vgnd vpwr scs8hd_decap_3
XPHY_841 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_830 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_95 vgnd vpwr scs8hd_decap_4
XFILLER_42_186 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_94 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_80 vgnd vpwr scs8hd_decap_12
XFILLER_65_245 vgnd vpwr scs8hd_decap_4
XFILLER_80_215 vgnd vpwr scs8hd_decap_12
XFILLER_61_451 vpwr vgnd scs8hd_fill_2
XFILLER_33_153 vgnd vpwr scs8hd_fill_1
XFILLER_21_315 vpwr vgnd scs8hd_fill_2
XFILLER_33_164 vpwr vgnd scs8hd_fill_2
XFILLER_33_197 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _594_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_267 vgnd vpwr scs8hd_decap_8
XFILLER_71_248 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_72_27 vgnd vpwr scs8hd_decap_4
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_decap_3
XPHY_137 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XFILLER_52_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_decap_3
XFILLER_12_337 vgnd vpwr scs8hd_decap_8
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XANTENNA__299__D _259_/A vgnd vpwr scs8hd_diode_2
XANTENNA__596__B _581_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_223 vgnd vpwr scs8hd_fill_1
XFILLER_47_245 vgnd vpwr scs8hd_fill_1
XFILLER_62_215 vgnd vpwr scs8hd_decap_3
XFILLER_46_61 vpwr vgnd scs8hd_fill_2
XFILLER_62_259 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XPHY_671 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_660 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_145 vgnd vpwr scs8hd_decap_8
XPHY_693 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_682 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_330 vgnd vpwr scs8hd_decap_12
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_510 vgnd vpwr scs8hd_decap_6
XFILLER_81_513 vgnd vpwr scs8hd_decap_3
XFILLER_26_407 vgnd vpwr scs8hd_decap_8
XFILLER_26_418 vgnd vpwr scs8hd_decap_6
XFILLER_21_145 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _601_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_17_407 vgnd vpwr scs8hd_fill_1
XFILLER_44_215 vpwr vgnd scs8hd_fill_2
X_480_ _447_/A _481_/B _480_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_101 vpwr vgnd scs8hd_fill_2
XFILLER_25_462 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_134 vgnd vpwr scs8hd_decap_4
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_8_138 vgnd vpwr scs8hd_decap_4
XFILLER_32_74 vpwr vgnd scs8hd_fill_2
XFILLER_4_300 vgnd vpwr scs8hd_decap_12
XFILLER_32_96 vpwr vgnd scs8hd_fill_2
XFILLER_79_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__400__A _325_/X vgnd vpwr scs8hd_diode_2
XFILLER_63_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_SLEEPB _335_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_443 vgnd vpwr scs8hd_decap_4
XFILLER_31_476 vgnd vpwr scs8hd_fill_1
XFILLER_31_487 vgnd vpwr scs8hd_fill_1
XFILLER_78_3 vgnd vpwr scs8hd_decap_12
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_182 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _298_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_58_307 vpwr vgnd scs8hd_fill_2
XANTENNA__310__A _575_/A vgnd vpwr scs8hd_diode_2
XFILLER_66_362 vpwr vgnd scs8hd_fill_2
XFILLER_66_351 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_354 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_410 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _624_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
X_601_ _575_/A _600_/X _601_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_513 vgnd vpwr scs8hd_decap_3
XFILLER_27_85 vpwr vgnd scs8hd_fill_2
X_532_ _584_/A _529_/X _532_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_398 vgnd vpwr scs8hd_decap_8
X_463_ _441_/A _467_/B _463_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_281 vpwr vgnd scs8hd_fill_2
XFILLER_43_40 vpwr vgnd scs8hd_fill_2
XFILLER_9_403 vgnd vpwr scs8hd_decap_12
X_394_ _340_/X _387_/A _394_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_43_51 vpwr vgnd scs8hd_fill_2
XFILLER_13_487 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _633_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XFILLER_67_126 vpwr vgnd scs8hd_fill_2
XFILLER_82_118 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_48_373 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__305__A _282_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_SLEEPB _444_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_340 vgnd vpwr scs8hd_decap_4
XFILLER_39_362 vpwr vgnd scs8hd_fill_2
XFILLER_27_513 vgnd vpwr scs8hd_decap_3
XFILLER_54_365 vgnd vpwr scs8hd_decap_6
XFILLER_81_184 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_22_273 vpwr vgnd scs8hd_fill_2
XFILLER_10_446 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_107 vgnd vpwr scs8hd_decap_3
XFILLER_38_62 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_73 vpwr vgnd scs8hd_fill_2
XFILLER_38_84 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _244_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _556_/Y vgnd vpwr scs8hd_diode_2
X_515_ _409_/A _382_/A _515_/C _515_/D _516_/A vgnd vpwr scs8hd_or4_4
XFILLER_60_346 vgnd vpwr scs8hd_decap_3
XFILLER_54_72 vpwr vgnd scs8hd_fill_2
XFILLER_45_398 vgnd vpwr scs8hd_decap_4
X_446_ _457_/A _445_/B _446_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
X_377_ _404_/A _376_/B _377_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _596_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_295 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_70_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q
+ _474_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_118 vpwr vgnd scs8hd_fill_2
XFILLER_51_313 vpwr vgnd scs8hd_fill_2
XFILLER_63_195 vpwr vgnd scs8hd_fill_2
XFILLER_63_184 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_SLEEPB _402_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q
+ _431_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_28 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_435 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q
+ _374_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_27 vgnd vpwr scs8hd_decap_12
XFILLER_74_405 vpwr vgnd scs8hd_fill_2
XFILLER_46_107 vgnd vpwr scs8hd_decap_12
XFILLER_46_129 vpwr vgnd scs8hd_fill_2
XFILLER_27_343 vpwr vgnd scs8hd_fill_2
XFILLER_54_151 vpwr vgnd scs8hd_fill_2
XFILLER_27_354 vpwr vgnd scs8hd_fill_2
XFILLER_27_376 vpwr vgnd scs8hd_fill_2
X_300_ _299_/X _597_/A vgnd vpwr scs8hd_buf_1
XFILLER_42_346 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_231_ address[6] _471_/B _515_/C _515_/D _231_/X vgnd vpwr scs8hd_or4_4
XFILLER_10_276 vpwr vgnd scs8hd_fill_2
XFILLER_40_41 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__599__B _578_/X vgnd vpwr scs8hd_diode_2
XFILLER_77_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_83 vgnd vpwr scs8hd_fill_1
XFILLER_65_438 vpwr vgnd scs8hd_fill_2
XFILLER_18_310 vpwr vgnd scs8hd_fill_2
XFILLER_37_118 vgnd vpwr scs8hd_decap_4
XFILLER_37_129 vpwr vgnd scs8hd_fill_2
XFILLER_18_332 vpwr vgnd scs8hd_fill_2
XFILLER_73_471 vgnd vpwr scs8hd_decap_12
XFILLER_60_154 vgnd vpwr scs8hd_fill_1
XFILLER_33_379 vpwr vgnd scs8hd_fill_2
X_429_ _429_/A _429_/X vgnd vpwr scs8hd_buf_1
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XANTENNA__302__B _302_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_SLEEPB _364_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _310_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_313 vgnd vpwr scs8hd_decap_12
XFILLER_51_132 vpwr vgnd scs8hd_fill_2
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_346 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y _607_/A vgnd vpwr scs8hd_inv_1
XFILLER_74_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_55_471 vpwr vgnd scs8hd_fill_2
XFILLER_15_302 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _570_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_313 vpwr vgnd scs8hd_fill_2
XFILLER_27_195 vpwr vgnd scs8hd_fill_2
XFILLER_35_30 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_SLEEPB _498_/Y vgnd vpwr scs8hd_diode_2
XPHY_820 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_463 vgnd vpwr scs8hd_decap_12
XFILLER_42_143 vpwr vgnd scs8hd_fill_2
XPHY_842 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_831 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_165 vpwr vgnd scs8hd_fill_2
XFILLER_51_62 vgnd vpwr scs8hd_decap_4
XFILLER_7_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__403__A _392_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_213 vpwr vgnd scs8hd_fill_2
XFILLER_38_427 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_227 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_327 vgnd vpwr scs8hd_decap_3
XFILLER_33_176 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__313__A _313_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_213 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_decap_3
XPHY_138 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XFILLER_12_327 vgnd vpwr scs8hd_decap_8
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XFILLER_12_349 vgnd vpwr scs8hd_decap_4
XFILLER_20_393 vgnd vpwr scs8hd_decap_4
XFILLER_4_515 vgnd vpwr scs8hd_fill_1
XFILLER_21_54 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_SLEEPB _465_/Y vgnd vpwr scs8hd_diode_2
XFILLER_62_205 vgnd vpwr scs8hd_decap_8
XFILLER_35_419 vpwr vgnd scs8hd_fill_2
XFILLER_46_51 vgnd vpwr scs8hd_fill_1
XFILLER_62_238 vgnd vpwr scs8hd_decap_8
XFILLER_62_227 vpwr vgnd scs8hd_fill_2
XFILLER_28_471 vgnd vpwr scs8hd_decap_12
XFILLER_46_73 vpwr vgnd scs8hd_fill_2
XFILLER_46_84 vgnd vpwr scs8hd_decap_8
XFILLER_55_290 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_187 vgnd vpwr scs8hd_decap_3
XFILLER_62_61 vgnd vpwr scs8hd_decap_4
XPHY_661 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_650 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_113 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y _625_/A vgnd vpwr scs8hd_inv_1
XPHY_694 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_683 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_672 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_342 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_246 vgnd vpwr scs8hd_decap_8
XFILLER_53_205 vpwr vgnd scs8hd_fill_2
XFILLER_53_216 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _539_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_249 vgnd vpwr scs8hd_fill_1
XFILLER_61_271 vpwr vgnd scs8hd_fill_2
XFILLER_61_260 vpwr vgnd scs8hd_fill_2
XANTENNA__308__A _599_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_179 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _544_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_279 vpwr vgnd scs8hd_fill_2
XFILLER_44_227 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_SLEEPB _432_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_157 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XFILLER_4_312 vgnd vpwr scs8hd_decap_12
XFILLER_79_135 vgnd vpwr scs8hd_decap_12
XANTENNA__400__B _404_/B vgnd vpwr scs8hd_diode_2
XFILLER_57_83 vgnd vpwr scs8hd_decap_3
XFILLER_75_374 vgnd vpwr scs8hd_decap_12
XFILLER_28_290 vpwr vgnd scs8hd_fill_2
XFILLER_43_271 vpwr vgnd scs8hd_fill_2
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_330 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__310__B _309_/X vgnd vpwr scs8hd_diode_2
XFILLER_78_190 vgnd vpwr scs8hd_decap_12
XFILLER_66_341 vgnd vpwr scs8hd_fill_1
XFILLER_26_205 vgnd vpwr scs8hd_decap_4
XFILLER_34_271 vpwr vgnd scs8hd_fill_2
XFILLER_22_466 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _531_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q
+ _510_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__501__A _523_/A vgnd vpwr scs8hd_diode_2
XFILLER_76_105 vgnd vpwr scs8hd_decap_12
XFILLER_57_330 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
X_600_ _599_/X _600_/X vgnd vpwr scs8hd_buf_1
XFILLER_72_311 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ _467_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_374 vgnd vpwr scs8hd_decap_4
X_531_ _583_/A _529_/X _531_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_42 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_72_388 vgnd vpwr scs8hd_decap_8
XFILLER_72_366 vgnd vpwr scs8hd_fill_1
X_462_ _462_/A _467_/B vgnd vpwr scs8hd_buf_1
XFILLER_13_400 vpwr vgnd scs8hd_fill_2
XFILLER_32_208 vgnd vpwr scs8hd_decap_6
XFILLER_25_293 vgnd vpwr scs8hd_fill_1
X_393_ _404_/A _387_/X _393_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_415 vgnd vpwr scs8hd_decap_12
XFILLER_40_252 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ _422_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__411__A _411_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_68_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ _367_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_48_341 vpwr vgnd scs8hd_fill_2
XFILLER_75_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_SLEEPB _519_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_399 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vpwr vgnd scs8hd_fill_2
XFILLER_31_241 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__305__B _241_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__321__A _320_/X vgnd vpwr scs8hd_diode_2
XFILLER_48_19 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_333 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q
+ _485_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_81_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_296 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q
+ _442_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_99 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_77_403 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__231__A address[6] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_41 vpwr vgnd scs8hd_fill_2
XFILLER_64_119 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q
+ _390_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_72_141 vgnd vpwr scs8hd_decap_12
XFILLER_60_303 vgnd vpwr scs8hd_decap_4
X_514_ _425_/A _505_/X _514_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_54_84 vgnd vpwr scs8hd_decap_6
XFILLER_54_62 vgnd vpwr scs8hd_fill_1
X_445_ _456_/A _445_/B _445_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_230 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_274 vpwr vgnd scs8hd_fill_2
X_376_ _392_/A _376_/B _376_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__406__A _395_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q
+ _332_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_440 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_108 vgnd vpwr scs8hd_decap_4
XFILLER_48_182 vgnd vpwr scs8hd_decap_4
XFILLER_36_377 vgnd vpwr scs8hd_fill_1
XFILLER_51_336 vgnd vpwr scs8hd_fill_1
XFILLER_51_358 vpwr vgnd scs8hd_fill_2
XANTENNA__316__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _575_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_458 vpwr vgnd scs8hd_fill_2
XFILLER_75_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_311 vpwr vgnd scs8hd_fill_2
XFILLER_46_119 vgnd vpwr scs8hd_fill_1
XFILLER_39_193 vpwr vgnd scs8hd_fill_2
XFILLER_54_196 vgnd vpwr scs8hd_fill_1
XFILLER_42_325 vpwr vgnd scs8hd_fill_2
X_230_ _230_/A address[5] _515_/D vgnd vpwr scs8hd_or2_4
XFILLER_10_222 vgnd vpwr scs8hd_decap_12
XANTENNA__226__A address[7] vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _572_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_410 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_95 vpwr vgnd scs8hd_fill_2
XFILLER_65_428 vgnd vpwr scs8hd_decap_3
XFILLER_58_480 vgnd vpwr scs8hd_decap_12
XFILLER_73_483 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_336 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_428_ _428_/A _429_/A vgnd vpwr scs8hd_buf_1
XFILLER_60_199 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_380 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_359_ _358_/X _367_/B vgnd vpwr scs8hd_buf_1
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_281 vgnd vpwr scs8hd_decap_12
XFILLER_64_450 vgnd vpwr scs8hd_decap_8
XFILLER_24_303 vgnd vpwr scs8hd_fill_1
XFILLER_36_163 vgnd vpwr scs8hd_decap_12
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_369 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_233 vpwr vgnd scs8hd_fill_2
XFILLER_47_417 vpwr vgnd scs8hd_fill_2
XFILLER_19_76 vpwr vgnd scs8hd_fill_2
XFILLER_47_439 vgnd vpwr scs8hd_fill_1
XFILLER_74_269 vgnd vpwr scs8hd_decap_6
XFILLER_62_409 vgnd vpwr scs8hd_decap_3
XFILLER_55_461 vgnd vpwr scs8hd_fill_1
XFILLER_82_280 vgnd vpwr scs8hd_decap_12
XFILLER_35_20 vgnd vpwr scs8hd_decap_4
XPHY_810 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_358 vpwr vgnd scs8hd_fill_2
XFILLER_15_347 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XPHY_843 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_832 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_821 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_475 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_328 vpwr vgnd scs8hd_fill_2
XFILLER_23_380 vgnd vpwr scs8hd_fill_1
XFILLER_7_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__403__B _404_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_76_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_450 vgnd vpwr scs8hd_decap_8
XFILLER_80_239 vgnd vpwr scs8hd_decap_12
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
XFILLER_33_111 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_464 vpwr vgnd scs8hd_fill_2
XFILLER_14_391 vpwr vgnd scs8hd_fill_2
XFILLER_21_339 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y _622_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_406 vpwr vgnd scs8hd_fill_2
XFILLER_29_439 vgnd vpwr scs8hd_decap_4
XFILLER_44_409 vpwr vgnd scs8hd_fill_2
XFILLER_71_228 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_431 vpwr vgnd scs8hd_fill_2
XPHY_106 vgnd vpwr scs8hd_decap_3
XFILLER_24_122 vpwr vgnd scs8hd_fill_2
XPHY_139 vgnd vpwr scs8hd_decap_3
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_350 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_33 vpwr vgnd scs8hd_fill_2
XANTENNA__504__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_88 vpwr vgnd scs8hd_fill_2
XFILLER_79_306 vgnd vpwr scs8hd_decap_12
XFILLER_75_501 vgnd vpwr scs8hd_decap_12
XFILLER_47_203 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_483 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_43_431 vpwr vgnd scs8hd_fill_2
XFILLER_43_453 vpwr vgnd scs8hd_fill_2
XFILLER_70_272 vgnd vpwr scs8hd_decap_3
XFILLER_70_261 vgnd vpwr scs8hd_fill_1
XFILLER_43_464 vpwr vgnd scs8hd_fill_2
XFILLER_43_475 vgnd vpwr scs8hd_decap_12
XFILLER_70_294 vgnd vpwr scs8hd_decap_8
XFILLER_70_283 vpwr vgnd scs8hd_fill_2
XFILLER_62_40 vgnd vpwr scs8hd_fill_1
XPHY_662 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_651 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_640 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_136 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_695 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_684 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_673 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__414__A _442_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ _503_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_361 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_239 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _289_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__308__B _231_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__324__A _324_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _535_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_501 vgnd vpwr scs8hd_decap_12
XFILLER_29_225 vpwr vgnd scs8hd_fill_2
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
XFILLER_72_515 vgnd vpwr scs8hd_fill_1
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_291 vgnd vpwr scs8hd_fill_1
XFILLER_25_475 vpwr vgnd scs8hd_fill_2
XFILLER_40_401 vpwr vgnd scs8hd_fill_2
XFILLER_40_456 vpwr vgnd scs8hd_fill_2
XFILLER_8_129 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_3
XFILLER_32_54 vgnd vpwr scs8hd_decap_3
XFILLER_20_191 vgnd vpwr scs8hd_decap_4
XFILLER_32_87 vpwr vgnd scs8hd_fill_2
XANTENNA__234__A _301_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_324 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _310_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_95 vpwr vgnd scs8hd_fill_2
XFILLER_57_73 vpwr vgnd scs8hd_fill_2
XFILLER_75_386 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_217 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__409__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_453 vpwr vgnd scs8hd_fill_2
XFILLER_31_401 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_423 vpwr vgnd scs8hd_fill_2
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_489 vgnd vpwr scs8hd_decap_12
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_191 vgnd vpwr scs8hd_decap_3
XFILLER_7_184 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _619_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_501 vgnd vpwr scs8hd_decap_12
XFILLER_54_504 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__319__A _482_/D vgnd vpwr scs8hd_diode_2
XFILLER_81_367 vgnd vpwr scs8hd_decap_12
XFILLER_41_209 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_SLEEPB _514_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_434 vgnd vpwr scs8hd_decap_3
XFILLER_22_456 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_478 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__501__B _499_/B vgnd vpwr scs8hd_diode_2
XFILLER_49_309 vpwr vgnd scs8hd_fill_2
XFILLER_76_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_353 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_364 vpwr vgnd scs8hd_fill_2
XFILLER_17_217 vpwr vgnd scs8hd_fill_2
X_530_ _582_/A _529_/X _530_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_345 vgnd vpwr scs8hd_decap_8
XFILLER_17_239 vpwr vgnd scs8hd_fill_2
XFILLER_27_76 vgnd vpwr scs8hd_decap_6
X_461_ _461_/A _462_/A vgnd vpwr scs8hd_buf_1
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XANTENNA__229__A enable vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_423 vgnd vpwr scs8hd_fill_1
X_392_ _392_/A _387_/X _392_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_489 vgnd vpwr scs8hd_decap_12
XFILLER_40_264 vgnd vpwr scs8hd_decap_8
XFILLER_43_75 vpwr vgnd scs8hd_fill_2
XFILLER_43_86 vgnd vpwr scs8hd_decap_3
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_36_515 vgnd vpwr scs8hd_fill_1
XFILLER_63_367 vgnd vpwr scs8hd_decap_4
XFILLER_63_356 vgnd vpwr scs8hd_decap_8
XFILLER_16_250 vpwr vgnd scs8hd_fill_2
XFILLER_31_264 vpwr vgnd scs8hd_fill_2
XFILLER_8_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__602__A _270_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_SLEEPB _481_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_128 vgnd vpwr scs8hd_decap_4
XFILLER_66_194 vgnd vpwr scs8hd_fill_1
XFILLER_39_397 vgnd vpwr scs8hd_fill_1
XFILLER_22_253 vgnd vpwr scs8hd_decap_4
XFILLER_10_459 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__512__A _523_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XANTENNA__231__B _471_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_415 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_139 vpwr vgnd scs8hd_fill_2
XFILLER_18_504 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_54_41 vgnd vpwr scs8hd_decap_6
XFILLER_45_356 vgnd vpwr scs8hd_decap_4
XFILLER_45_367 vgnd vpwr scs8hd_decap_3
X_513_ _423_/A _505_/X _513_/Y vgnd vpwr scs8hd_nor2_4
X_444_ _466_/A _445_/B _444_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_326 vgnd vpwr scs8hd_decap_6
XFILLER_54_52 vpwr vgnd scs8hd_fill_2
X_375_ _391_/A _376_/B _375_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__406__B _405_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__422__A _457_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_452 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_415 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _638_/HI ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_161 vgnd vpwr scs8hd_decap_4
XFILLER_36_312 vgnd vpwr scs8hd_decap_4
XFILLER_51_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__332__A _391_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_59_426 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_27_301 vpwr vgnd scs8hd_fill_2
XFILLER_54_120 vgnd vpwr scs8hd_decap_3
XFILLER_27_367 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_54_186 vgnd vpwr scs8hd_decap_8
XFILLER_42_359 vgnd vpwr scs8hd_decap_6
XANTENNA__507__A _407_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_234 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _616_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_2_422 vgnd vpwr scs8hd_decap_12
XFILLER_40_98 vpwr vgnd scs8hd_fill_2
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_30 vpwr vgnd scs8hd_fill_2
XFILLER_77_245 vgnd vpwr scs8hd_decap_12
XFILLER_65_407 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_65_51 vgnd vpwr scs8hd_decap_8
XFILLER_58_492 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_65_62 vgnd vpwr scs8hd_decap_6
XFILLER_45_153 vpwr vgnd scs8hd_fill_2
XFILLER_18_389 vpwr vgnd scs8hd_fill_2
XFILLER_33_315 vpwr vgnd scs8hd_fill_2
XFILLER_45_164 vpwr vgnd scs8hd_fill_2
XFILLER_45_175 vpwr vgnd scs8hd_fill_2
XFILLER_45_197 vgnd vpwr scs8hd_decap_6
XANTENNA__417__A _510_/A vgnd vpwr scs8hd_diode_2
X_427_ _409_/A _382_/X _409_/C _471_/D _428_/A vgnd vpwr scs8hd_or4_4
X_358_ address[8] _383_/B _358_/C _409_/D _358_/X vgnd vpwr scs8hd_or4_4
X_289_ _277_/A _593_/A _289_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_293 vgnd vpwr scs8hd_decap_12
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_223 vpwr vgnd scs8hd_fill_2
XFILLER_68_289 vgnd vpwr scs8hd_decap_4
XFILLER_64_462 vgnd vpwr scs8hd_decap_12
XFILLER_36_175 vgnd vpwr scs8hd_decap_6
XFILLER_51_123 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_167 vgnd vpwr scs8hd_decap_4
XANTENNA__327__A _327_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _277_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_510 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_59_201 vgnd vpwr scs8hd_fill_1
XFILLER_59_256 vpwr vgnd scs8hd_fill_2
XFILLER_74_215 vgnd vpwr scs8hd_decap_12
XFILLER_70_421 vgnd vpwr scs8hd_fill_1
XFILLER_27_164 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
XFILLER_82_292 vgnd vpwr scs8hd_decap_12
XPHY_811 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_800 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_76 vpwr vgnd scs8hd_fill_2
XFILLER_42_123 vgnd vpwr scs8hd_decap_8
XPHY_844 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_833 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_822 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_487 vgnd vpwr scs8hd_decap_12
XFILLER_30_318 vpwr vgnd scs8hd_fill_2
XFILLER_35_87 vpwr vgnd scs8hd_fill_2
XANTENNA__237__A address[2] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y _613_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_237 vgnd vpwr scs8hd_decap_4
XFILLER_18_164 vpwr vgnd scs8hd_fill_2
XFILLER_46_462 vgnd vpwr scs8hd_decap_12
XFILLER_61_432 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
XFILLER_33_134 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _248_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_156 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _634_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__610__A _610_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_215 vgnd vpwr scs8hd_decap_4
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XFILLER_56_259 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
XFILLER_20_373 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__504__B _382_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_318 vgnd vpwr scs8hd_decap_12
XANTENNA__520__A _509_/A vgnd vpwr scs8hd_diode_2
XFILLER_75_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_215 vpwr vgnd scs8hd_fill_2
XFILLER_47_237 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_4
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_28_495 vgnd vpwr scs8hd_decap_12
XFILLER_70_240 vpwr vgnd scs8hd_fill_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XFILLER_43_487 vgnd vpwr scs8hd_fill_1
XPHY_652 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_641 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_630 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_696 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_685 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_674 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_663 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_159 vpwr vgnd scs8hd_fill_2
XFILLER_11_384 vgnd vpwr scs8hd_fill_1
XFILLER_11_362 vpwr vgnd scs8hd_fill_2
XFILLER_11_351 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__414__B _422_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ _616_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__430__A _441_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_SLEEPB _389_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_373 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _590_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_440 vpwr vgnd scs8hd_fill_2
XFILLER_34_410 vpwr vgnd scs8hd_fill_2
XFILLER_61_284 vpwr vgnd scs8hd_fill_2
XFILLER_21_126 vpwr vgnd scs8hd_fill_2
XFILLER_21_137 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y _631_/A vgnd vpwr scs8hd_inv_1
XANTENNA__605__A _605_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__340__A _423_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_384 vpwr vgnd scs8hd_fill_2
XFILLER_57_513 vgnd vpwr scs8hd_decap_3
XFILLER_29_204 vpwr vgnd scs8hd_fill_2
XFILLER_44_207 vgnd vpwr scs8hd_decap_6
XFILLER_25_443 vpwr vgnd scs8hd_fill_2
XFILLER_37_270 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_262 vpwr vgnd scs8hd_fill_2
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_487 vgnd vpwr scs8hd_fill_1
XFILLER_40_413 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_468 vgnd vpwr scs8hd_decap_8
XANTENNA__515__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_479 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__250__A _249_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_354 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_398 vgnd vpwr scs8hd_decap_12
XFILLER_73_62 vgnd vpwr scs8hd_decap_12
XFILLER_73_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _640_/HI
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__409__B _382_/X vgnd vpwr scs8hd_diode_2
XFILLER_43_240 vgnd vpwr scs8hd_decap_4
XFILLER_43_284 vpwr vgnd scs8hd_fill_2
XFILLER_43_295 vgnd vpwr scs8hd_decap_4
XFILLER_31_468 vgnd vpwr scs8hd_decap_8
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__425__A _425_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_SLEEPB _350_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_479 vgnd vpwr scs8hd_decap_8
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_163 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_391 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _564_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_229 vgnd vpwr scs8hd_decap_4
XFILLER_81_379 vgnd vpwr scs8hd_decap_12
XFILLER_34_251 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__335__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_306 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_SLEEPB _485_/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_129 vgnd vpwr scs8hd_decap_12
XFILLER_72_379 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
X_460_ _409_/A _471_/B _471_/C _409_/D _461_/A vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_391_ _391_/A _387_/X _391_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_43_21 vgnd vpwr scs8hd_fill_1
XFILLER_9_428 vgnd vpwr scs8hd_decap_12
XANTENNA__245__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_287 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _564_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_118 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_321 vgnd vpwr scs8hd_decap_4
XFILLER_48_332 vgnd vpwr scs8hd_decap_4
XFILLER_63_302 vgnd vpwr scs8hd_fill_1
XFILLER_48_387 vpwr vgnd scs8hd_fill_2
XFILLER_75_184 vgnd vpwr scs8hd_decap_12
XFILLER_48_398 vgnd vpwr scs8hd_decap_4
X_589_ _589_/A _594_/B _589_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_262 vpwr vgnd scs8hd_fill_2
XFILLER_31_210 vpwr vgnd scs8hd_fill_2
XFILLER_76_3 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_298 vgnd vpwr scs8hd_decap_4
XFILLER_8_483 vgnd vpwr scs8hd_decap_12
XANTENNA__602__B _600_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_310 vgnd vpwr scs8hd_fill_1
XFILLER_39_376 vpwr vgnd scs8hd_fill_2
XFILLER_81_110 vgnd vpwr scs8hd_decap_12
XFILLER_54_324 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_SLEEPB _452_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_232 vpwr vgnd scs8hd_fill_2
XFILLER_22_243 vgnd vpwr scs8hd_decap_8
XFILLER_22_265 vgnd vpwr scs8hd_decap_8
XANTENNA__512__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XANTENNA__231__C _515_/C vgnd vpwr scs8hd_diode_2
XFILLER_49_118 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vpwr vgnd scs8hd_fill_2
XFILLER_57_162 vpwr vgnd scs8hd_fill_2
XFILLER_45_302 vgnd vpwr scs8hd_fill_1
XFILLER_57_184 vgnd vpwr scs8hd_decap_4
XFILLER_57_173 vgnd vpwr scs8hd_fill_1
XFILLER_45_313 vpwr vgnd scs8hd_fill_2
XFILLER_45_335 vpwr vgnd scs8hd_fill_2
XFILLER_72_154 vgnd vpwr scs8hd_decap_12
X_512_ _523_/A _511_/B _512_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_379 vpwr vgnd scs8hd_fill_2
X_443_ _454_/A _445_/B _443_/Y vgnd vpwr scs8hd_nor2_4
X_374_ _328_/X _376_/B _374_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_254 vgnd vpwr scs8hd_decap_3
XFILLER_9_214 vgnd vpwr scs8hd_fill_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_12
XFILLER_5_464 vgnd vpwr scs8hd_decap_12
XANTENNA__422__B _422_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_438 vgnd vpwr scs8hd_fill_1
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_76_471 vgnd vpwr scs8hd_decap_12
XFILLER_36_302 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_165 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__613__A _613_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__332__B _322_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_SLEEPB _412_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_405 vpwr vgnd scs8hd_fill_2
XFILLER_67_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_54_110 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_154 vgnd vpwr scs8hd_decap_4
XFILLER_54_143 vgnd vpwr scs8hd_decap_8
XFILLER_54_165 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_45 vgnd vpwr scs8hd_decap_12
XANTENNA__507__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_89 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _538_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_246 vgnd vpwr scs8hd_decap_12
XANTENNA__523__A _523_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _584_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_40_22 vpwr vgnd scs8hd_fill_2
XFILLER_40_77 vgnd vpwr scs8hd_decap_4
XANTENNA__242__B _313_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_434 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_53 vpwr vgnd scs8hd_fill_2
XFILLER_49_75 vpwr vgnd scs8hd_fill_2
XFILLER_77_257 vgnd vpwr scs8hd_decap_12
XFILLER_65_419 vpwr vgnd scs8hd_fill_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_110 vpwr vgnd scs8hd_fill_2
XFILLER_18_346 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_132 vgnd vpwr scs8hd_decap_4
XFILLER_65_96 vpwr vgnd scs8hd_fill_2
XFILLER_60_102 vgnd vpwr scs8hd_decap_3
XFILLER_18_379 vgnd vpwr scs8hd_fill_1
XFILLER_60_124 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_81_62 vgnd vpwr scs8hd_decap_12
XFILLER_81_51 vgnd vpwr scs8hd_decap_8
X_426_ _448_/A _411_/A _426_/Y vgnd vpwr scs8hd_nor2_4
X_357_ address[6] address[7] _358_/C vgnd vpwr scs8hd_or2_4
XFILLER_41_393 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_288_ _288_/A _593_/A vgnd vpwr scs8hd_buf_1
XANTENNA__433__A _466_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _559_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_68_213 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_3 vgnd vpwr scs8hd_decap_4
XFILLER_68_268 vgnd vpwr scs8hd_decap_6
XFILLER_56_419 vgnd vpwr scs8hd_decap_8
XFILLER_64_430 vgnd vpwr scs8hd_fill_1
XFILLER_64_474 vgnd vpwr scs8hd_decap_12
XANTENNA__608__A _608_/A vgnd vpwr scs8hd_diode_2
XFILLER_51_157 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_SLEEPB _372_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_371 vgnd vpwr scs8hd_decap_8
XANTENNA__343__A _425_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_45 vgnd vpwr scs8hd_fill_1
XFILLER_47_408 vpwr vgnd scs8hd_fill_2
XFILLER_74_227 vgnd vpwr scs8hd_decap_4
XFILLER_19_89 vpwr vgnd scs8hd_fill_2
XFILLER_55_441 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_3
XFILLER_27_143 vgnd vpwr scs8hd_decap_4
XFILLER_42_102 vpwr vgnd scs8hd_fill_2
XPHY_801 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_433 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _597_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__518__A _407_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XPHY_845 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_834 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_823 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_812 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_308 vgnd vpwr scs8hd_decap_3
XFILLER_42_157 vgnd vpwr scs8hd_decap_8
XFILLER_70_499 vgnd vpwr scs8hd_decap_12
XFILLER_23_393 vpwr vgnd scs8hd_fill_2
XFILLER_51_32 vpwr vgnd scs8hd_fill_2
XANTENNA__253__A _253_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_98 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_38_408 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vgnd vpwr scs8hd_fill_1
XFILLER_46_474 vgnd vpwr scs8hd_decap_12
XFILLER_73_282 vpwr vgnd scs8hd_fill_2
XANTENNA__428__A _428_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_319 vpwr vgnd scs8hd_fill_2
X_409_ _409_/A _382_/X _409_/C _409_/D _409_/X vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q
+ _361_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_205 vpwr vgnd scs8hd_fill_2
XFILLER_37_452 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_71_208 vgnd vpwr scs8hd_decap_12
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XANTENNA__338__A _404_/A vgnd vpwr scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_24_168 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_507 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__504__C _515_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__520__B _523_/B vgnd vpwr scs8hd_diode_2
XFILLER_46_43 vgnd vpwr scs8hd_decap_8
XFILLER_47_249 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_65 vpwr vgnd scs8hd_fill_2
XANTENNA__248__A _257_/A vgnd vpwr scs8hd_diode_2
XPHY_620 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_146 vgnd vpwr scs8hd_fill_1
XPHY_653 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_642 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_631 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XPHY_686 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_675 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_664 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_697 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_367 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__430__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_78_385 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_inv_1
XFILLER_61_241 vgnd vpwr scs8hd_fill_1
XANTENNA__621__A _621_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_SLEEPB _344_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_1_0_clk/X ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XFILLER_44_219 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_285 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_fill_1
XFILLER_40_425 vgnd vpwr scs8hd_decap_8
XFILLER_32_23 vgnd vpwr scs8hd_decap_6
XANTENNA__515__B _382_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_171 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_337 vgnd vpwr scs8hd_decap_12
XANTENNA__531__A _583_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_57_53 vpwr vgnd scs8hd_fill_2
XFILLER_75_333 vgnd vpwr scs8hd_decap_6
XFILLER_28_271 vpwr vgnd scs8hd_fill_2
XFILLER_73_74 vgnd vpwr scs8hd_decap_12
XANTENNA__409__C _409_/C vgnd vpwr scs8hd_diode_2
XFILLER_43_263 vpwr vgnd scs8hd_fill_2
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_182 vgnd vpwr scs8hd_fill_1
XFILLER_7_175 vgnd vpwr scs8hd_decap_4
XANTENNA__441__A _441_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_66_366 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_414 vgnd vpwr scs8hd_decap_4
XFILLER_34_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__616__A _616_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_296 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__335__B _322_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_480 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XANTENNA__351__A _328_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_318 vgnd vpwr scs8hd_decap_12
XFILLER_69_182 vgnd vpwr scs8hd_fill_1
XFILLER_72_369 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_285 vpwr vgnd scs8hd_fill_2
X_390_ _328_/X _387_/X _390_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__526__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_233 vpwr vgnd scs8hd_fill_2
XFILLER_40_244 vpwr vgnd scs8hd_fill_2
XFILLER_43_55 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_SLEEPB _447_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__261__A _261_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_48_377 vgnd vpwr scs8hd_fill_1
XFILLER_75_196 vgnd vpwr scs8hd_decap_12
XFILLER_63_347 vpwr vgnd scs8hd_fill_2
X_588_ _581_/A _594_/B vgnd vpwr scs8hd_buf_1
XFILLER_71_380 vgnd vpwr scs8hd_decap_4
XANTENNA__436__A _447_/A vgnd vpwr scs8hd_diode_2
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _266_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_69_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_495 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ _522_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _559_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_66_163 vgnd vpwr scs8hd_decap_8
XFILLER_66_174 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_509 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ _479_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__346__A address[8] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ _436_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__231__D _515_/D vgnd vpwr scs8hd_diode_2
XFILLER_77_428 vgnd vpwr scs8hd_decap_12
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_11 vpwr vgnd scs8hd_fill_2
XFILLER_38_22 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_141 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_SLEEPB _405_/Y vgnd vpwr scs8hd_diode_2
X_511_ _522_/A _511_/B _511_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_166 vgnd vpwr scs8hd_decap_12
X_442_ _442_/A _445_/B _442_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ _379_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_76 vpwr vgnd scs8hd_fill_2
XFILLER_53_380 vpwr vgnd scs8hd_fill_2
XANTENNA__256__A _255_/X vgnd vpwr scs8hd_diode_2
X_373_ _325_/X _376_/B _373_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_299 vgnd vpwr scs8hd_decap_4
XFILLER_79_62 vgnd vpwr scs8hd_decap_12
XFILLER_79_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _609_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _644_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_483 vgnd vpwr scs8hd_decap_12
XFILLER_36_347 vgnd vpwr scs8hd_decap_8
XFILLER_51_317 vpwr vgnd scs8hd_fill_2
XFILLER_63_199 vpwr vgnd scs8hd_fill_2
XFILLER_51_339 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q
+ _497_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q
+ _454_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_439 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_409 vgnd vpwr scs8hd_decap_12
XFILLER_67_450 vpwr vgnd scs8hd_fill_2
XFILLER_39_130 vgnd vpwr scs8hd_decap_4
XFILLER_67_483 vgnd vpwr scs8hd_decap_4
XFILLER_54_133 vgnd vpwr scs8hd_fill_1
XFILLER_27_347 vpwr vgnd scs8hd_fill_2
XFILLER_27_358 vgnd vpwr scs8hd_decap_6
XFILLER_82_497 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q
+ _402_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_380 vpwr vgnd scs8hd_fill_2
XFILLER_50_361 vpwr vgnd scs8hd_fill_2
XFILLER_50_372 vpwr vgnd scs8hd_fill_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_3
XFILLER_24_79 vgnd vpwr scs8hd_decap_4
XFILLER_10_258 vgnd vpwr scs8hd_decap_12
XANTENNA__523__B _523_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_45 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_SLEEPB _367_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_89 vgnd vpwr scs8hd_decap_3
XFILLER_2_446 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ _353_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_77_269 vgnd vpwr scs8hd_decap_12
XFILLER_58_450 vpwr vgnd scs8hd_fill_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_314 vgnd vpwr scs8hd_decap_4
XFILLER_73_431 vpwr vgnd scs8hd_fill_2
XFILLER_18_358 vpwr vgnd scs8hd_fill_2
XFILLER_18_369 vpwr vgnd scs8hd_fill_2
XFILLER_26_391 vgnd vpwr scs8hd_decap_6
X_425_ _425_/A _448_/A vgnd vpwr scs8hd_buf_1
XFILLER_81_74 vgnd vpwr scs8hd_decap_12
X_356_ _395_/A _356_/B _356_/Y vgnd vpwr scs8hd_nor2_4
X_287_ _278_/X _327_/A _288_/A vgnd vpwr scs8hd_or2_4
XANTENNA__433__B _429_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_SLEEPB _501_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_236 vpwr vgnd scs8hd_fill_2
XFILLER_56_409 vgnd vpwr scs8hd_fill_1
XFILLER_49_461 vpwr vgnd scs8hd_fill_2
XFILLER_64_442 vpwr vgnd scs8hd_fill_2
XFILLER_64_486 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_114 vpwr vgnd scs8hd_fill_2
XFILLER_24_328 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_147 vgnd vpwr scs8hd_decap_4
XANTENNA__624__A _624_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_269 vpwr vgnd scs8hd_fill_2
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_82_261 vgnd vpwr scs8hd_decap_12
XFILLER_55_475 vgnd vpwr scs8hd_decap_12
XFILLER_15_317 vpwr vgnd scs8hd_fill_2
XFILLER_15_306 vpwr vgnd scs8hd_fill_2
XFILLER_35_12 vgnd vpwr scs8hd_fill_1
XFILLER_35_34 vpwr vgnd scs8hd_fill_2
XPHY_802 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__518__B _523_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_114 vpwr vgnd scs8hd_fill_2
XPHY_835 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_824 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_813 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_147 vgnd vpwr scs8hd_decap_6
XFILLER_11_501 vgnd vpwr scs8hd_decap_12
XFILLER_23_361 vgnd vpwr scs8hd_decap_3
XFILLER_23_383 vgnd vpwr scs8hd_fill_1
XFILLER_50_180 vgnd vpwr scs8hd_decap_6
XANTENNA__534__A _586_/A vgnd vpwr scs8hd_diode_2
XFILLER_51_77 vpwr vgnd scs8hd_fill_2
XFILLER_51_55 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_217 vgnd vpwr scs8hd_decap_3
XFILLER_46_486 vgnd vpwr scs8hd_decap_12
XFILLER_61_423 vpwr vgnd scs8hd_fill_2
XFILLER_61_489 vgnd vpwr scs8hd_decap_12
X_408_ address[6] _409_/A vgnd vpwr scs8hd_buf_1
XANTENNA__444__A _466_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_SLEEPB _468_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_180 vgnd vpwr scs8hd_decap_3
XFILLER_41_191 vpwr vgnd scs8hd_fill_2
X_339_ _271_/B _423_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XANTENNA__619__A _619_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_431 vpwr vgnd scs8hd_fill_2
XFILLER_37_442 vpwr vgnd scs8hd_fill_2
XFILLER_64_261 vgnd vpwr scs8hd_decap_12
XFILLER_52_401 vpwr vgnd scs8hd_fill_2
XFILLER_37_475 vgnd vpwr scs8hd_fill_1
XFILLER_52_423 vgnd vpwr scs8hd_decap_8
XFILLER_52_412 vpwr vgnd scs8hd_fill_2
XANTENNA__338__B _322_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_114 vpwr vgnd scs8hd_fill_2
XFILLER_37_486 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_12_309 vpwr vgnd scs8hd_fill_2
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XANTENNA__354__A _404_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__504__D _482_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _542_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__529__A _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_453 vgnd vpwr scs8hd_decap_4
XFILLER_55_294 vgnd vpwr scs8hd_decap_4
XFILLER_43_423 vgnd vpwr scs8hd_decap_4
XANTENNA__248__B _583_/A vgnd vpwr scs8hd_diode_2
XPHY_610 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_70_264 vgnd vpwr scs8hd_decap_8
XFILLER_62_32 vgnd vpwr scs8hd_decap_6
XPHY_643 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_632 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_621 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_489 vgnd vpwr scs8hd_decap_12
XPHY_687 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_676 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_665 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_654 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_180 vgnd vpwr scs8hd_fill_1
XFILLER_23_191 vgnd vpwr scs8hd_decap_3
XANTENNA__264__A _242_/A vgnd vpwr scs8hd_diode_2
XPHY_698 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_379 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_SLEEPB _435_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__439__A _438_/X vgnd vpwr scs8hd_diode_2
XFILLER_53_209 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_261 vpwr vgnd scs8hd_fill_2
XFILLER_61_231 vgnd vpwr scs8hd_decap_4
XFILLER_61_264 vgnd vpwr scs8hd_decap_4
XFILLER_21_106 vpwr vgnd scs8hd_fill_2
XFILLER_61_297 vpwr vgnd scs8hd_fill_2
XFILLER_14_180 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_507 vgnd vpwr scs8hd_decap_8
XANTENNA__349__A _314_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_401 vgnd vpwr scs8hd_fill_1
XFILLER_25_423 vpwr vgnd scs8hd_fill_2
XFILLER_37_294 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_489 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_297 vgnd vpwr scs8hd_decap_4
XFILLER_40_448 vgnd vpwr scs8hd_decap_8
XFILLER_32_46 vgnd vpwr scs8hd_decap_8
XANTENNA__515__C _515_/C vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_4
XFILLER_32_79 vgnd vpwr scs8hd_decap_8
XFILLER_4_349 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__531__B _529_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_75_312 vgnd vpwr scs8hd_fill_1
XFILLER_48_515 vgnd vpwr scs8hd_fill_1
XANTENNA__259__A _259_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_412 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _534_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_283 vgnd vpwr scs8hd_decap_4
XFILLER_16_445 vgnd vpwr scs8hd_decap_8
XANTENNA__409__D _409_/D vgnd vpwr scs8hd_diode_2
XFILLER_73_86 vgnd vpwr scs8hd_decap_12
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _641_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__441__B _445_/B vgnd vpwr scs8hd_diode_2
XFILLER_66_312 vgnd vpwr scs8hd_decap_3
XFILLER_66_345 vgnd vpwr scs8hd_decap_4
XFILLER_66_323 vgnd vpwr scs8hd_decap_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_209 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_66_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_283 vgnd vpwr scs8hd_decap_3
XFILLER_34_220 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_448 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y _614_/A vgnd vpwr scs8hd_buf_1
XFILLER_30_492 vgnd vpwr scs8hd_decap_12
XANTENNA__632__A _632_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__351__B _348_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_SLEEPB _522_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_301 vpwr vgnd scs8hd_fill_2
XFILLER_57_378 vgnd vpwr scs8hd_fill_1
XFILLER_72_337 vgnd vpwr scs8hd_decap_4
XFILLER_72_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_46 vpwr vgnd scs8hd_fill_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _633_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_404 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _583_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_426 vgnd vpwr scs8hd_fill_1
XFILLER_25_297 vpwr vgnd scs8hd_fill_2
XANTENNA__526__B address[7] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ _490_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__542__A _594_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ _447_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_345 vgnd vpwr scs8hd_decap_4
XFILLER_63_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_587_ _587_/A _587_/B _587_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__436__B _429_/A vgnd vpwr scs8hd_diode_2
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ _395_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _589_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__452__A _441_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_39_323 vpwr vgnd scs8hd_fill_2
XFILLER_66_131 vgnd vpwr scs8hd_decap_4
XFILLER_66_186 vgnd vpwr scs8hd_decap_8
XFILLER_54_337 vpwr vgnd scs8hd_fill_2
XFILLER_54_304 vpwr vgnd scs8hd_fill_2
XFILLER_81_123 vgnd vpwr scs8hd_decap_12
XFILLER_54_348 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__627__A _627_/A vgnd vpwr scs8hd_diode_2
XANTENNA__346__B _383_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XANTENNA__362__A _325_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_45 vpwr vgnd scs8hd_fill_2
X_510_ _510_/A _511_/B _510_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_89 vgnd vpwr scs8hd_decap_3
XFILLER_45_348 vpwr vgnd scs8hd_fill_2
XFILLER_72_178 vgnd vpwr scs8hd_decap_12
X_441_ _441_/A _445_/B _441_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_318 vpwr vgnd scs8hd_fill_2
XANTENNA__537__A _589_/A vgnd vpwr scs8hd_diode_2
X_372_ _314_/X _376_/B _372_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_234 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_70_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_278 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__272__A _271_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_495 vgnd vpwr scs8hd_decap_12
XFILLER_63_112 vpwr vgnd scs8hd_fill_2
XFILLER_63_123 vgnd vpwr scs8hd_decap_4
XFILLER_36_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__447__A _447_/A vgnd vpwr scs8hd_diode_2
X_639_ _639_/HI _639_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_81_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_418 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_326 vgnd vpwr scs8hd_decap_6
XFILLER_39_164 vpwr vgnd scs8hd_fill_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_197 vgnd vpwr scs8hd_decap_4
XANTENNA__357__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_42_329 vpwr vgnd scs8hd_fill_2
XFILLER_58_440 vgnd vpwr scs8hd_fill_1
XFILLER_49_99 vgnd vpwr scs8hd_decap_6
XFILLER_73_487 vgnd vpwr scs8hd_fill_1
XANTENNA__267__A _301_/A vgnd vpwr scs8hd_diode_2
XFILLER_60_137 vpwr vgnd scs8hd_fill_2
X_424_ _447_/A _411_/A _424_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_81_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_355_ _340_/X _356_/B _355_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
X_286_ _286_/A _286_/B address[1] _327_/A vgnd vpwr scs8hd_or3_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_215 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_134 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_145 vgnd vpwr scs8hd_decap_8
XFILLER_64_498 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_237 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_454 vgnd vpwr scs8hd_decap_4
XFILLER_35_24 vgnd vpwr scs8hd_fill_1
XFILLER_82_273 vgnd vpwr scs8hd_decap_6
XFILLER_70_413 vgnd vpwr scs8hd_decap_8
XFILLER_55_487 vgnd vpwr scs8hd_fill_1
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XPHY_836 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_825 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_814 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_803 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_457 vgnd vpwr scs8hd_fill_1
XFILLER_11_513 vgnd vpwr scs8hd_decap_3
XANTENNA__534__B _529_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__550__A _270_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_2_288 vgnd vpwr scs8hd_decap_12
XFILLER_46_432 vgnd vpwr scs8hd_decap_6
XFILLER_73_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XFILLER_33_115 vpwr vgnd scs8hd_fill_2
XFILLER_46_498 vgnd vpwr scs8hd_decap_12
XFILLER_61_468 vgnd vpwr scs8hd_decap_12
XFILLER_14_340 vpwr vgnd scs8hd_fill_2
X_407_ _407_/A _441_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA__444__B _445_/B vgnd vpwr scs8hd_diode_2
X_338_ _404_/A _322_/X _338_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_395 vpwr vgnd scs8hd_fill_2
X_269_ _268_/X _270_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _648_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__460__A _409_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_465 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_273 vpwr vgnd scs8hd_fill_2
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__635__A _635_/A vgnd vpwr scs8hd_diode_2
XANTENNA__354__B _348_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_332 vpwr vgnd scs8hd_fill_2
XFILLER_20_365 vpwr vgnd scs8hd_fill_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_48 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__370__A _369_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _298_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_23 vgnd vpwr scs8hd_decap_3
XFILLER_55_273 vgnd vpwr scs8hd_decap_3
XFILLER_15_115 vgnd vpwr scs8hd_decap_4
XFILLER_43_413 vgnd vpwr scs8hd_decap_4
XFILLER_43_435 vgnd vpwr scs8hd_decap_3
XPHY_611 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_600 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_276 vgnd vpwr scs8hd_decap_4
XFILLER_62_44 vpwr vgnd scs8hd_fill_2
XPHY_644 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_633 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_622 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__545__A _597_/A vgnd vpwr scs8hd_diode_2
XPHY_677 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_666 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_655 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_699 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_688 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__264__B _336_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_387 vgnd vpwr scs8hd_decap_12
XFILLER_11_376 vgnd vpwr scs8hd_decap_8
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__280__A _280_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_218 vpwr vgnd scs8hd_fill_2
XFILLER_78_398 vgnd vpwr scs8hd_decap_12
XFILLER_38_229 vgnd vpwr scs8hd_decap_8
XFILLER_19_465 vpwr vgnd scs8hd_fill_2
XFILLER_46_240 vgnd vpwr scs8hd_decap_4
XFILLER_19_476 vpwr vgnd scs8hd_fill_2
XFILLER_46_273 vpwr vgnd scs8hd_fill_2
XFILLER_34_446 vgnd vpwr scs8hd_decap_12
XFILLER_34_468 vgnd vpwr scs8hd_decap_8
XANTENNA__455__A _466_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_118 vgnd vpwr scs8hd_fill_1
XFILLER_34_479 vgnd vpwr scs8hd_decap_12
XFILLER_14_192 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_332 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__349__B _348_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_52_232 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_254 vpwr vgnd scs8hd_fill_2
XANTENNA__365__A _392_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_479 vgnd vpwr scs8hd_decap_8
XFILLER_40_405 vpwr vgnd scs8hd_fill_2
XANTENNA__515__D _515_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_151 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_77 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XANTENNA__259__B _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_424 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_16_457 vgnd vpwr scs8hd_fill_1
XFILLER_43_232 vpwr vgnd scs8hd_fill_2
XFILLER_73_98 vgnd vpwr scs8hd_decap_12
XFILLER_16_468 vgnd vpwr scs8hd_decap_12
XFILLER_31_405 vgnd vpwr scs8hd_decap_3
XANTENNA__275__A _242_/A vgnd vpwr scs8hd_diode_2
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_188 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_232 vgnd vpwr scs8hd_decap_4
XFILLER_34_243 vpwr vgnd scs8hd_fill_2
XFILLER_34_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_69_184 vgnd vpwr scs8hd_decap_12
XFILLER_57_335 vpwr vgnd scs8hd_fill_2
XFILLER_57_313 vpwr vgnd scs8hd_fill_2
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XFILLER_25_210 vpwr vgnd scs8hd_fill_2
XFILLER_25_254 vpwr vgnd scs8hd_fill_2
XFILLER_40_202 vpwr vgnd scs8hd_fill_2
XANTENNA__526__C _515_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__542__B _542_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_75_110 vgnd vpwr scs8hd_decap_12
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_327 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_390 vgnd vpwr scs8hd_decap_6
X_655_ _655_/HI _655_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_586_ _586_/A _587_/B _586_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XFILLER_16_254 vpwr vgnd scs8hd_fill_2
XFILLER_16_287 vgnd vpwr scs8hd_decap_12
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_268 vpwr vgnd scs8hd_fill_2
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_471 vgnd vpwr scs8hd_decap_12
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_279 vpwr vgnd scs8hd_fill_2
XANTENNA__452__B _456_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_313 vgnd vpwr scs8hd_decap_3
XFILLER_39_346 vgnd vpwr scs8hd_decap_3
XFILLER_81_135 vgnd vpwr scs8hd_decap_12
XFILLER_66_198 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_224 vgnd vpwr scs8hd_decap_8
XANTENNA__346__C _320_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_257 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_22_279 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_290 vpwr vgnd scs8hd_fill_2
XANTENNA__362__B _360_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _551_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_176 vpwr vgnd scs8hd_fill_2
X_440_ _448_/B _445_/B vgnd vpwr scs8hd_buf_1
XFILLER_54_56 vgnd vpwr scs8hd_decap_6
XFILLER_53_360 vgnd vpwr scs8hd_decap_4
XANTENNA__537__B _542_/B vgnd vpwr scs8hd_diode_2
XFILLER_53_393 vgnd vpwr scs8hd_decap_4
X_371_ _378_/B _376_/B vgnd vpwr scs8hd_buf_1
XFILLER_13_213 vpwr vgnd scs8hd_fill_2
XFILLER_80_190 vgnd vpwr scs8hd_decap_12
XFILLER_70_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_217 vgnd vpwr scs8hd_decap_12
XANTENNA__553__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_21_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_489 vgnd vpwr scs8hd_decap_12
XFILLER_79_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_110 vpwr vgnd scs8hd_fill_2
XFILLER_48_121 vpwr vgnd scs8hd_fill_2
XFILLER_36_316 vgnd vpwr scs8hd_fill_1
XFILLER_48_165 vgnd vpwr scs8hd_fill_1
XFILLER_63_135 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_179 vpwr vgnd scs8hd_fill_2
XANTENNA__447__B _448_/B vgnd vpwr scs8hd_diode_2
X_638_ _638_/HI _638_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _645_/HI
+ vgnd vpwr scs8hd_diode_2
X_569_ _294_/X _562_/A _569_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__463__A _441_/A vgnd vpwr scs8hd_diode_2
XFILLER_74_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_54_102 vgnd vpwr scs8hd_decap_8
XFILLER_82_466 vgnd vpwr scs8hd_decap_12
XANTENNA__357__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_190 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__373__A _325_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_58 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _295_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_459 vgnd vpwr scs8hd_decap_12
XFILLER_49_45 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__548__A _547_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_327 vgnd vpwr scs8hd_decap_3
XFILLER_45_157 vpwr vgnd scs8hd_fill_2
XFILLER_45_168 vpwr vgnd scs8hd_fill_2
XFILLER_60_116 vgnd vpwr scs8hd_decap_8
XFILLER_33_319 vpwr vgnd scs8hd_fill_2
XFILLER_45_179 vpwr vgnd scs8hd_fill_2
X_423_ _423_/A _447_/A vgnd vpwr scs8hd_buf_1
XFILLER_53_190 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
X_354_ _404_/A _348_/X _354_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_81_98 vgnd vpwr scs8hd_decap_12
X_285_ _277_/A _592_/A _285_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__283__A _278_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_68_205 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_441 vpwr vgnd scs8hd_fill_2
XFILLER_49_485 vgnd vpwr scs8hd_decap_3
XANTENNA__458__A _447_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_102 vgnd vpwr scs8hd_fill_1
XFILLER_36_124 vgnd vpwr scs8hd_fill_1
XFILLER_17_382 vgnd vpwr scs8hd_decap_4
XFILLER_32_330 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_190 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_216 vpwr vgnd scs8hd_fill_2
XFILLER_59_205 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _262_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_37 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_67_282 vpwr vgnd scs8hd_fill_2
XANTENNA__368__A _395_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_102 vpwr vgnd scs8hd_fill_2
XFILLER_27_113 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _632_/Y vgnd vpwr scs8hd_diode_2
XFILLER_82_230 vgnd vpwr scs8hd_decap_12
XFILLER_27_168 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_70_425 vpwr vgnd scs8hd_fill_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XPHY_826 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_815 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_804 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_837 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_width_0_height_0__pin_12_ vgnd vpwr scs8hd_inv_1
XANTENNA__550__B _548_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_76_32 vgnd vpwr scs8hd_decap_12
XFILLER_65_208 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XANTENNA__278__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_46_411 vpwr vgnd scs8hd_fill_2
XFILLER_18_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_168 vgnd vpwr scs8hd_decap_12
XFILLER_73_274 vpwr vgnd scs8hd_fill_2
XFILLER_61_447 vpwr vgnd scs8hd_fill_2
XFILLER_33_149 vgnd vpwr scs8hd_decap_4
XFILLER_14_363 vgnd vpwr scs8hd_decap_4
X_406_ _395_/A _405_/B _406_/Y vgnd vpwr scs8hd_nor2_4
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _617_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_337_ _523_/A _404_/A vgnd vpwr scs8hd_buf_1
X_268_ _286_/B address[1] _268_/X vgnd vpwr scs8hd_or2_4
XANTENNA__460__B _471_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_6
XFILLER_56_219 vgnd vpwr scs8hd_fill_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_clkbuf_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_400 vpwr vgnd scs8hd_fill_2
XFILLER_49_260 vpwr vgnd scs8hd_fill_2
XFILLER_37_422 vgnd vpwr scs8hd_decap_3
XFILLER_64_241 vgnd vpwr scs8hd_decap_8
XFILLER_64_230 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_190 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _595_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_20_311 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_SLEEPB _392_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_219 vpwr vgnd scs8hd_fill_2
XFILLER_28_433 vpwr vgnd scs8hd_fill_2
XFILLER_28_444 vgnd vpwr scs8hd_decap_3
XFILLER_70_244 vgnd vpwr scs8hd_decap_4
XPHY_601 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_149 vpwr vgnd scs8hd_fill_2
XFILLER_15_127 vgnd vpwr scs8hd_fill_1
XPHY_634 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_623 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_612 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__545__B _528_/X vgnd vpwr scs8hd_diode_2
XPHY_678 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_78 vgnd vpwr scs8hd_decap_12
XFILLER_62_67 vpwr vgnd scs8hd_fill_2
XPHY_667 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_656 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_645 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q
+ _430_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_689 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_399 vgnd vpwr scs8hd_decap_12
XANTENNA__561__A _587_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_300 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q
+ _373_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _603_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_444 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_230 vpwr vgnd scs8hd_fill_2
XFILLER_61_211 vgnd vpwr scs8hd_fill_1
XFILLER_34_414 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__455__B _456_/B vgnd vpwr scs8hd_diode_2
XFILLER_61_288 vgnd vpwr scs8hd_decap_4
XANTENNA__471__A _409_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_208 vpwr vgnd scs8hd_fill_2
XFILLER_69_399 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_SLEEPB _353_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_252 vpwr vgnd scs8hd_fill_2
XFILLER_37_263 vpwr vgnd scs8hd_fill_2
XFILLER_37_274 vpwr vgnd scs8hd_fill_2
XFILLER_52_244 vgnd vpwr scs8hd_fill_1
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_458 vpwr vgnd scs8hd_fill_2
XANTENNA__365__B _360_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_480 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _567_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__381__A _471_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_34 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_358 vgnd vpwr scs8hd_decap_8
XFILLER_28_241 vpwr vgnd scs8hd_fill_2
XANTENNA__259__C _286_/B vgnd vpwr scs8hd_diode_2
XANTENNA__556__A _582_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_222 vgnd vpwr scs8hd_fill_1
XANTENNA__275__B _302_/B vgnd vpwr scs8hd_diode_2
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_439 vpwr vgnd scs8hd_fill_2
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_288 vpwr vgnd scs8hd_fill_2
XFILLER_24_491 vgnd vpwr scs8hd_decap_12
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_SLEEPB _488_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_196 vpwr vgnd scs8hd_fill_2
XANTENNA__291__A _291_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_167 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _642_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_230 vgnd vpwr scs8hd_fill_1
XFILLER_81_306 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _569_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_200 vpwr vgnd scs8hd_fill_2
XANTENNA__466__A _466_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _652_/HI
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_69_130 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_15 vgnd vpwr scs8hd_decap_8
XFILLER_72_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__376__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_361 vgnd vpwr scs8hd_decap_12
XFILLER_25_266 vpwr vgnd scs8hd_fill_2
XFILLER_13_439 vgnd vpwr scs8hd_decap_12
XANTENNA__526__D _482_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_225 vgnd vpwr scs8hd_decap_8
XFILLER_43_25 vpwr vgnd scs8hd_fill_2
XFILLER_43_36 vpwr vgnd scs8hd_fill_2
XFILLER_43_47 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_SLEEPB _455_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_509 vgnd vpwr scs8hd_decap_6
XFILLER_48_358 vgnd vpwr scs8hd_decap_8
XFILLER_48_369 vpwr vgnd scs8hd_fill_2
X_654_ _654_/HI _654_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_233 vgnd vpwr scs8hd_decap_4
XANTENNA__286__A _286_/A vgnd vpwr scs8hd_diode_2
X_585_ _585_/A _587_/B _585_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_70 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_299 vgnd vpwr scs8hd_fill_1
XFILLER_31_214 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_410 vgnd vpwr scs8hd_decap_12
XFILLER_12_483 vgnd vpwr scs8hd_decap_12
XFILLER_39_336 vpwr vgnd scs8hd_fill_2
XFILLER_39_358 vpwr vgnd scs8hd_fill_2
XFILLER_81_147 vgnd vpwr scs8hd_decap_12
XFILLER_62_350 vgnd vpwr scs8hd_decap_4
XANTENNA__346__D _471_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_58 vpwr vgnd scs8hd_fill_2
XFILLER_38_69 vpwr vgnd scs8hd_fill_2
XFILLER_45_317 vgnd vpwr scs8hd_decap_3
X_370_ _369_/X _378_/B vgnd vpwr scs8hd_buf_1
XFILLER_41_501 vgnd vpwr scs8hd_decap_12
XFILLER_9_229 vgnd vpwr scs8hd_decap_12
XFILLER_70_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_SLEEPB _418_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__553__B _552_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _543_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_79_98 vgnd vpwr scs8hd_decap_12
XFILLER_48_133 vgnd vpwr scs8hd_decap_3
XFILLER_63_103 vgnd vpwr scs8hd_decap_6
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XFILLER_36_328 vgnd vpwr scs8hd_decap_8
XFILLER_63_169 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _587_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_309 vpwr vgnd scs8hd_fill_2
X_637_ _637_/HI _637_/LO vgnd vpwr scs8hd_conb_1
X_568_ _594_/A _568_/B _568_/Y vgnd vpwr scs8hd_nor2_4
X_499_ _510_/A _499_/B _499_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__463__B _467_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_67_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_100 vpwr vgnd scs8hd_fill_2
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_27_306 vgnd vpwr scs8hd_decap_3
XFILLER_54_125 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_478 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_350 vgnd vpwr scs8hd_decap_4
XFILLER_23_501 vgnd vpwr scs8hd_decap_12
XFILLER_35_361 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__373__B _376_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_26 vgnd vpwr scs8hd_decap_3
XFILLER_49_57 vpwr vgnd scs8hd_fill_2
XFILLER_49_79 vgnd vpwr scs8hd_decap_4
XFILLER_73_401 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_SLEEPB _375_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_73_423 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_114 vpwr vgnd scs8hd_fill_2
XFILLER_73_489 vgnd vpwr scs8hd_decap_12
X_422_ _457_/A _422_/B _422_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__564__A _590_/A vgnd vpwr scs8hd_diode_2
X_353_ _392_/A _348_/X _353_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_353 vpwr vgnd scs8hd_fill_2
XANTENNA__283__B _324_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_397 vgnd vpwr scs8hd_decap_4
X_284_ _283_/X _592_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q
+ _509_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_93 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q
+ _466_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__458__B _451_/A vgnd vpwr scs8hd_diode_2
XFILLER_51_128 vpwr vgnd scs8hd_fill_2
XANTENNA__474__A _441_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_SLEEPB _509_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_353 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ _420_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _637_/HI ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ _366_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_423 vpwr vgnd scs8hd_fill_2
XANTENNA__368__B _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_82_242 vgnd vpwr scs8hd_decap_6
XFILLER_55_489 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_8
XPHY_827 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_816 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_805 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_459 vpwr vgnd scs8hd_fill_2
XFILLER_70_437 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__384__A _471_/C vgnd vpwr scs8hd_diode_2
XPHY_838 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_36 vpwr vgnd scs8hd_fill_2
XFILLER_23_397 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_78_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_250 vpwr vgnd scs8hd_fill_2
XANTENNA__559__A _585_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_114 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_147 vgnd vpwr scs8hd_decap_4
XFILLER_73_264 vgnd vpwr scs8hd_fill_1
XFILLER_61_415 vpwr vgnd scs8hd_fill_2
XFILLER_61_404 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_73_297 vgnd vpwr scs8hd_decap_4
XFILLER_14_320 vpwr vgnd scs8hd_fill_2
XFILLER_25_81 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_decap_3
X_405_ _340_/X _405_/B _405_/Y vgnd vpwr scs8hd_nor2_4
XPHY_81 vgnd vpwr scs8hd_decap_3
XANTENNA__294__A _294_/A vgnd vpwr scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_decap_3
XFILLER_14_375 vgnd vpwr scs8hd_fill_1
X_336_ _336_/A _523_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q
+ _441_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_267_ _301_/A _277_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_91 vpwr vgnd scs8hd_fill_2
XANTENNA__460__C _471_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_SLEEPB _476_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__469__A _447_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _649_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_209 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q
+ _389_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_49_294 vpwr vgnd scs8hd_fill_2
XFILLER_24_106 vgnd vpwr scs8hd_decap_8
XFILLER_37_478 vgnd vpwr scs8hd_decap_8
XFILLER_37_489 vgnd vpwr scs8hd_decap_12
XFILLER_52_459 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y _634_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_183 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q
+ _329_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_20_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__379__A _395_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_242 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_46_69 vpwr vgnd scs8hd_fill_2
XFILLER_70_223 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XPHY_602 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_635 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_624 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_613 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_668 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_657 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_646 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
XPHY_679 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__561__B _561_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_78_312 vgnd vpwr scs8hd_decap_12
XFILLER_38_209 vgnd vpwr scs8hd_decap_3
XANTENNA__289__A _277_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_401 vgnd vpwr scs8hd_decap_6
XFILLER_19_423 vpwr vgnd scs8hd_fill_2
XFILLER_19_489 vgnd vpwr scs8hd_decap_12
XFILLER_36_91 vgnd vpwr scs8hd_fill_1
XFILLER_61_245 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_161 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_319_ _482_/D _409_/D vgnd vpwr scs8hd_buf_1
XANTENNA__471__B _471_/B vgnd vpwr scs8hd_diode_2
XFILLER_69_301 vpwr vgnd scs8hd_fill_2
XFILLER_69_367 vpwr vgnd scs8hd_fill_2
XFILLER_69_345 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_404 vpwr vgnd scs8hd_fill_2
XFILLER_52_212 vpwr vgnd scs8hd_fill_2
XFILLER_52_267 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_507 vgnd vpwr scs8hd_decap_8
XFILLER_75_304 vgnd vpwr scs8hd_fill_1
XFILLER_57_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_201 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__556__B _561_/B vgnd vpwr scs8hd_diode_2
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_245 vgnd vpwr scs8hd_decap_3
XFILLER_43_267 vpwr vgnd scs8hd_fill_2
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _611_/Y vgnd vpwr scs8hd_diode_2
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_153 vgnd vpwr scs8hd_decap_3
XANTENNA__572__A _304_/B vgnd vpwr scs8hd_diode_2
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_clkbuf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_179 vgnd vpwr scs8hd_fill_1
XFILLER_22_71 vgnd vpwr scs8hd_decap_8
XFILLER_22_82 vpwr vgnd scs8hd_fill_2
XFILLER_22_93 vgnd vpwr scs8hd_decap_4
XFILLER_3_330 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_337 vgnd vpwr scs8hd_decap_4
XFILLER_81_318 vgnd vpwr scs8hd_decap_12
XFILLER_47_90 vpwr vgnd scs8hd_fill_2
XANTENNA__466__B _467_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_510 vgnd vpwr scs8hd_decap_6
XFILLER_19_297 vgnd vpwr scs8hd_decap_3
XFILLER_34_267 vpwr vgnd scs8hd_fill_2
XFILLER_15_470 vgnd vpwr scs8hd_decap_12
XFILLER_22_429 vgnd vpwr scs8hd_decap_3
XFILLER_34_289 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_451 vgnd vpwr scs8hd_decap_6
XANTENNA__482__A _385_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_69_142 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__376__B _376_/B vgnd vpwr scs8hd_diode_2
XFILLER_80_373 vgnd vpwr scs8hd_decap_12
XFILLER_25_289 vgnd vpwr scs8hd_decap_4
XFILLER_40_215 vgnd vpwr scs8hd_fill_1
XFILLER_43_15 vgnd vpwr scs8hd_decap_6
XFILLER_40_248 vgnd vpwr scs8hd_decap_4
XANTENNA__392__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_311 vgnd vpwr scs8hd_decap_12
XFILLER_68_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
XFILLER_75_123 vgnd vpwr scs8hd_decap_12
XFILLER_48_337 vgnd vpwr scs8hd_fill_1
X_653_ _653_/HI _653_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__567__A _593_/A vgnd vpwr scs8hd_diode_2
XANTENNA__286__B _286_/B vgnd vpwr scs8hd_diode_2
X_584_ _584_/A _587_/B _584_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_362 vpwr vgnd scs8hd_fill_2
XFILLER_16_267 vpwr vgnd scs8hd_fill_2
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_237 vpwr vgnd scs8hd_fill_2
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_422 vgnd vpwr scs8hd_decap_12
XFILLER_12_495 vgnd vpwr scs8hd_decap_12
XFILLER_33_81 vpwr vgnd scs8hd_fill_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_79_440 vgnd vpwr scs8hd_decap_12
XFILLER_39_304 vgnd vpwr scs8hd_fill_1
XFILLER_66_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XANTENNA__477__A _466_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_370 vpwr vgnd scs8hd_fill_2
XFILLER_81_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_204 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ _502_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_26 vgnd vpwr scs8hd_decap_3
XFILLER_57_123 vgnd vpwr scs8hd_decap_3
XANTENNA__387__A _387_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ _459_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_513 vgnd vpwr scs8hd_decap_3
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_70_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_403 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _534_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_410 vgnd vpwr scs8hd_decap_12
XANTENNA__297__A _297_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_145 vgnd vpwr scs8hd_decap_8
XFILLER_48_178 vpwr vgnd scs8hd_fill_2
XFILLER_48_189 vgnd vpwr scs8hd_decap_8
XFILLER_63_148 vgnd vpwr scs8hd_decap_6
X_636_ _636_/HI _636_/LO vgnd vpwr scs8hd_conb_1
X_567_ _593_/A _568_/B _567_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_373 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_498_ _509_/A _499_/B _498_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _646_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_79_281 vgnd vpwr scs8hd_decap_12
XFILLER_67_421 vpwr vgnd scs8hd_fill_2
XFILLER_67_454 vpwr vgnd scs8hd_fill_2
XFILLER_39_145 vpwr vgnd scs8hd_fill_2
XFILLER_82_435 vgnd vpwr scs8hd_decap_12
XFILLER_67_487 vgnd vpwr scs8hd_fill_1
XFILLER_54_137 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y _606_/A vgnd vpwr scs8hd_buf_1
XFILLER_35_384 vpwr vgnd scs8hd_fill_2
XFILLER_50_376 vpwr vgnd scs8hd_fill_2
XFILLER_50_398 vgnd vpwr scs8hd_decap_8
XFILLER_10_218 vpwr vgnd scs8hd_fill_2
XFILLER_40_16 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_443 vgnd vpwr scs8hd_decap_4
XFILLER_58_454 vgnd vpwr scs8hd_decap_4
XFILLER_73_435 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_79 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_107 vgnd vpwr scs8hd_decap_6
X_421_ _523_/A _457_/A vgnd vpwr scs8hd_buf_1
X_352_ _391_/A _348_/X _352_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__564__B _568_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_332 vgnd vpwr scs8hd_decap_4
XFILLER_41_376 vpwr vgnd scs8hd_fill_2
X_283_ _278_/X _324_/A _283_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _625_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__580__A _579_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_3
XFILLER_49_421 vgnd vpwr scs8hd_decap_4
XFILLER_76_251 vgnd vpwr scs8hd_decap_8
XFILLER_49_454 vgnd vpwr scs8hd_decap_4
XFILLER_49_465 vgnd vpwr scs8hd_decap_12
XFILLER_64_402 vgnd vpwr scs8hd_decap_6
XFILLER_64_446 vpwr vgnd scs8hd_fill_2
XFILLER_51_118 vpwr vgnd scs8hd_fill_2
XFILLER_17_362 vpwr vgnd scs8hd_fill_2
X_619_ _619_/A _619_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__474__B _476_/B vgnd vpwr scs8hd_diode_2
XANTENNA__490__A _523_/A vgnd vpwr scs8hd_diode_2
XFILLER_67_240 vpwr vgnd scs8hd_fill_2
XFILLER_67_273 vgnd vpwr scs8hd_decap_3
XFILLER_55_413 vgnd vpwr scs8hd_decap_3
XFILLER_27_137 vgnd vpwr scs8hd_decap_3
XFILLER_35_16 vpwr vgnd scs8hd_fill_2
XFILLER_70_405 vpwr vgnd scs8hd_fill_2
XFILLER_35_49 vpwr vgnd scs8hd_fill_2
XPHY_817 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_806 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_449 vgnd vpwr scs8hd_decap_8
XFILLER_23_321 vgnd vpwr scs8hd_decap_4
XFILLER_23_332 vpwr vgnd scs8hd_fill_2
XPHY_839 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_828 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_343 vpwr vgnd scs8hd_fill_2
XFILLER_23_354 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_6
XFILLER_23_376 vgnd vpwr scs8hd_decap_4
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_76_56 vgnd vpwr scs8hd_decap_12
XANTENNA__559__B _561_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_262 vpwr vgnd scs8hd_fill_2
XFILLER_58_295 vgnd vpwr scs8hd_decap_3
XFILLER_73_254 vpwr vgnd scs8hd_fill_2
XANTENNA__575__A _575_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_60 vgnd vpwr scs8hd_decap_3
X_404_ _404_/A _404_/B _404_/Y vgnd vpwr scs8hd_nor2_4
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_14_387 vpwr vgnd scs8hd_fill_2
X_335_ _392_/A _322_/X _335_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_151 vpwr vgnd scs8hd_fill_2
XFILLER_41_162 vgnd vpwr scs8hd_decap_4
XPHY_93 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _545_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_195 vpwr vgnd scs8hd_fill_2
X_266_ _257_/A _587_/A _266_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__460__D _409_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__469__B _462_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_240 vpwr vgnd scs8hd_fill_2
XFILLER_37_435 vpwr vgnd scs8hd_fill_2
XFILLER_37_446 vgnd vpwr scs8hd_decap_4
XFILLER_64_276 vgnd vpwr scs8hd_decap_3
XFILLER_52_416 vgnd vpwr scs8hd_decap_4
XFILLER_52_405 vgnd vpwr scs8hd_decap_4
XANTENNA__485__A _407_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_52_438 vgnd vpwr scs8hd_decap_12
XFILLER_24_118 vgnd vpwr scs8hd_fill_1
XFILLER_20_346 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_379 vgnd vpwr scs8hd_fill_1
XFILLER_9_391 vgnd vpwr scs8hd_decap_12
XFILLER_21_29 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__379__B _378_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_402 vgnd vpwr scs8hd_decap_4
XFILLER_46_15 vgnd vpwr scs8hd_decap_8
XFILLER_55_232 vgnd vpwr scs8hd_decap_4
XFILLER_28_457 vgnd vpwr scs8hd_fill_1
XFILLER_70_202 vgnd vpwr scs8hd_decap_12
XFILLER_55_254 vpwr vgnd scs8hd_fill_2
XANTENNA__395__A _395_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_449 vpwr vgnd scs8hd_fill_2
XFILLER_70_257 vgnd vpwr scs8hd_decap_4
XPHY_625 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_614 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_603 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_140 vgnd vpwr scs8hd_decap_6
XPHY_669 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_658 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_647 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_636 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_471 vgnd vpwr scs8hd_decap_12
XFILLER_11_302 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_306 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_324 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__289__B _593_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_210 vgnd vpwr scs8hd_decap_4
XFILLER_46_265 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_287 vgnd vpwr scs8hd_fill_1
XFILLER_61_268 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_91 vgnd vpwr scs8hd_fill_1
X_318_ enable address[5] _482_/D vgnd vpwr scs8hd_nand2_4
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _618_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__471__C _471_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_249_ _249_/A _286_/A _286_/B address[1] _249_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_361 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_6
XFILLER_37_221 vgnd vpwr scs8hd_decap_4
XFILLER_37_287 vgnd vpwr scs8hd_decap_4
XFILLER_37_298 vgnd vpwr scs8hd_decap_4
XFILLER_20_176 vgnd vpwr scs8hd_decap_8
XFILLER_20_187 vpwr vgnd scs8hd_fill_2
XFILLER_0_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_75_316 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_232 vpwr vgnd scs8hd_fill_2
XFILLER_28_254 vpwr vgnd scs8hd_fill_2
XFILLER_28_287 vgnd vpwr scs8hd_fill_1
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_419 vpwr vgnd scs8hd_fill_2
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_SLEEPB _525_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _273_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__572__B _562_/A vgnd vpwr scs8hd_diode_2
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_342 vgnd vpwr scs8hd_decap_12
XFILLER_78_154 vgnd vpwr scs8hd_decap_12
XFILLER_66_327 vgnd vpwr scs8hd_fill_1
XFILLER_74_360 vgnd vpwr scs8hd_decap_8
XFILLER_19_254 vgnd vpwr scs8hd_decap_3
XFILLER_19_265 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _643_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_90 vpwr vgnd scs8hd_fill_2
XFILLER_15_482 vgnd vpwr scs8hd_decap_6
XANTENNA__482__B _382_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _653_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_154 vgnd vpwr scs8hd_decap_12
XFILLER_57_349 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_382 vpwr vgnd scs8hd_fill_2
XFILLER_65_360 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _592_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_224 vgnd vpwr scs8hd_fill_1
XFILLER_80_385 vgnd vpwr scs8hd_decap_12
XFILLER_13_419 vgnd vpwr scs8hd_decap_4
XFILLER_21_452 vpwr vgnd scs8hd_fill_2
XFILLER_21_463 vpwr vgnd scs8hd_fill_2
XANTENNA__392__B _387_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_68 vgnd vpwr scs8hd_decap_12
XFILLER_0_323 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_135 vgnd vpwr scs8hd_decap_12
XFILLER_63_319 vgnd vpwr scs8hd_decap_6
X_652_ _652_/HI _652_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__567__B _568_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_382 vpwr vgnd scs8hd_fill_2
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XFILLER_71_330 vpwr vgnd scs8hd_fill_2
X_583_ _583_/A _587_/B _583_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_83 vgnd vpwr scs8hd_decap_8
XANTENNA__286__C address[1] vgnd vpwr scs8hd_diode_2
XANTENNA__583__A _583_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_430 vpwr vgnd scs8hd_fill_2
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_227 vgnd vpwr scs8hd_decap_8
XFILLER_31_249 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_434 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_452 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_102 vgnd vpwr scs8hd_decap_3
XFILLER_66_135 vgnd vpwr scs8hd_fill_1
XFILLER_54_308 vgnd vpwr scs8hd_fill_1
XANTENNA__477__B _476_/B vgnd vpwr scs8hd_diode_2
XFILLER_74_190 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_393 vgnd vpwr scs8hd_decap_8
XFILLER_62_374 vpwr vgnd scs8hd_fill_2
XANTENNA__493__A _385_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_260 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_102 vpwr vgnd scs8hd_fill_2
XFILLER_38_16 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _589_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_72_105 vgnd vpwr scs8hd_decap_12
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_330 vpwr vgnd scs8hd_fill_2
XFILLER_38_393 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_415 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_76_422 vgnd vpwr scs8hd_decap_12
XANTENNA__578__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_48_102 vgnd vpwr scs8hd_decap_8
XFILLER_36_308 vpwr vgnd scs8hd_fill_2
XFILLER_48_157 vpwr vgnd scs8hd_fill_2
XFILLER_48_168 vgnd vpwr scs8hd_fill_1
XFILLER_63_116 vgnd vpwr scs8hd_decap_6
XFILLER_28_60 vgnd vpwr scs8hd_decap_3
X_635_ _635_/A _635_/Y vgnd vpwr scs8hd_inv_8
XFILLER_44_330 vgnd vpwr scs8hd_decap_4
XFILLER_44_341 vpwr vgnd scs8hd_fill_2
X_566_ _592_/A _568_/B _566_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_171 vgnd vpwr scs8hd_decap_12
X_497_ _413_/A _499_/B _497_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_SLEEPB _329_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_width_0_height_0__pin_11_ vgnd vpwr scs8hd_inv_1
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_79_293 vgnd vpwr scs8hd_decap_12
XFILLER_67_433 vpwr vgnd scs8hd_fill_2
XANTENNA__488__A _510_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_168 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_82_447 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_330 vgnd vpwr scs8hd_decap_4
XFILLER_62_171 vgnd vpwr scs8hd_decap_8
XFILLER_50_311 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _609_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_49_26 vpwr vgnd scs8hd_fill_2
XFILLER_77_208 vgnd vpwr scs8hd_decap_12
XANTENNA__398__A _405_/B vgnd vpwr scs8hd_diode_2
XFILLER_73_414 vpwr vgnd scs8hd_fill_2
XFILLER_73_447 vgnd vpwr scs8hd_decap_12
XFILLER_45_138 vpwr vgnd scs8hd_fill_2
X_420_ _456_/A _422_/B _420_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_352 vgnd vpwr scs8hd_decap_4
X_351_ _328_/X _348_/X _351_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_282_ _286_/A _241_/B _282_/C _324_/A vgnd vpwr scs8hd_or3_4
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_30_61 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_440 vgnd vpwr scs8hd_decap_12
XFILLER_76_263 vpwr vgnd scs8hd_fill_2
XFILLER_36_105 vpwr vgnd scs8hd_fill_2
XFILLER_36_116 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_477 vgnd vpwr scs8hd_decap_8
XFILLER_36_138 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
X_618_ _618_/A _618_/Y vgnd vpwr scs8hd_inv_8
X_549_ _575_/A _548_/X _549_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_366 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__490__B _490_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _563_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_67_230 vpwr vgnd scs8hd_fill_2
XFILLER_82_211 vgnd vpwr scs8hd_decap_6
XFILLER_67_263 vgnd vpwr scs8hd_fill_1
XFILLER_55_458 vgnd vpwr scs8hd_fill_1
XFILLER_27_149 vpwr vgnd scs8hd_fill_2
XPHY_818 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_807 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_829 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_193 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_163 vgnd vpwr scs8hd_decap_8
XFILLER_50_152 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_SLEEPB _442_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_49 vgnd vpwr scs8hd_decap_4
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_76_68 vgnd vpwr scs8hd_decap_12
XANTENNA__575__B _574_/X vgnd vpwr scs8hd_diode_2
XFILLER_61_428 vpwr vgnd scs8hd_fill_2
XFILLER_54_480 vgnd vpwr scs8hd_decap_12
XFILLER_26_171 vgnd vpwr scs8hd_fill_1
X_403_ _392_/A _404_/B _403_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_119 vgnd vpwr scs8hd_decap_3
XFILLER_14_344 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_25_50 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
X_334_ _522_/A _392_/A vgnd vpwr scs8hd_buf_1
XPHY_94 vgnd vpwr scs8hd_decap_3
XANTENNA__591__A _591_/A vgnd vpwr scs8hd_diode_2
X_265_ _264_/X _587_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_281 vgnd vpwr scs8hd_decap_12
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_37_414 vpwr vgnd scs8hd_fill_2
XFILLER_37_469 vgnd vpwr scs8hd_decap_6
XANTENNA__485__B _490_/B vgnd vpwr scs8hd_diode_2
XFILLER_64_299 vgnd vpwr scs8hd_decap_6
XFILLER_64_288 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _650_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_450 vpwr vgnd scs8hd_fill_2
XFILLER_20_303 vpwr vgnd scs8hd_fill_2
XFILLER_20_369 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_SLEEPB _400_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_211 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__395__B _387_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_119 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XPHY_626 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_615 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_604 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_48 vgnd vpwr scs8hd_decap_4
XPHY_659 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_648 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_637 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_483 vgnd vpwr scs8hd_decap_4
XFILLER_23_174 vgnd vpwr scs8hd_decap_6
XFILLER_23_196 vpwr vgnd scs8hd_fill_2
XFILLER_11_358 vpwr vgnd scs8hd_fill_2
XFILLER_7_318 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_513 vgnd vpwr scs8hd_decap_3
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__586__A _586_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_469 vgnd vpwr scs8hd_decap_4
XFILLER_34_406 vgnd vpwr scs8hd_fill_1
XFILLER_46_244 vgnd vpwr scs8hd_fill_1
XFILLER_61_214 vpwr vgnd scs8hd_fill_2
XFILLER_46_299 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _537_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_317_ _380_/A address[7] _320_/C vgnd vpwr scs8hd_or2_4
XFILLER_52_81 vpwr vgnd scs8hd_fill_2
X_248_ _257_/A _583_/A _248_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__471__D _471_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_373 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_69_358 vgnd vpwr scs8hd_decap_8
XFILLER_69_336 vgnd vpwr scs8hd_fill_1
XFILLER_77_391 vgnd vpwr scs8hd_decap_12
XANTENNA__496__A _407_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_480 vgnd vpwr scs8hd_decap_12
XFILLER_25_428 vpwr vgnd scs8hd_fill_2
XFILLER_25_439 vpwr vgnd scs8hd_fill_2
XFILLER_52_258 vpwr vgnd scs8hd_fill_2
XFILLER_52_236 vgnd vpwr scs8hd_decap_8
XFILLER_40_409 vgnd vpwr scs8hd_decap_4
XFILLER_20_100 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_SLEEPB _362_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _558_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_15 vgnd vpwr scs8hd_decap_8
XFILLER_75_306 vgnd vpwr scs8hd_decap_6
XFILLER_68_391 vgnd vpwr scs8hd_decap_6
XFILLER_71_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_472 vgnd vpwr scs8hd_decap_4
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y _611_/A vgnd vpwr scs8hd_inv_1
XFILLER_7_137 vgnd vpwr scs8hd_decap_12
XFILLER_7_159 vpwr vgnd scs8hd_fill_2
XFILLER_3_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_SLEEPB _496_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_166 vgnd vpwr scs8hd_decap_12
XFILLER_66_317 vgnd vpwr scs8hd_decap_3
XFILLER_19_222 vpwr vgnd scs8hd_fill_2
XFILLER_34_236 vgnd vpwr scs8hd_fill_1
XFILLER_34_247 vgnd vpwr scs8hd_decap_4
XFILLER_15_461 vpwr vgnd scs8hd_fill_2
XFILLER_30_442 vpwr vgnd scs8hd_fill_2
XANTENNA__482__C _515_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_69_166 vgnd vpwr scs8hd_decap_12
XFILLER_57_317 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_339 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_29 vpwr vgnd scs8hd_fill_2
XFILLER_53_501 vgnd vpwr scs8hd_decap_12
XFILLER_25_203 vgnd vpwr scs8hd_decap_4
XFILLER_25_214 vpwr vgnd scs8hd_fill_2
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_25_258 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_206 vgnd vpwr scs8hd_decap_8
XFILLER_21_420 vpwr vgnd scs8hd_fill_2
XFILLER_21_431 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_335 vgnd vpwr scs8hd_decap_6
XFILLER_48_317 vpwr vgnd scs8hd_fill_2
XFILLER_48_328 vpwr vgnd scs8hd_fill_2
XFILLER_75_147 vgnd vpwr scs8hd_decap_12
X_651_ _651_/HI _651_/LO vgnd vpwr scs8hd_conb_1
X_582_ _582_/A _587_/B _582_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_203 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XFILLER_16_258 vpwr vgnd scs8hd_fill_2
XFILLER_71_397 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_SLEEPB _463_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__583__B _587_/B vgnd vpwr scs8hd_diode_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_446 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_79_464 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_306 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_501 vgnd vpwr scs8hd_decap_12
XFILLER_47_350 vpwr vgnd scs8hd_fill_2
XFILLER_62_331 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_504 vgnd vpwr scs8hd_decap_12
XANTENNA__493__B _382_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _537_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_114 vpwr vgnd scs8hd_fill_2
XFILLER_57_169 vgnd vpwr scs8hd_decap_4
XFILLER_57_158 vpwr vgnd scs8hd_fill_2
XFILLER_45_309 vpwr vgnd scs8hd_fill_2
XFILLER_72_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_191 vgnd vpwr scs8hd_decap_4
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_397 vgnd vpwr scs8hd_fill_1
XFILLER_13_217 vpwr vgnd scs8hd_fill_2
XFILLER_70_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_SLEEPB _430_/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_434 vgnd vpwr scs8hd_decap_12
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XANTENNA__578__B address[7] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_125 vpwr vgnd scs8hd_fill_2
XFILLER_17_501 vgnd vpwr scs8hd_decap_12
XFILLER_28_83 vgnd vpwr scs8hd_decap_8
X_634_ _634_/A _634_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__594__A _594_/A vgnd vpwr scs8hd_diode_2
XFILLER_44_320 vgnd vpwr scs8hd_decap_3
XFILLER_32_504 vgnd vpwr scs8hd_decap_12
X_565_ _591_/A _568_/B _565_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_71 vgnd vpwr scs8hd_decap_8
X_496_ _407_/A _499_/B _496_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_93 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_471 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _647_/HI
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__488__B _490_/B vgnd vpwr scs8hd_diode_2
XFILLER_67_467 vpwr vgnd scs8hd_fill_2
XFILLER_82_404 vgnd vpwr scs8hd_decap_12
XFILLER_67_489 vgnd vpwr scs8hd_decap_12
XFILLER_82_459 vgnd vpwr scs8hd_decap_6
XFILLER_35_397 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_389 vgnd vpwr scs8hd_decap_8
XFILLER_49_49 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_106 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_459 vgnd vpwr scs8hd_decap_12
XFILLER_65_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_331 vgnd vpwr scs8hd_decap_3
XFILLER_38_180 vgnd vpwr scs8hd_decap_4
XFILLER_14_515 vgnd vpwr scs8hd_fill_1
X_350_ _325_/X _348_/X _350_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_301 vpwr vgnd scs8hd_fill_2
X_281_ _277_/A _591_/A _281_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_30_73 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_30_84 vgnd vpwr scs8hd_decap_8
XANTENNA__589__A _589_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_452 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_242 vgnd vpwr scs8hd_decap_3
XFILLER_49_489 vgnd vpwr scs8hd_decap_12
XFILLER_17_331 vpwr vgnd scs8hd_fill_2
XFILLER_55_70 vpwr vgnd scs8hd_fill_2
X_617_ _617_/A _617_/Y vgnd vpwr scs8hd_inv_8
X_548_ _547_/X _548_/X vgnd vpwr scs8hd_buf_1
XFILLER_32_334 vpwr vgnd scs8hd_fill_2
X_479_ _457_/A _476_/B _479_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_389 vgnd vpwr scs8hd_decap_8
XFILLER_65_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_209 vpwr vgnd scs8hd_fill_2
XANTENNA__499__A _510_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_117 vgnd vpwr scs8hd_decap_3
XFILLER_67_297 vpwr vgnd scs8hd_fill_2
XFILLER_55_437 vpwr vgnd scs8hd_fill_2
XPHY_808 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_429 vpwr vgnd scs8hd_fill_2
XFILLER_23_301 vpwr vgnd scs8hd_fill_2
XFILLER_35_150 vpwr vgnd scs8hd_fill_2
XPHY_819 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_142 vpwr vgnd scs8hd_fill_2
XFILLER_50_131 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _262_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_197 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q
+ _521_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XFILLER_78_507 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_106 vgnd vpwr scs8hd_decap_8
XFILLER_46_415 vgnd vpwr scs8hd_decap_4
XFILLER_73_223 vpwr vgnd scs8hd_fill_2
XFILLER_73_278 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ _478_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_301 vgnd vpwr scs8hd_decap_4
XPHY_40 vgnd vpwr scs8hd_decap_3
X_402_ _391_/A _404_/B _402_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_SLEEPB _395_/Y vgnd vpwr scs8hd_diode_2
XFILLER_54_492 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_26_183 vgnd vpwr scs8hd_fill_1
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_333_ _260_/B _522_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_175 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__591__B _594_/B vgnd vpwr scs8hd_diode_2
X_264_ _242_/A _336_/A _264_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ _435_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_293 vgnd vpwr scs8hd_decap_12
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_404 vgnd vpwr scs8hd_fill_1
XFILLER_49_275 vpwr vgnd scs8hd_fill_2
XFILLER_64_234 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ _378_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_45_481 vgnd vpwr scs8hd_decap_6
XFILLER_17_194 vpwr vgnd scs8hd_fill_2
XFILLER_32_131 vgnd vpwr scs8hd_decap_3
XFILLER_60_462 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_164 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_437 vgnd vpwr scs8hd_decap_4
XFILLER_46_28 vgnd vpwr scs8hd_decap_3
XFILLER_28_459 vgnd vpwr scs8hd_decap_12
XFILLER_70_215 vgnd vpwr scs8hd_decap_4
XFILLER_55_278 vgnd vpwr scs8hd_decap_3
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XPHY_616 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_605 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _608_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q
+ _496_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_649 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_638 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_627 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_315 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q
+ _453_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_SLEEPB _356_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_337 vgnd vpwr scs8hd_decap_12
XANTENNA__586__B _587_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_448 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _570_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_234 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q
+ _401_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_429 vgnd vpwr scs8hd_decap_6
XFILLER_36_72 vgnd vpwr scs8hd_decap_4
XFILLER_61_237 vgnd vpwr scs8hd_decap_4
XFILLER_36_83 vgnd vpwr scs8hd_decap_8
XFILLER_42_462 vgnd vpwr scs8hd_decap_8
XFILLER_42_473 vgnd vpwr scs8hd_decap_12
XFILLER_14_186 vgnd vpwr scs8hd_decap_6
X_316_ address[6] _380_/A vgnd vpwr scs8hd_inv_8
XFILLER_52_93 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_247_ _247_/A _583_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_385 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q
+ _352_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_315 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_SLEEPB _491_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__496__B _499_/B vgnd vpwr scs8hd_diode_2
XFILLER_52_204 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_492 vgnd vpwr scs8hd_decap_12
XFILLER_33_473 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_19 vgnd vpwr scs8hd_fill_1
XFILLER_33_484 vgnd vpwr scs8hd_decap_4
XFILLER_20_134 vgnd vpwr scs8hd_decap_8
XFILLER_20_145 vgnd vpwr scs8hd_decap_4
XFILLER_57_38 vpwr vgnd scs8hd_fill_2
XFILLER_73_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_513 vgnd vpwr scs8hd_decap_3
XFILLER_16_407 vgnd vpwr scs8hd_decap_3
XFILLER_28_267 vpwr vgnd scs8hd_fill_2
XFILLER_43_215 vgnd vpwr scs8hd_decap_4
XFILLER_73_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_259 vpwr vgnd scs8hd_fill_2
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_112 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_178 vpwr vgnd scs8hd_fill_2
XFILLER_7_149 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_178 vgnd vpwr scs8hd_decap_12
XANTENNA__597__A _597_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_370 vpwr vgnd scs8hd_fill_2
XFILLER_34_204 vgnd vpwr scs8hd_decap_8
XFILLER_34_215 vgnd vpwr scs8hd_decap_3
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__482__D _482_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_SLEEPB _458_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _654_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_178 vgnd vpwr scs8hd_decap_4
XANTENNA__300__A _299_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y _626_/A vgnd vpwr scs8hd_buf_1
XFILLER_53_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_29 vpwr vgnd scs8hd_fill_2
XFILLER_80_398 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_487 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _635_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_650_ _650_/HI _650_/LO vgnd vpwr scs8hd_conb_1
X_581_ _581_/A _587_/B vgnd vpwr scs8hd_buf_1
XFILLER_71_343 vpwr vgnd scs8hd_fill_2
XFILLER_71_310 vgnd vpwr scs8hd_decap_3
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XFILLER_16_226 vgnd vpwr scs8hd_fill_1
XFILLER_71_376 vpwr vgnd scs8hd_fill_2
XFILLER_71_354 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XFILLER_79_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_SLEEPB _424_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__493__C _515_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_292 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _281_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_137 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_373 vpwr vgnd scs8hd_fill_2
XFILLER_72_129 vgnd vpwr scs8hd_decap_12
XFILLER_53_343 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_376 vpwr vgnd scs8hd_fill_2
XFILLER_70_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XFILLER_21_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_428 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__578__C _578_/C vgnd vpwr scs8hd_diode_2
XFILLER_76_446 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_17_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_362 vpwr vgnd scs8hd_fill_2
XFILLER_29_373 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_633_ _633_/A _633_/Y vgnd vpwr scs8hd_inv_8
XFILLER_63_129 vgnd vpwr scs8hd_decap_4
XFILLER_56_192 vpwr vgnd scs8hd_fill_2
XANTENNA__594__B _594_/B vgnd vpwr scs8hd_diode_2
X_564_ _590_/A _568_/B _564_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_184 vgnd vpwr scs8hd_decap_12
X_495_ _495_/A _499_/B vgnd vpwr scs8hd_buf_1
XFILLER_44_398 vpwr vgnd scs8hd_fill_2
XFILLER_12_240 vgnd vpwr scs8hd_decap_4
XFILLER_12_273 vpwr vgnd scs8hd_fill_2
XFILLER_60_82 vpwr vgnd scs8hd_fill_2
XFILLER_8_288 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_SLEEPB _378_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ _514_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_115 vgnd vpwr scs8hd_decap_4
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_126 vpwr vgnd scs8hd_fill_2
XFILLER_82_416 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_321 vpwr vgnd scs8hd_fill_2
XFILLER_35_365 vgnd vpwr scs8hd_fill_1
XFILLER_62_195 vgnd vpwr scs8hd_decap_3
XFILLER_50_357 vpwr vgnd scs8hd_fill_2
XFILLER_50_346 vgnd vpwr scs8hd_decap_8
XFILLER_50_368 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_SLEEPB _512_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_65_27 vgnd vpwr scs8hd_decap_12
XFILLER_58_468 vgnd vpwr scs8hd_decap_12
XFILLER_45_118 vpwr vgnd scs8hd_fill_2
XFILLER_81_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_184 vgnd vpwr scs8hd_decap_4
XFILLER_26_387 vpwr vgnd scs8hd_fill_2
XFILLER_81_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_357 vgnd vpwr scs8hd_decap_3
X_280_ _280_/A _591_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_97 vgnd vpwr scs8hd_fill_1
XFILLER_30_41 vgnd vpwr scs8hd_decap_4
XFILLER_5_269 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__589__B _594_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_1_464 vgnd vpwr scs8hd_decap_12
XFILLER_49_413 vpwr vgnd scs8hd_fill_2
XFILLER_39_83 vpwr vgnd scs8hd_fill_2
XFILLER_76_276 vgnd vpwr scs8hd_decap_12
XFILLER_64_427 vgnd vpwr scs8hd_fill_1
XFILLER_17_321 vpwr vgnd scs8hd_fill_2
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
XFILLER_17_343 vgnd vpwr scs8hd_decap_4
XFILLER_29_192 vpwr vgnd scs8hd_fill_2
X_616_ _616_/A _616_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _582_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_547_ _599_/A _526_/X _547_/X vgnd vpwr scs8hd_or2_4
XFILLER_32_302 vpwr vgnd scs8hd_fill_2
XFILLER_44_173 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_478_ _456_/A _476_/B _478_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_379 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ _489_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_390 vgnd vpwr scs8hd_decap_6
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__499__B _499_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ _446_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_254 vpwr vgnd scs8hd_fill_2
XFILLER_55_405 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_809 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ _394_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_SLEEPB _479_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ _344_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y _628_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_276 vpwr vgnd scs8hd_fill_2
XFILLER_58_254 vgnd vpwr scs8hd_decap_8
XFILLER_58_243 vpwr vgnd scs8hd_fill_2
XFILLER_58_287 vgnd vpwr scs8hd_decap_8
XFILLER_18_118 vgnd vpwr scs8hd_decap_8
XFILLER_46_438 vgnd vpwr scs8hd_fill_1
XFILLER_61_408 vpwr vgnd scs8hd_fill_2
XFILLER_61_419 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_25_30 vpwr vgnd scs8hd_fill_2
X_401_ _328_/X _404_/B _401_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_324 vgnd vpwr scs8hd_decap_12
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
X_332_ _391_/A _322_/X _332_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_85 vgnd vpwr scs8hd_fill_1
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_263_ _259_/A _241_/B _282_/C _336_/A vgnd vpwr scs8hd_or3_4
XFILLER_41_187 vpwr vgnd scs8hd_fill_2
XFILLER_41_40 vpwr vgnd scs8hd_fill_2
XFILLER_41_62 vgnd vpwr scs8hd_decap_3
XFILLER_41_95 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_64_202 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_298 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_60_474 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_32_154 vgnd vpwr scs8hd_fill_1
XFILLER_32_187 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _651_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__303__A _302_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_416 vgnd vpwr scs8hd_decap_8
XFILLER_28_449 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_419 vpwr vgnd scs8hd_fill_2
XPHY_617 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_606 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_639 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_628 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_11_327 vgnd vpwr scs8hd_decap_12
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_98 vgnd vpwr scs8hd_decap_8
XFILLER_78_349 vgnd vpwr scs8hd_decap_12
XFILLER_46_257 vpwr vgnd scs8hd_fill_2
XFILLER_36_40 vpwr vgnd scs8hd_fill_2
XFILLER_46_279 vgnd vpwr scs8hd_decap_8
XFILLER_61_227 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_4
X_315_ address[9] _383_/B vgnd vpwr scs8hd_inv_8
XFILLER_42_485 vgnd vpwr scs8hd_decap_12
XFILLER_10_371 vgnd vpwr scs8hd_decap_12
X_246_ _249_/A _286_/A _282_/C _241_/B _247_/A vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _550_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _609_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_419 vpwr vgnd scs8hd_fill_2
XFILLER_33_452 vpwr vgnd scs8hd_fill_2
XFILLER_60_271 vpwr vgnd scs8hd_fill_2
XFILLER_60_293 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ _632_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_224 vgnd vpwr scs8hd_decap_8
XFILLER_73_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_430 vpwr vgnd scs8hd_fill_2
XFILLER_24_441 vgnd vpwr scs8hd_decap_6
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_271 vpwr vgnd scs8hd_fill_2
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_86 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_367 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__597__B _581_/A vgnd vpwr scs8hd_diode_2
XFILLER_59_382 vpwr vgnd scs8hd_fill_2
XFILLER_47_72 vpwr vgnd scs8hd_fill_2
XFILLER_19_279 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
X_229_ enable _230_/A vgnd vpwr scs8hd_inv_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y _617_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_330 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_80_300 vgnd vpwr scs8hd_decap_12
XFILLER_65_352 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_290 vgnd vpwr scs8hd_decap_8
XFILLER_33_260 vgnd vpwr scs8hd_decap_3
XFILLER_68_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_304 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _627_/Y vgnd vpwr scs8hd_diode_2
X_580_ _579_/X _581_/A vgnd vpwr scs8hd_buf_1
XFILLER_56_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_width_0_height_0__pin_10_ vgnd vpwr scs8hd_inv_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_260 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_30 vpwr vgnd scs8hd_fill_2
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_85 vpwr vgnd scs8hd_fill_2
XFILLER_8_459 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__401__A _328_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_319 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_47_374 vpwr vgnd scs8hd_fill_2
XFILLER_15_271 vgnd vpwr scs8hd_decap_4
XFILLER_22_208 vgnd vpwr scs8hd_decap_6
XANTENNA__493__D _515_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__311__A _270_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_330 vgnd vpwr scs8hd_decap_6
XFILLER_26_503 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_352 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y _635_/A vgnd vpwr scs8hd_inv_1
XFILLER_65_182 vgnd vpwr scs8hd_fill_1
XFILLER_53_300 vgnd vpwr scs8hd_decap_3
XFILLER_80_141 vgnd vpwr scs8hd_decap_12
XFILLER_21_252 vpwr vgnd scs8hd_fill_2
XFILLER_79_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA__578__D _482_/D vgnd vpwr scs8hd_diode_2
XFILLER_28_41 vgnd vpwr scs8hd_decap_8
XFILLER_28_52 vgnd vpwr scs8hd_decap_8
XFILLER_28_74 vpwr vgnd scs8hd_fill_2
X_632_ _632_/A _632_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_385 vpwr vgnd scs8hd_fill_2
XFILLER_29_396 vpwr vgnd scs8hd_fill_2
X_563_ _589_/A _568_/B _563_/Y vgnd vpwr scs8hd_nor2_4
X_494_ _494_/A _495_/A vgnd vpwr scs8hd_buf_1
XFILLER_44_377 vgnd vpwr scs8hd_fill_1
XFILLER_71_196 vgnd vpwr scs8hd_decap_12
XFILLER_44_84 vgnd vpwr scs8hd_decap_8
XFILLER_12_285 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_495 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_67_425 vpwr vgnd scs8hd_fill_2
XFILLER_39_149 vpwr vgnd scs8hd_fill_2
XFILLER_82_428 vgnd vpwr scs8hd_decap_6
XFILLER_35_300 vgnd vpwr scs8hd_decap_3
XFILLER_47_171 vgnd vpwr scs8hd_fill_1
XFILLER_62_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_303 vgnd vpwr scs8hd_decap_8
XANTENNA__306__A _305_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_414 vpwr vgnd scs8hd_fill_2
XFILLER_58_436 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_300 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_27 vgnd vpwr scs8hd_decap_12
XFILLER_53_152 vpwr vgnd scs8hd_fill_2
XFILLER_41_336 vgnd vpwr scs8hd_fill_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_20 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_476 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vpwr vgnd scs8hd_fill_2
XFILLER_39_62 vpwr vgnd scs8hd_fill_2
XFILLER_49_458 vgnd vpwr scs8hd_fill_1
XFILLER_76_288 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _576_/Y vgnd vpwr scs8hd_diode_2
X_615_ _615_/A _615_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_72_483 vgnd vpwr scs8hd_decap_12
XFILLER_17_388 vpwr vgnd scs8hd_fill_2
X_546_ _304_/B _528_/X _546_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_152 vgnd vpwr scs8hd_fill_1
XFILLER_44_163 vgnd vpwr scs8hd_decap_8
XFILLER_17_399 vpwr vgnd scs8hd_fill_2
X_477_ _466_/A _476_/B _477_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_409 vpwr vgnd scs8hd_fill_2
XFILLER_35_130 vpwr vgnd scs8hd_fill_2
XFILLER_63_461 vgnd vpwr scs8hd_decap_12
XFILLER_23_336 vpwr vgnd scs8hd_fill_2
XFILLER_23_347 vpwr vgnd scs8hd_fill_2
XFILLER_23_358 vgnd vpwr scs8hd_fill_1
XFILLER_31_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_480 vpwr vgnd scs8hd_fill_2
XFILLER_46_428 vpwr vgnd scs8hd_fill_2
XFILLER_73_258 vgnd vpwr scs8hd_decap_4
XFILLER_73_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_450 vgnd vpwr scs8hd_decap_8
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XFILLER_25_20 vgnd vpwr scs8hd_decap_8
XFILLER_26_163 vgnd vpwr scs8hd_decap_8
X_400_ _325_/X _404_/B _400_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_26_196 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
X_331_ _510_/A _391_/A vgnd vpwr scs8hd_buf_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XFILLER_14_369 vgnd vpwr scs8hd_decap_6
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_41_155 vpwr vgnd scs8hd_fill_2
XFILLER_41_166 vgnd vpwr scs8hd_fill_1
XPHY_86 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XFILLER_41_199 vgnd vpwr scs8hd_fill_1
X_262_ _257_/A _586_/A _262_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_74 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _550_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_49_222 vgnd vpwr scs8hd_decap_3
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_152 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_450 vpwr vgnd scs8hd_fill_2
XFILLER_45_461 vpwr vgnd scs8hd_fill_2
XFILLER_32_100 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_529_ _528_/X _529_/X vgnd vpwr scs8hd_buf_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_486 vgnd vpwr scs8hd_decap_12
XFILLER_20_317 vgnd vpwr scs8hd_decap_8
XFILLER_20_328 vpwr vgnd scs8hd_fill_2
XFILLER_70_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_406 vgnd vpwr scs8hd_fill_1
XFILLER_55_258 vpwr vgnd scs8hd_fill_2
XFILLER_43_409 vpwr vgnd scs8hd_fill_2
XFILLER_63_291 vgnd vpwr scs8hd_decap_4
XPHY_607 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_100 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_629 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_618 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_339 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _636_/HI ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_428 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _582_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_247 vgnd vpwr scs8hd_fill_1
XFILLER_27_450 vgnd vpwr scs8hd_decap_6
XFILLER_36_96 vgnd vpwr scs8hd_decap_6
XFILLER_14_133 vgnd vpwr scs8hd_decap_3
XFILLER_42_442 vpwr vgnd scs8hd_fill_2
XFILLER_52_51 vpwr vgnd scs8hd_fill_2
XFILLER_14_166 vgnd vpwr scs8hd_decap_3
X_314_ _407_/A _314_/X vgnd vpwr scs8hd_buf_1
XFILLER_42_497 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_245_ address[0] _282_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_361 vgnd vpwr scs8hd_decap_4
XFILLER_10_383 vgnd vpwr scs8hd_decap_12
XANTENNA__404__A _404_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _292_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_398 vgnd vpwr scs8hd_decap_12
XFILLER_69_339 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_0_0_clk/X ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_203 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_236 vpwr vgnd scs8hd_fill_2
XFILLER_80_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_228 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_20_103 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__314__A _407_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_258 vgnd vpwr scs8hd_decap_4
XFILLER_73_39 vgnd vpwr scs8hd_decap_12
XFILLER_36_280 vpwr vgnd scs8hd_fill_2
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _595_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_361 vpwr vgnd scs8hd_fill_2
XFILLER_59_350 vpwr vgnd scs8hd_fill_2
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_47_62 vgnd vpwr scs8hd_decap_3
XFILLER_34_239 vgnd vpwr scs8hd_fill_1
XFILLER_15_431 vgnd vpwr scs8hd_decap_4
XFILLER_27_291 vgnd vpwr scs8hd_fill_1
XFILLER_30_412 vgnd vpwr scs8hd_decap_3
XFILLER_42_272 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
X_228_ _578_/C _515_/C vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_309 vpwr vgnd scs8hd_fill_2
XFILLER_80_312 vgnd vpwr scs8hd_decap_12
XFILLER_65_386 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _655_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__309__A _308_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_412 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_467 vgnd vpwr scs8hd_decap_12
XFILLER_21_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_504 vgnd vpwr scs8hd_decap_12
XFILLER_56_386 vpwr vgnd scs8hd_fill_2
XFILLER_16_239 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_412 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_272 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _594_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_434 vgnd vpwr scs8hd_decap_12
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vgnd vpwr scs8hd_decap_8
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _602_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__401__B _404_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_489 vgnd vpwr scs8hd_decap_12
XFILLER_59_180 vgnd vpwr scs8hd_fill_1
XFILLER_62_312 vpwr vgnd scs8hd_fill_2
XFILLER_74_93 vgnd vpwr scs8hd_decap_12
XFILLER_62_334 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_62_389 vgnd vpwr scs8hd_decap_8
XFILLER_62_378 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_790 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_286 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q
+ _372_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__311__B _309_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_106 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _602_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_65_150 vpwr vgnd scs8hd_fill_2
XFILLER_26_515 vgnd vpwr scs8hd_fill_1
XFILLER_53_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_SLEEPB _338_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_286 vpwr vgnd scs8hd_fill_2
XFILLER_21_297 vpwr vgnd scs8hd_fill_2
XFILLER_79_27 vgnd vpwr scs8hd_decap_12
XANTENNA__502__A _423_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_76_459 vgnd vpwr scs8hd_decap_12
XFILLER_63_109 vgnd vpwr scs8hd_fill_1
X_631_ _631_/A _631_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_342 vgnd vpwr scs8hd_decap_4
X_562_ _562_/A _568_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_345 vgnd vpwr scs8hd_decap_4
X_493_ _385_/A _382_/X _515_/C _515_/D _494_/A vgnd vpwr scs8hd_or4_4
XFILLER_44_41 vgnd vpwr scs8hd_decap_8
XFILLER_44_52 vgnd vpwr scs8hd_decap_8
XFILLER_44_389 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_297 vgnd vpwr scs8hd_decap_3
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA__412__A _441_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_220 vgnd vpwr scs8hd_decap_12
XFILLER_67_404 vpwr vgnd scs8hd_fill_2
XFILLER_67_437 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_334 vgnd vpwr scs8hd_fill_1
XFILLER_47_194 vgnd vpwr scs8hd_decap_3
XFILLER_50_315 vgnd vpwr scs8hd_decap_4
XFILLER_35_367 vpwr vgnd scs8hd_fill_2
XANTENNA__322__A _344_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_426 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _568_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_73_418 vgnd vpwr scs8hd_decap_3
XFILLER_26_312 vgnd vpwr scs8hd_decap_4
XFILLER_81_440 vgnd vpwr scs8hd_decap_12
XFILLER_26_356 vgnd vpwr scs8hd_fill_1
XFILLER_53_175 vpwr vgnd scs8hd_fill_2
XFILLER_14_507 vgnd vpwr scs8hd_decap_8
XFILLER_41_315 vpwr vgnd scs8hd_fill_2
XFILLER_81_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_3
XFILLER_30_54 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__232__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_98 vgnd vpwr scs8hd_decap_4
XFILLER_49_437 vpwr vgnd scs8hd_fill_2
XFILLER_76_267 vgnd vpwr scs8hd_decap_8
XFILLER_39_96 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_SLEEPB _445_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_301 vpwr vgnd scs8hd_fill_2
XFILLER_36_109 vgnd vpwr scs8hd_decap_4
X_614_ _614_/A _614_/Y vgnd vpwr scs8hd_inv_8
XFILLER_44_131 vpwr vgnd scs8hd_fill_2
XFILLER_17_367 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_545_ _597_/A _528_/X _545_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _616_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_495 vgnd vpwr scs8hd_decap_12
XFILLER_32_315 vpwr vgnd scs8hd_fill_2
XFILLER_32_326 vpwr vgnd scs8hd_fill_2
XFILLER_32_337 vgnd vpwr scs8hd_fill_1
XFILLER_44_186 vpwr vgnd scs8hd_fill_2
X_476_ _454_/A _476_/B _476_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__407__A _407_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_234 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_278 vpwr vgnd scs8hd_fill_2
XFILLER_27_109 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_473 vgnd vpwr scs8hd_decap_12
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XANTENNA__317__A _380_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _557_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_267 vgnd vpwr scs8hd_decap_6
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XFILLER_26_131 vgnd vpwr scs8hd_decap_4
XFILLER_81_281 vgnd vpwr scs8hd_decap_12
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_54 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vgnd vpwr scs8hd_fill_1
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_41_112 vgnd vpwr scs8hd_decap_4
XFILLER_41_123 vpwr vgnd scs8hd_fill_2
X_330_ _330_/A _510_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_348 vgnd vpwr scs8hd_decap_4
XANTENNA__227__A address[8] vgnd vpwr scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XFILLER_41_134 vpwr vgnd scs8hd_fill_2
XPHY_87 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_decap_3
X_261_ _261_/A _586_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_53 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_SLEEPB _403_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_245 vpwr vgnd scs8hd_fill_2
XFILLER_49_256 vpwr vgnd scs8hd_fill_2
XFILLER_66_72 vgnd vpwr scs8hd_decap_12
XFILLER_64_215 vgnd vpwr scs8hd_decap_4
XFILLER_37_418 vpwr vgnd scs8hd_fill_2
XFILLER_64_237 vgnd vpwr scs8hd_fill_1
XFILLER_60_432 vgnd vpwr scs8hd_decap_4
XFILLER_60_421 vgnd vpwr scs8hd_decap_8
XFILLER_60_454 vgnd vpwr scs8hd_decap_4
X_528_ _527_/X _528_/X vgnd vpwr scs8hd_buf_1
XFILLER_32_145 vgnd vpwr scs8hd_decap_8
X_459_ _448_/A _451_/A _459_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_498 vgnd vpwr scs8hd_decap_12
XFILLER_20_307 vpwr vgnd scs8hd_fill_2
XFILLER_9_330 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _542_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_68_510 vgnd vpwr scs8hd_decap_6
XANTENNA__600__A _599_/X vgnd vpwr scs8hd_diode_2
XFILLER_55_215 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_462 vpwr vgnd scs8hd_fill_2
XFILLER_63_270 vpwr vgnd scs8hd_fill_2
XPHY_608 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_473 vgnd vpwr scs8hd_decap_12
XPHY_619 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_487 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__510__A _510_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_407 vgnd vpwr scs8hd_fill_1
XFILLER_46_226 vpwr vgnd scs8hd_fill_2
XFILLER_61_207 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_SLEEPB _365_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_112 vgnd vpwr scs8hd_decap_3
XFILLER_42_410 vgnd vpwr scs8hd_decap_8
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _311_/Y vgnd vpwr scs8hd_diode_2
X_313_ _313_/A _407_/A vgnd vpwr scs8hd_buf_1
XFILLER_52_85 vgnd vpwr scs8hd_decap_6
X_244_ _257_/A _582_/A _244_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_300 vgnd vpwr scs8hd_decap_12
XFILLER_10_395 vpwr vgnd scs8hd_fill_2
XANTENNA__404__B _404_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__420__A _456_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_340 vgnd vpwr scs8hd_decap_8
XFILLER_77_351 vpwr vgnd scs8hd_fill_2
XFILLER_65_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_248 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y _605_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_259 vpwr vgnd scs8hd_fill_2
XFILLER_52_218 vgnd vpwr scs8hd_decap_8
XFILLER_45_270 vpwr vgnd scs8hd_fill_2
XFILLER_33_432 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_SLEEPB _499_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q
+ _508_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_509 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__330__A _330_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q
+ _465_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_373 vgnd vpwr scs8hd_decap_3
XFILLER_28_237 vpwr vgnd scs8hd_fill_2
XFILLER_51_240 vpwr vgnd scs8hd_fill_2
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q
+ _418_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_51_295 vpwr vgnd scs8hd_fill_2
XFILLER_51_284 vpwr vgnd scs8hd_fill_2
XANTENNA__505__A _504_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_99 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__240__A address[0] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ _365_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_226 vgnd vpwr scs8hd_decap_4
XFILLER_74_343 vgnd vpwr scs8hd_decap_8
XFILLER_19_259 vgnd vpwr scs8hd_decap_6
XFILLER_47_85 vgnd vpwr scs8hd_decap_3
XFILLER_74_398 vgnd vpwr scs8hd_decap_4
XFILLER_63_62 vgnd vpwr scs8hd_decap_3
XFILLER_42_295 vpwr vgnd scs8hd_fill_2
XFILLER_30_457 vgnd vpwr scs8hd_fill_1
XFILLER_30_468 vgnd vpwr scs8hd_decap_12
XANTENNA__415__A _509_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
X_227_ address[8] address[9] _578_/C vgnd vpwr scs8hd_or2_4
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XFILLER_69_126 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_SLEEPB _466_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_8
XFILLER_65_310 vgnd vpwr scs8hd_decap_3
XFILLER_80_324 vgnd vpwr scs8hd_decap_12
XFILLER_65_376 vgnd vpwr scs8hd_decap_4
XFILLER_18_270 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_218 vgnd vpwr scs8hd_decap_6
XFILLER_33_240 vpwr vgnd scs8hd_fill_2
XFILLER_21_424 vgnd vpwr scs8hd_decap_3
XFILLER_21_435 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_479 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__325__A _413_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y _623_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q
+ _388_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_68_181 vgnd vpwr scs8hd_decap_12
XFILLER_56_365 vgnd vpwr scs8hd_decap_8
XFILLER_16_229 vgnd vpwr scs8hd_fill_1
XFILLER_16_218 vgnd vpwr scs8hd_decap_8
XFILLER_16_207 vgnd vpwr scs8hd_decap_6
XFILLER_17_99 vgnd vpwr scs8hd_decap_6
XFILLER_17_66 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_446 vgnd vpwr scs8hd_decap_12
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _540_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q
+ _326_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__235__A address[3] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_66_107 vgnd vpwr scs8hd_decap_3
XFILLER_58_73 vgnd vpwr scs8hd_decap_4
XFILLER_59_170 vpwr vgnd scs8hd_fill_2
XFILLER_58_84 vgnd vpwr scs8hd_decap_8
XFILLER_47_321 vgnd vpwr scs8hd_decap_4
XFILLER_47_354 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_357 vgnd vpwr scs8hd_decap_8
XFILLER_62_346 vpwr vgnd scs8hd_fill_2
XFILLER_62_368 vgnd vpwr scs8hd_decap_4
XFILLER_15_240 vgnd vpwr scs8hd_fill_1
XPHY_780 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_243 vpwr vgnd scs8hd_fill_2
XPHY_791 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_SLEEPB _433_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_118 vpwr vgnd scs8hd_fill_2
XFILLER_38_321 vpwr vgnd scs8hd_fill_2
XFILLER_38_365 vpwr vgnd scs8hd_fill_2
XFILLER_38_398 vgnd vpwr scs8hd_fill_1
XFILLER_80_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_39 vgnd vpwr scs8hd_decap_12
XANTENNA__502__B _495_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_48_129 vpwr vgnd scs8hd_fill_2
XFILLER_56_140 vgnd vpwr scs8hd_decap_6
X_630_ _630_/A _630_/Y vgnd vpwr scs8hd_inv_8
XFILLER_56_173 vpwr vgnd scs8hd_fill_2
X_561_ _587_/A _561_/B _561_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_110 vgnd vpwr scs8hd_decap_12
X_492_ _425_/A _491_/B _492_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_97 vpwr vgnd scs8hd_fill_2
XFILLER_12_265 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__412__B _422_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _532_/Y vgnd vpwr scs8hd_diode_2
XFILLER_79_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_151 vpwr vgnd scs8hd_fill_2
XFILLER_35_346 vpwr vgnd scs8hd_fill_2
XFILLER_47_184 vgnd vpwr scs8hd_fill_1
XFILLER_62_154 vpwr vgnd scs8hd_fill_2
XFILLER_35_357 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__603__A _274_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _610_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y _618_/A vgnd vpwr scs8hd_buf_1
XFILLER_38_140 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_132 vpwr vgnd scs8hd_fill_2
XFILLER_26_346 vgnd vpwr scs8hd_decap_4
XFILLER_81_452 vgnd vpwr scs8hd_decap_12
XFILLER_53_165 vpwr vgnd scs8hd_fill_2
XFILLER_26_368 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_SLEEPB _520_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_349 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XANTENNA__513__A _423_/A vgnd vpwr scs8hd_diode_2
XANTENNA__232__B _231_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_202 vgnd vpwr scs8hd_decap_12
XFILLER_1_489 vgnd vpwr scs8hd_decap_12
XFILLER_64_419 vgnd vpwr scs8hd_decap_8
XFILLER_57_460 vpwr vgnd scs8hd_fill_2
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
X_613_ _613_/A _613_/Y vgnd vpwr scs8hd_inv_8
XFILLER_55_41 vpwr vgnd scs8hd_fill_2
XFILLER_17_335 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vgnd vpwr scs8hd_fill_1
XFILLER_44_110 vgnd vpwr scs8hd_decap_8
XFILLER_55_85 vpwr vgnd scs8hd_fill_2
X_544_ _596_/A _528_/X _544_/Y vgnd vpwr scs8hd_nor2_4
X_475_ _442_/A _476_/B _475_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_501 vgnd vpwr scs8hd_decap_12
XFILLER_32_349 vpwr vgnd scs8hd_fill_2
XFILLER_71_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_51 vgnd vpwr scs8hd_decap_8
XANTENNA__423__A _423_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_55_419 vpwr vgnd scs8hd_fill_2
XFILLER_48_471 vgnd vpwr scs8hd_decap_12
XFILLER_82_249 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_441 vpwr vgnd scs8hd_fill_2
XFILLER_35_154 vpwr vgnd scs8hd_fill_2
XFILLER_63_485 vgnd vpwr scs8hd_decap_3
XFILLER_23_327 vpwr vgnd scs8hd_fill_2
XFILLER_35_198 vpwr vgnd scs8hd_fill_2
XFILLER_50_146 vgnd vpwr scs8hd_decap_6
XFILLER_50_135 vpwr vgnd scs8hd_fill_2
XANTENNA__317__B address[7] vgnd vpwr scs8hd_diode_2
XANTENNA__333__A _260_/B vgnd vpwr scs8hd_diode_2
XFILLER_58_224 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_235 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XFILLER_25_11 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_14_305 vgnd vpwr scs8hd_fill_1
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XANTENNA__508__A _413_/A vgnd vpwr scs8hd_diode_2
XFILLER_81_293 vgnd vpwr scs8hd_decap_12
XFILLER_25_66 vpwr vgnd scs8hd_fill_2
XFILLER_25_88 vpwr vgnd scs8hd_fill_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XANTENNA__227__B address[9] vgnd vpwr scs8hd_diode_2
X_260_ _242_/A _260_/B _261_/A vgnd vpwr scs8hd_or2_4
XPHY_99 vgnd vpwr scs8hd_decap_3
XFILLER_41_10 vpwr vgnd scs8hd_fill_2
XFILLER_6_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ _501_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_49_213 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ _458_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_279 vpwr vgnd scs8hd_fill_2
XFILLER_66_84 vgnd vpwr scs8hd_decap_6
XFILLER_64_249 vgnd vpwr scs8hd_fill_1
XFILLER_57_290 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_411 vgnd vpwr scs8hd_fill_1
XANTENNA__418__A _466_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_165 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_527_ address[4] _526_/X _527_/X vgnd vpwr scs8hd_or2_4
XFILLER_17_198 vpwr vgnd scs8hd_fill_2
XFILLER_82_94 vgnd vpwr scs8hd_decap_12
X_458_ _447_/A _451_/A _458_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_360 vpwr vgnd scs8hd_fill_2
XFILLER_9_342 vgnd vpwr scs8hd_decap_12
X_389_ _325_/X _387_/X _389_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ _406_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _533_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_238 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_430 vgnd vpwr scs8hd_decap_6
XFILLER_70_219 vgnd vpwr scs8hd_fill_1
XFILLER_51_422 vgnd vpwr scs8hd_decap_4
XFILLER_51_400 vpwr vgnd scs8hd_fill_2
XFILLER_23_113 vgnd vpwr scs8hd_decap_3
XANTENNA__328__A _509_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_485 vgnd vpwr scs8hd_decap_12
XPHY_609 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_455 vpwr vgnd scs8hd_fill_2
XFILLER_51_444 vgnd vpwr scs8hd_decap_8
XFILLER_23_157 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__510__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_419 vpwr vgnd scs8hd_fill_2
XFILLER_27_463 vgnd vpwr scs8hd_decap_12
XFILLER_36_32 vgnd vpwr scs8hd_fill_1
XFILLER_36_76 vgnd vpwr scs8hd_fill_1
XANTENNA__238__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_124 vgnd vpwr scs8hd_decap_3
X_312_ _274_/B _309_/X _312_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_64 vpwr vgnd scs8hd_fill_2
X_243_ _243_/A _582_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_312 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_319 vpwr vgnd scs8hd_fill_2
XANTENNA__420__B _422_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_363 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_18_430 vpwr vgnd scs8hd_fill_2
XFILLER_60_230 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_285 vgnd vpwr scs8hd_decap_8
XFILLER_9_172 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__611__A _611_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _624_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_352 vpwr vgnd scs8hd_fill_2
XFILLER_56_514 vpwr vgnd scs8hd_fill_2
XFILLER_43_219 vgnd vpwr scs8hd_fill_1
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_263 vgnd vpwr scs8hd_fill_1
XFILLER_24_455 vgnd vpwr scs8hd_fill_1
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_149 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y _620_/A vgnd vpwr scs8hd_buf_1
XANTENNA__521__A _510_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_105 vgnd vpwr scs8hd_decap_12
XFILLER_59_330 vgnd vpwr scs8hd_fill_1
XFILLER_74_311 vgnd vpwr scs8hd_decap_8
XFILLER_59_374 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_53 vgnd vpwr scs8hd_decap_4
XFILLER_47_97 vpwr vgnd scs8hd_fill_2
XFILLER_74_377 vgnd vpwr scs8hd_decap_12
XFILLER_15_400 vpwr vgnd scs8hd_fill_2
XFILLER_27_271 vgnd vpwr scs8hd_fill_1
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_63_74 vpwr vgnd scs8hd_fill_2
XFILLER_63_52 vgnd vpwr scs8hd_decap_3
XFILLER_15_466 vpwr vgnd scs8hd_fill_2
XFILLER_15_455 vgnd vpwr scs8hd_decap_4
XFILLER_42_252 vgnd vpwr scs8hd_decap_3
XFILLER_30_436 vgnd vpwr scs8hd_decap_4
XFILLER_30_447 vpwr vgnd scs8hd_fill_2
XFILLER_10_160 vpwr vgnd scs8hd_fill_2
X_226_ address[7] _471_/B vgnd vpwr scs8hd_buf_1
XANTENNA__431__A _442_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_503 vgnd vpwr scs8hd_decap_12
XFILLER_77_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_252 vpwr vgnd scs8hd_fill_2
XANTENNA__606__A _606_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_274 vpwr vgnd scs8hd_fill_2
XFILLER_33_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__341__A _340_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_56_311 vpwr vgnd scs8hd_fill_2
XFILLER_56_300 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_193 vgnd vpwr scs8hd_decap_12
XFILLER_17_56 vpwr vgnd scs8hd_fill_2
XFILLER_71_358 vpwr vgnd scs8hd_fill_2
XFILLER_71_347 vpwr vgnd scs8hd_fill_2
XFILLER_17_78 vgnd vpwr scs8hd_decap_3
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__516__A _516_/A vgnd vpwr scs8hd_diode_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _292_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__251__A _257_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_79_403 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_119 vgnd vpwr scs8hd_decap_12
XFILLER_74_141 vgnd vpwr scs8hd_decap_12
XFILLER_59_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_252 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_15_296 vgnd vpwr scs8hd_decap_4
XFILLER_30_222 vgnd vpwr scs8hd_decap_8
XPHY_781 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_770 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__426__A _448_/A vgnd vpwr scs8hd_diode_2
XPHY_792 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_440 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_130 vgnd vpwr scs8hd_decap_4
XFILLER_65_174 vpwr vgnd scs8hd_fill_2
XFILLER_65_163 vgnd vpwr scs8hd_decap_8
XFILLER_38_377 vgnd vpwr scs8hd_decap_3
XFILLER_53_347 vgnd vpwr scs8hd_decap_4
XFILLER_80_166 vgnd vpwr scs8hd_decap_12
XANTENNA__336__A _336_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_130 vgnd vpwr scs8hd_fill_1
X_560_ _586_/A _561_/B _560_/Y vgnd vpwr scs8hd_nor2_4
X_491_ _423_/A _491_/B _491_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_358 vgnd vpwr scs8hd_decap_8
XFILLER_44_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_244 vgnd vpwr scs8hd_fill_1
XANTENNA__246__A _249_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_255 vpwr vgnd scs8hd_fill_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_60_86 vgnd vpwr scs8hd_decap_6
XFILLER_4_410 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_69_62 vgnd vpwr scs8hd_decap_12
XFILLER_69_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_428 vpwr vgnd scs8hd_fill_2
XFILLER_67_417 vpwr vgnd scs8hd_fill_2
XFILLER_39_119 vgnd vpwr scs8hd_fill_1
XFILLER_50_328 vgnd vpwr scs8hd_decap_6
XFILLER_43_391 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _587_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__603__B _600_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_281 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XFILLER_38_163 vgnd vpwr scs8hd_decap_8
XFILLER_53_100 vgnd vpwr scs8hd_decap_3
XFILLER_81_464 vgnd vpwr scs8hd_decap_12
XFILLER_53_144 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _611_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_339 vgnd vpwr scs8hd_fill_1
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XANTENNA__513__B _505_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _636_/HI vgnd vpwr scs8hd_diode_2
XFILLER_49_417 vpwr vgnd scs8hd_fill_2
XFILLER_76_247 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_612_ _612_/A _612_/Y vgnd vpwr scs8hd_inv_8
XFILLER_55_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_325 vgnd vpwr scs8hd_decap_3
XFILLER_29_174 vpwr vgnd scs8hd_fill_2
XFILLER_29_196 vpwr vgnd scs8hd_fill_2
XFILLER_44_122 vpwr vgnd scs8hd_fill_2
XFILLER_17_358 vpwr vgnd scs8hd_fill_2
X_543_ _294_/X _528_/X _543_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_144 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
X_474_ _441_/A _476_/B _474_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_258 vgnd vpwr scs8hd_decap_3
XFILLER_0_490 vgnd vpwr scs8hd_decap_6
XFILLER_55_409 vpwr vgnd scs8hd_fill_2
XFILLER_48_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_483 vgnd vpwr scs8hd_decap_12
XFILLER_50_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_317 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_31_350 vpwr vgnd scs8hd_fill_2
XFILLER_31_361 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__614__A _614_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__508__B _511_/B vgnd vpwr scs8hd_diode_2
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_169 vgnd vpwr scs8hd_decap_3
XFILLER_41_44 vgnd vpwr scs8hd_decap_3
XANTENNA__524__A _423_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_77_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_49_236 vpwr vgnd scs8hd_fill_2
XFILLER_64_206 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_72_272 vgnd vpwr scs8hd_fill_1
XANTENNA__418__B _422_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_526_ _380_/A address[7] _515_/C _482_/D _526_/X vgnd vpwr scs8hd_or4_4
X_457_ _457_/A _456_/B _457_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_388_ _314_/X _387_/X _388_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__434__A _456_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_228 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__609__A _609_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_497 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_51_489 vgnd vpwr scs8hd_decap_12
XANTENNA__344__A _395_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_180 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _633_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_515 vgnd vpwr scs8hd_fill_1
XFILLER_46_206 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_431 vpwr vgnd scs8hd_fill_2
XFILLER_27_442 vpwr vgnd scs8hd_fill_2
XFILLER_36_55 vpwr vgnd scs8hd_fill_2
XFILLER_39_291 vgnd vpwr scs8hd_fill_1
XANTENNA__519__A _413_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_475 vgnd vpwr scs8hd_decap_12
XFILLER_52_32 vpwr vgnd scs8hd_fill_2
X_311_ _270_/B _309_/X _311_/Y vgnd vpwr scs8hd_nor2_4
X_242_ _242_/A _313_/A _243_/A vgnd vpwr scs8hd_or2_4
XFILLER_22_180 vgnd vpwr scs8hd_decap_4
XANTENNA__254__A _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_324 vgnd vpwr scs8hd_decap_12
XFILLER_35_9 vgnd vpwr scs8hd_fill_1
XFILLER_77_62 vgnd vpwr scs8hd_decap_12
XFILLER_77_51 vgnd vpwr scs8hd_decap_8
XFILLER_37_217 vpwr vgnd scs8hd_fill_2
XFILLER_80_507 vgnd vpwr scs8hd_decap_8
XANTENNA__429__A _429_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_423 vpwr vgnd scs8hd_fill_2
XFILLER_33_445 vgnd vpwr scs8hd_decap_4
XFILLER_45_283 vpwr vgnd scs8hd_fill_2
XFILLER_45_294 vpwr vgnd scs8hd_fill_2
X_509_ _509_/A _511_/B _509_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_456 vpwr vgnd scs8hd_fill_2
XFILLER_20_117 vgnd vpwr scs8hd_decap_6
XFILLER_33_489 vgnd vpwr scs8hd_decap_12
XFILLER_13_191 vgnd vpwr scs8hd_decap_4
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_8
XANTENNA__339__A _271_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _251_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__521__B _523_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_301 vgnd vpwr scs8hd_fill_1
XFILLER_59_386 vpwr vgnd scs8hd_fill_2
XFILLER_47_43 vgnd vpwr scs8hd_fill_1
XANTENNA__249__A _249_/A vgnd vpwr scs8hd_diode_2
XFILLER_74_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_423 vpwr vgnd scs8hd_fill_2
XFILLER_27_283 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_242 vpwr vgnd scs8hd_fill_2
XFILLER_42_264 vgnd vpwr scs8hd_decap_8
XFILLER_63_86 vpwr vgnd scs8hd_fill_2
XFILLER_15_489 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XANTENNA__431__B _429_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _625_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_515 vgnd vpwr scs8hd_fill_1
XFILLER_65_356 vpwr vgnd scs8hd_fill_2
XFILLER_18_250 vpwr vgnd scs8hd_fill_2
XFILLER_80_337 vgnd vpwr scs8hd_decap_12
XFILLER_33_231 vgnd vpwr scs8hd_decap_6
XFILLER_33_297 vpwr vgnd scs8hd_fill_2
XFILLER_21_448 vpwr vgnd scs8hd_fill_2
XFILLER_21_459 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__622__A _622_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__341__B _344_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_71_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_SLEEPB _390_/Y vgnd vpwr scs8hd_diode_2
XFILLER_71_326 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_426 vpwr vgnd scs8hd_fill_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_264 vgnd vpwr scs8hd_decap_6
XFILLER_12_459 vgnd vpwr scs8hd_decap_12
XFILLER_33_45 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__532__A _584_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y _629_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_79_415 vgnd vpwr scs8hd_decap_12
XANTENNA__251__B _584_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_64 vpwr vgnd scs8hd_fill_2
XFILLER_47_301 vpwr vgnd scs8hd_fill_2
XFILLER_47_378 vpwr vgnd scs8hd_fill_2
XFILLER_70_370 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vgnd vpwr scs8hd_fill_1
XPHY_771 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_760 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__426__B _411_/A vgnd vpwr scs8hd_diode_2
XPHY_793 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_782 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_256 vpwr vgnd scs8hd_fill_2
XFILLER_30_267 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__442__A _442_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_452 vgnd vpwr scs8hd_decap_12
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_53_315 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_389 vpwr vgnd scs8hd_fill_2
XFILLER_65_197 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_326 vpwr vgnd scs8hd_fill_2
XANTENNA__617__A _617_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ _608_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_245 vgnd vpwr scs8hd_decap_4
XFILLER_21_256 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__352__A _391_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_SLEEPB _351_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_29_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_323 vpwr vgnd scs8hd_fill_2
XFILLER_28_78 vgnd vpwr scs8hd_decap_3
XFILLER_29_367 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _565_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_71_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_44_326 vpwr vgnd scs8hd_fill_2
XFILLER_44_337 vgnd vpwr scs8hd_fill_1
XANTENNA__527__A address[4] vgnd vpwr scs8hd_diode_2
X_490_ _523_/A _490_/B _490_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__246__B _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_60_65 vpwr vgnd scs8hd_fill_2
XFILLER_60_32 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _557_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__262__A _257_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_422 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_69_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_SLEEPB _486_/Y vgnd vpwr scs8hd_diode_2
XFILLER_75_440 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_142 vpwr vgnd scs8hd_fill_2
XFILLER_47_164 vgnd vpwr scs8hd_decap_4
XFILLER_62_123 vgnd vpwr scs8hd_decap_4
XFILLER_35_315 vgnd vpwr scs8hd_decap_4
XFILLER_35_326 vpwr vgnd scs8hd_fill_2
XFILLER_47_175 vpwr vgnd scs8hd_fill_2
XANTENNA__437__A _448_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_370 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_3 vgnd vpwr scs8hd_decap_12
XPHY_590 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_293 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_418 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_66_462 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_304 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_186 vpwr vgnd scs8hd_fill_2
XFILLER_38_197 vgnd vpwr scs8hd_decap_12
XFILLER_81_476 vgnd vpwr scs8hd_decap_12
XANTENNA__347__A _346_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_392 vgnd vpwr scs8hd_decap_4
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_1_403 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_215 vgnd vpwr scs8hd_decap_12
XFILLER_39_55 vgnd vpwr scs8hd_decap_4
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XFILLER_76_259 vgnd vpwr scs8hd_fill_1
X_611_ _611_/A _611_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_153 vgnd vpwr scs8hd_decap_6
XFILLER_55_21 vgnd vpwr scs8hd_fill_1
XFILLER_55_65 vgnd vpwr scs8hd_decap_3
X_542_ _594_/A _542_/B _542_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_473_ _481_/B _476_/B vgnd vpwr scs8hd_buf_1
XANTENNA__257__A _257_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_351 vgnd vpwr scs8hd_decap_4
XFILLER_71_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_SLEEPB _453_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_67_215 vpwr vgnd scs8hd_fill_2
XFILLER_67_226 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _637_/HI vgnd vpwr scs8hd_diode_2
XFILLER_82_218 vgnd vpwr scs8hd_decap_12
XFILLER_35_101 vpwr vgnd scs8hd_fill_2
XFILLER_48_495 vgnd vpwr scs8hd_decap_12
XFILLER_63_454 vgnd vpwr scs8hd_decap_4
XFILLER_35_134 vgnd vpwr scs8hd_decap_3
XFILLER_35_167 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_384 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__630__A _630_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_484 vgnd vpwr scs8hd_decap_4
XFILLER_54_432 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_373 vgnd vpwr scs8hd_decap_6
XFILLER_41_23 vpwr vgnd scs8hd_fill_2
XANTENNA__524__B _517_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_78 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__540__A _592_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_SLEEPB _414_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_421 vpwr vgnd scs8hd_fill_2
XFILLER_17_134 vgnd vpwr scs8hd_decap_3
XFILLER_45_454 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _655_/HI ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_32_104 vpwr vgnd scs8hd_fill_2
XFILLER_45_465 vpwr vgnd scs8hd_fill_2
XFILLER_45_487 vgnd vpwr scs8hd_fill_1
X_525_ _425_/A _517_/A _525_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_82_63 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_126 vgnd vpwr scs8hd_decap_3
X_456_ _456_/A _456_/B _456_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_373 vpwr vgnd scs8hd_fill_2
X_387_ _387_/A _387_/X vgnd vpwr scs8hd_buf_1
XANTENNA__434__B _429_/X vgnd vpwr scs8hd_diode_2
XANTENNA__450__A _450_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _585_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_240 vpwr vgnd scs8hd_fill_2
XFILLER_63_295 vgnd vpwr scs8hd_fill_1
XANTENNA__625__A _625_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_170 vgnd vpwr scs8hd_decap_4
XANTENNA__344__B _344_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XANTENNA__360__A _367_/B vgnd vpwr scs8hd_diode_2
XFILLER_59_513 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_27_410 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__519__B _523_/B vgnd vpwr scs8hd_diode_2
XFILLER_54_262 vpwr vgnd scs8hd_fill_2
XFILLER_27_487 vgnd vpwr scs8hd_fill_1
XFILLER_42_402 vpwr vgnd scs8hd_fill_2
X_310_ _575_/A _309_/X _310_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_457 vgnd vpwr scs8hd_fill_1
XANTENNA__535__A _587_/A vgnd vpwr scs8hd_diode_2
X_241_ _286_/A _241_/B _286_/B _313_/A vgnd vpwr scs8hd_or3_4
XFILLER_52_99 vgnd vpwr scs8hd_decap_6
XANTENNA__254__B _274_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_SLEEPB _373_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_398 vgnd vpwr scs8hd_decap_12
XANTENNA__270__A _259_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_413 vgnd vpwr scs8hd_fill_1
X_508_ _413_/A _511_/B _508_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__445__A _456_/A vgnd vpwr scs8hd_diode_2
X_439_ _438_/X _448_/B vgnd vpwr scs8hd_buf_1
XFILLER_20_107 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _598_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_391 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_SLEEPB _507_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_365 vgnd vpwr scs8hd_decap_6
XFILLER_68_332 vgnd vpwr scs8hd_decap_4
XFILLER_68_398 vgnd vpwr scs8hd_decap_8
XFILLER_68_387 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_402 vpwr vgnd scs8hd_fill_2
XFILLER_51_221 vpwr vgnd scs8hd_fill_2
XFILLER_24_413 vgnd vpwr scs8hd_decap_8
XFILLER_24_424 vgnd vpwr scs8hd_decap_4
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_468 vpwr vgnd scs8hd_fill_2
XFILLER_24_479 vgnd vpwr scs8hd_decap_12
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__355__A _340_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_47 vgnd vpwr scs8hd_decap_12
XFILLER_3_306 vgnd vpwr scs8hd_decap_12
XFILLER_78_129 vgnd vpwr scs8hd_decap_12
XFILLER_59_365 vgnd vpwr scs8hd_fill_1
XFILLER_19_218 vpwr vgnd scs8hd_fill_2
XANTENNA__249__B _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_435 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _257_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__265__A _264_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_276 vgnd vpwr scs8hd_decap_6
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q
+ _520_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_2_361 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q
+ _477_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_80_349 vgnd vpwr scs8hd_decap_12
XFILLER_33_210 vgnd vpwr scs8hd_decap_6
XFILLER_21_416 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_SLEEPB _474_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ _434_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_151 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_47 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ _377_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_243 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_287 vgnd vpwr scs8hd_decap_12
XFILLER_33_68 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__532__B _529_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_32 vpwr vgnd scs8hd_fill_2
XFILLER_47_335 vpwr vgnd scs8hd_fill_2
XFILLER_74_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_327 vgnd vpwr scs8hd_decap_4
XFILLER_62_316 vpwr vgnd scs8hd_fill_2
XFILLER_55_390 vpwr vgnd scs8hd_fill_2
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
XPHY_772 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_761 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_750 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_794 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_783 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__442__B _445_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_464 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q
+ _452_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_78_471 vgnd vpwr scs8hd_decap_12
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_65_187 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q
+ _400_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_61_371 vgnd vpwr scs8hd_decap_3
XANTENNA__633__A _633_/A vgnd vpwr scs8hd_diode_2
XANTENNA__352__B _348_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q
+ _351_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_346 vgnd vpwr scs8hd_fill_1
XFILLER_56_165 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_135 vgnd vpwr scs8hd_decap_12
XANTENNA__527__B _526_/X vgnd vpwr scs8hd_diode_2
XFILLER_52_382 vpwr vgnd scs8hd_fill_2
XFILLER_12_235 vgnd vpwr scs8hd_decap_3
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XANTENNA__246__C _282_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA__543__A _294_/X vgnd vpwr scs8hd_diode_2
XANTENNA__262__B _586_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_434 vgnd vpwr scs8hd_decap_12
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_79_257 vgnd vpwr scs8hd_decap_12
XFILLER_69_86 vgnd vpwr scs8hd_decap_12
XFILLER_75_452 vgnd vpwr scs8hd_decap_12
XANTENNA__437__B _429_/A vgnd vpwr scs8hd_diode_2
XFILLER_70_190 vgnd vpwr scs8hd_decap_12
XPHY_580 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__453__A _442_/A vgnd vpwr scs8hd_diode_2
XPHY_591 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_SLEEPB _448_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_452 vgnd vpwr scs8hd_decap_6
XFILLER_38_154 vpwr vgnd scs8hd_fill_2
XFILLER_66_474 vgnd vpwr scs8hd_decap_12
XANTENNA__628__A _628_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_327 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_179 vgnd vpwr scs8hd_decap_4
XFILLER_41_319 vpwr vgnd scs8hd_fill_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_371 vgnd vpwr scs8hd_decap_8
XFILLER_61_190 vpwr vgnd scs8hd_fill_2
XANTENNA__363__A _328_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_58 vgnd vpwr scs8hd_fill_1
XFILLER_1_415 vgnd vpwr scs8hd_decap_12
XFILLER_39_12 vpwr vgnd scs8hd_fill_2
XFILLER_39_34 vpwr vgnd scs8hd_fill_2
XFILLER_76_227 vgnd vpwr scs8hd_decap_12
XFILLER_57_441 vpwr vgnd scs8hd_fill_2
X_610_ _610_/A _610_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XFILLER_57_485 vgnd vpwr scs8hd_decap_3
XANTENNA__538__A _590_/A vgnd vpwr scs8hd_diode_2
X_541_ _593_/A _542_/B _541_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _560_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_32_319 vpwr vgnd scs8hd_fill_2
X_472_ _471_/X _481_/B vgnd vpwr scs8hd_buf_1
XANTENNA__257__B _585_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_393 vpwr vgnd scs8hd_fill_2
XFILLER_71_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_40_396 vgnd vpwr scs8hd_fill_1
XANTENNA__273__A _277_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_411 vpwr vgnd scs8hd_fill_2
XANTENNA__448__A _448_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XFILLER_16_393 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_SLEEPB _406_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XFILLER_73_208 vgnd vpwr scs8hd_decap_8
XFILLER_39_452 vpwr vgnd scs8hd_fill_2
XFILLER_73_219 vpwr vgnd scs8hd_fill_2
XANTENNA__358__A address[8] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_14_308 vgnd vpwr scs8hd_fill_1
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_179 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_58 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_41_138 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _638_/HI vgnd vpwr scs8hd_diode_2
XFILLER_6_507 vgnd vpwr scs8hd_decap_8
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XANTENNA__540__B _542_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_66_32 vgnd vpwr scs8hd_decap_12
XFILLER_49_249 vpwr vgnd scs8hd_fill_2
XFILLER_17_113 vpwr vgnd scs8hd_fill_2
XANTENNA__268__A _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_45_433 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
X_524_ _423_/A _517_/A _524_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_82_75 vgnd vpwr scs8hd_decap_12
XFILLER_72_285 vgnd vpwr scs8hd_decap_12
X_455_ _466_/A _456_/B _455_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_171 vgnd vpwr scs8hd_fill_1
X_386_ _385_/X _387_/A vgnd vpwr scs8hd_buf_1
XFILLER_13_396 vpwr vgnd scs8hd_fill_2
XFILLER_9_367 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_SLEEPB _368_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_252 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_455 vgnd vpwr scs8hd_fill_1
XFILLER_36_466 vpwr vgnd scs8hd_fill_2
XFILLER_63_274 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ _513_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y _610_/A vgnd vpwr scs8hd_buf_1
XFILLER_39_271 vgnd vpwr scs8hd_fill_1
XFILLER_27_422 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_SLEEPB _502_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_79 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ _470_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_296 vgnd vpwr scs8hd_decap_8
XFILLER_54_285 vpwr vgnd scs8hd_fill_2
XFILLER_54_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_45 vgnd vpwr scs8hd_decap_4
XANTENNA__535__B _529_/X vgnd vpwr scs8hd_diode_2
X_240_ address[0] _286_/B vgnd vpwr scs8hd_inv_8
XFILLER_50_480 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__551__A _274_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_337 vgnd vpwr scs8hd_decap_12
XANTENNA__270__B _270_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_355 vgnd vpwr scs8hd_decap_8
XFILLER_77_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_455 vgnd vpwr scs8hd_fill_1
XFILLER_33_403 vgnd vpwr scs8hd_decap_4
XFILLER_45_241 vgnd vpwr scs8hd_fill_1
XFILLER_60_211 vgnd vpwr scs8hd_fill_1
XFILLER_33_469 vpwr vgnd scs8hd_fill_2
X_507_ _407_/A _511_/B _507_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__445__B _445_/B vgnd vpwr scs8hd_diode_2
X_438_ _385_/A _471_/B _409_/C _409_/D _438_/X vgnd vpwr scs8hd_or4_4
XFILLER_60_299 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vgnd vpwr scs8hd_fill_1
X_369_ address[8] _383_/B _358_/C _471_/D _369_/X vgnd vpwr scs8hd_or4_4
XANTENNA__461__A _461_/A vgnd vpwr scs8hd_diode_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_311 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_506 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_200 vpwr vgnd scs8hd_fill_2
XFILLER_36_285 vpwr vgnd scs8hd_fill_2
XFILLER_51_255 vpwr vgnd scs8hd_fill_2
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q
+ _488_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_51_288 vpwr vgnd scs8hd_fill_2
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
XANTENNA__355__B _356_/B vgnd vpwr scs8hd_diode_2
XFILLER_51_299 vgnd vpwr scs8hd_decap_3
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_480 vgnd vpwr scs8hd_decap_12
XANTENNA__371__A _378_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_59 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_SLEEPB _469_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_318 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _634_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ _445_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_333 vpwr vgnd scs8hd_fill_2
XFILLER_47_23 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_241 vgnd vpwr scs8hd_fill_1
XANTENNA__249__C _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_263 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__546__A _304_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ _393_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_417 vgnd vpwr scs8hd_decap_6
XFILLER_23_480 vpwr vgnd scs8hd_fill_2
XFILLER_42_299 vgnd vpwr scs8hd_decap_4
XFILLER_10_141 vgnd vpwr scs8hd_fill_1
XANTENNA__281__A _277_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ _341_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_373 vgnd vpwr scs8hd_decap_12
XFILLER_77_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _543_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_285 vgnd vpwr scs8hd_decap_3
XANTENNA__456__A _456_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_306 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_SLEEPB _436_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__366__A _404_/A vgnd vpwr scs8hd_diode_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_299 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_79_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_174 vgnd vpwr scs8hd_decap_6
XFILLER_74_166 vgnd vpwr scs8hd_decap_12
XFILLER_74_32 vgnd vpwr scs8hd_decap_12
XFILLER_47_358 vgnd vpwr scs8hd_decap_6
XFILLER_15_211 vgnd vpwr scs8hd_decap_4
XANTENNA__276__A _276_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_762 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_751 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_740 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_288 vpwr vgnd scs8hd_fill_2
XPHY_795 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_784 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_773 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_303 vgnd vpwr scs8hd_decap_3
XFILLER_78_483 vgnd vpwr scs8hd_decap_12
XFILLER_65_100 vgnd vpwr scs8hd_decap_3
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_314 vgnd vpwr scs8hd_decap_4
XFILLER_38_369 vpwr vgnd scs8hd_fill_2
XFILLER_46_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_203 vpwr vgnd scs8hd_fill_2
XFILLER_21_214 vpwr vgnd scs8hd_fill_2
XFILLER_21_225 vpwr vgnd scs8hd_fill_2
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _535_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_358 vpwr vgnd scs8hd_fill_2
XFILLER_56_188 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _654_/HI ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_71_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
XFILLER_52_394 vgnd vpwr scs8hd_decap_3
XANTENNA__246__D _241_/B vgnd vpwr scs8hd_diode_2
XFILLER_44_79 vpwr vgnd scs8hd_fill_2
XFILLER_12_247 vgnd vpwr scs8hd_decap_8
XFILLER_8_207 vgnd vpwr scs8hd_decap_6
XANTENNA__543__B _528_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _608_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y _612_/A vgnd vpwr scs8hd_buf_1
XFILLER_4_446 vgnd vpwr scs8hd_decap_12
XFILLER_69_98 vgnd vpwr scs8hd_decap_12
XFILLER_79_269 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_SLEEPB _523_/Y vgnd vpwr scs8hd_diode_2
XFILLER_75_464 vgnd vpwr scs8hd_decap_12
XFILLER_18_80 vgnd vpwr scs8hd_fill_1
XFILLER_28_380 vgnd vpwr scs8hd_decap_4
XFILLER_28_391 vgnd vpwr scs8hd_decap_6
XFILLER_47_199 vgnd vpwr scs8hd_decap_4
XFILLER_62_158 vgnd vpwr scs8hd_decap_4
XFILLER_31_501 vgnd vpwr scs8hd_decap_12
XFILLER_43_361 vgnd vpwr scs8hd_decap_4
XPHY_570 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__453__B _456_/B vgnd vpwr scs8hd_diode_2
XPHY_592 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_581 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_280 vpwr vgnd scs8hd_fill_2
XFILLER_7_240 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_409 vgnd vpwr scs8hd_decap_3
XFILLER_38_100 vgnd vpwr scs8hd_decap_4
XFILLER_38_144 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_486 vgnd vpwr scs8hd_decap_12
XFILLER_53_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_136 vgnd vpwr scs8hd_decap_8
XFILLER_81_489 vgnd vpwr scs8hd_decap_12
XFILLER_53_169 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XANTENNA__363__B _360_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_3
XFILLER_30_37 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _590_/Y vgnd vpwr scs8hd_diode_2
XFILLER_69_280 vpwr vgnd scs8hd_fill_2
XFILLER_39_79 vpwr vgnd scs8hd_fill_2
XFILLER_57_464 vpwr vgnd scs8hd_fill_2
XFILLER_17_317 vpwr vgnd scs8hd_fill_2
XANTENNA__538__B _542_/B vgnd vpwr scs8hd_diode_2
X_540_ _592_/A _542_/B _540_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_445 vpwr vgnd scs8hd_fill_2
XFILLER_72_434 vgnd vpwr scs8hd_decap_8
XFILLER_72_423 vpwr vgnd scs8hd_fill_2
XFILLER_55_45 vgnd vpwr scs8hd_decap_3
XFILLER_17_339 vpwr vgnd scs8hd_fill_2
XFILLER_55_89 vpwr vgnd scs8hd_fill_2
XFILLER_13_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_471_ _409_/A _471_/B _471_/C _471_/D _471_/X vgnd vpwr scs8hd_or4_4
XANTENNA__554__A _553_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_342 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_40_375 vgnd vpwr scs8hd_decap_8
XFILLER_40_386 vpwr vgnd scs8hd_fill_2
XANTENNA__273__B _589_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ _625_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_423 vpwr vgnd scs8hd_fill_2
XANTENNA__448__B _448_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XFILLER_63_489 vgnd vpwr scs8hd_decap_12
XANTENNA__464__A _442_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_320 vpwr vgnd scs8hd_fill_2
XFILLER_31_331 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _626_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_397 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_206 vgnd vpwr scs8hd_decap_8
XFILLER_58_228 vgnd vpwr scs8hd_decap_4
XFILLER_39_420 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _651_/HI ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_39_442 vpwr vgnd scs8hd_fill_2
XFILLER_66_272 vgnd vpwr scs8hd_fill_1
XFILLER_66_261 vgnd vpwr scs8hd_decap_3
XFILLER_81_220 vgnd vpwr scs8hd_decap_12
XFILLER_26_114 vpwr vgnd scs8hd_fill_2
XANTENNA__358__B _383_/B vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA__374__A _328_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_515 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_44 vgnd vpwr scs8hd_decap_12
XANTENNA__549__A _575_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__268__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_82_32 vgnd vpwr scs8hd_decap_12
XFILLER_72_264 vpwr vgnd scs8hd_fill_2
XFILLER_72_253 vgnd vpwr scs8hd_decap_8
XFILLER_60_404 vgnd vpwr scs8hd_decap_4
X_523_ _523_/A _523_/B _523_/Y vgnd vpwr scs8hd_nor2_4
X_454_ _454_/A _456_/B _454_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_297 vgnd vpwr scs8hd_decap_3
XFILLER_45_489 vgnd vpwr scs8hd_decap_12
XFILLER_82_87 vgnd vpwr scs8hd_decap_6
XANTENNA__284__A _283_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
XFILLER_13_364 vpwr vgnd scs8hd_fill_2
X_385_ _385_/A _382_/X _409_/C _409_/D _385_/X vgnd vpwr scs8hd_or4_4
XFILLER_9_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _639_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__459__A _448_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_401 vgnd vpwr scs8hd_decap_4
XFILLER_36_445 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_SLEEPB _323_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_426 vgnd vpwr scs8hd_fill_1
XFILLER_51_459 vgnd vpwr scs8hd_decap_12
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XANTENNA__369__A address[8] vgnd vpwr scs8hd_diode_2
XFILLER_74_507 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_250 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_36 vpwr vgnd scs8hd_fill_2
XFILLER_39_294 vpwr vgnd scs8hd_fill_2
XFILLER_27_489 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_150 vgnd vpwr scs8hd_decap_3
XFILLER_22_161 vgnd vpwr scs8hd_decap_4
XFILLER_52_68 vpwr vgnd scs8hd_fill_2
XFILLER_50_492 vgnd vpwr scs8hd_decap_12
XFILLER_10_312 vgnd vpwr scs8hd_decap_12
XFILLER_22_194 vgnd vpwr scs8hd_fill_1
XFILLER_10_367 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__551__B _548_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_349 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__279__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_77_367 vgnd vpwr scs8hd_decap_12
XFILLER_77_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_401 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_18_412 vgnd vpwr scs8hd_decap_6
XFILLER_18_434 vpwr vgnd scs8hd_fill_2
X_506_ _505_/X _511_/B vgnd vpwr scs8hd_buf_1
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_437_ _448_/A _429_/A _437_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_110 vgnd vpwr scs8hd_decap_8
X_368_ _395_/A _367_/B _368_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_176 vpwr vgnd scs8hd_fill_2
X_299_ _286_/B address[1] address[3] _259_/A _299_/X vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_245 vgnd vpwr scs8hd_fill_1
XFILLER_51_267 vpwr vgnd scs8hd_fill_2
XFILLER_32_492 vgnd vpwr scs8hd_decap_12
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_59_301 vpwr vgnd scs8hd_fill_2
XFILLER_59_378 vpwr vgnd scs8hd_fill_2
XFILLER_47_35 vpwr vgnd scs8hd_fill_2
XFILLER_74_337 vgnd vpwr scs8hd_decap_3
XFILLER_47_68 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__249__D address[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_404 vgnd vpwr scs8hd_decap_4
XANTENNA__546__B _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_297 vpwr vgnd scs8hd_fill_2
XFILLER_63_78 vgnd vpwr scs8hd_decap_6
XFILLER_30_407 vgnd vpwr scs8hd_decap_3
XANTENNA__562__A _562_/A vgnd vpwr scs8hd_diode_2
XANTENNA__281__B _591_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_385 vgnd vpwr scs8hd_decap_12
XFILLER_65_326 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _301_/Y vgnd vpwr scs8hd_diode_2
XFILLER_73_370 vpwr vgnd scs8hd_fill_2
XFILLER_73_381 vpwr vgnd scs8hd_fill_2
XANTENNA__456__B _456_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_256 vpwr vgnd scs8hd_fill_2
XFILLER_33_278 vpwr vgnd scs8hd_fill_2
XFILLER_33_289 vgnd vpwr scs8hd_decap_3
XANTENNA__472__A _471_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _549_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_315 vgnd vpwr scs8hd_decap_4
XFILLER_56_348 vgnd vpwr scs8hd_decap_8
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_392 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__366__B _360_/X vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_26 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__382__A _382_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_462 vgnd vpwr scs8hd_decap_12
XFILLER_58_56 vgnd vpwr scs8hd_decap_8
XFILLER_58_45 vgnd vpwr scs8hd_decap_8
XFILLER_59_153 vpwr vgnd scs8hd_fill_2
XFILLER_59_197 vgnd vpwr scs8hd_decap_4
XFILLER_74_178 vgnd vpwr scs8hd_decap_12
XFILLER_74_44 vgnd vpwr scs8hd_decap_12
XANTENNA__557__A _583_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_15_223 vpwr vgnd scs8hd_fill_2
XFILLER_70_340 vgnd vpwr scs8hd_decap_8
XFILLER_15_278 vgnd vpwr scs8hd_fill_1
XFILLER_15_256 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_763 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_752 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_741 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_395 vpwr vgnd scs8hd_fill_2
XPHY_730 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_796 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_785 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_774 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_440 vgnd vpwr scs8hd_decap_12
XANTENNA__292__A _277_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_92 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_495 vgnd vpwr scs8hd_decap_12
XFILLER_38_326 vpwr vgnd scs8hd_fill_2
XFILLER_65_134 vgnd vpwr scs8hd_fill_1
XFILLER_38_348 vpwr vgnd scs8hd_fill_2
XANTENNA__467__A _456_/A vgnd vpwr scs8hd_diode_2
XFILLER_65_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_61_362 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _289_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_315 vpwr vgnd scs8hd_fill_2
XFILLER_56_123 vgnd vpwr scs8hd_decap_4
XANTENNA__377__A _404_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_370 vpwr vgnd scs8hd_fill_2
XFILLER_71_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_259 vgnd vpwr scs8hd_decap_4
XFILLER_60_46 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_410 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_101 vpwr vgnd scs8hd_fill_2
XFILLER_47_123 vpwr vgnd scs8hd_fill_2
XFILLER_75_476 vgnd vpwr scs8hd_decap_12
XANTENNA__287__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_62_137 vgnd vpwr scs8hd_fill_1
XFILLER_43_340 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_513 vgnd vpwr scs8hd_decap_3
XFILLER_43_395 vgnd vpwr scs8hd_decap_3
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_571 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_593 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_582 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_123 vgnd vpwr scs8hd_decap_8
XFILLER_66_498 vgnd vpwr scs8hd_decap_12
XFILLER_53_148 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_502 vgnd vpwr scs8hd_decap_12
XFILLER_61_181 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_428 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_55_24 vpwr vgnd scs8hd_fill_2
XFILLER_29_178 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_57 vpwr vgnd scs8hd_fill_2
XFILLER_72_457 vgnd vpwr scs8hd_fill_1
X_470_ _448_/A _462_/A _470_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_148 vgnd vpwr scs8hd_decap_4
XFILLER_13_513 vgnd vpwr scs8hd_decap_3
XFILLER_25_362 vpwr vgnd scs8hd_fill_2
XFILLER_52_181 vgnd vpwr scs8hd_decap_6
XFILLER_40_332 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__570__A _596_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_288 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_75_273 vgnd vpwr scs8hd_decap_12
XFILLER_75_262 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_126 vpwr vgnd scs8hd_fill_2
XFILLER_16_351 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _593_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_118 vgnd vpwr scs8hd_decap_4
XFILLER_16_373 vgnd vpwr scs8hd_decap_6
X_599_ _599_/A _578_/X _599_/X vgnd vpwr scs8hd_or2_4
XANTENNA__464__B _467_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__480__A _447_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_410 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_465 vpwr vgnd scs8hd_fill_2
XFILLER_39_476 vpwr vgnd scs8hd_fill_2
XFILLER_66_295 vgnd vpwr scs8hd_decap_8
XFILLER_54_413 vgnd vpwr scs8hd_decap_4
XFILLER_26_137 vgnd vpwr scs8hd_decap_3
XANTENNA__358__C _358_/C vgnd vpwr scs8hd_diode_2
XFILLER_81_232 vgnd vpwr scs8hd_decap_12
XFILLER_54_468 vgnd vpwr scs8hd_decap_12
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XFILLER_26_159 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__374__B _376_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_332 vpwr vgnd scs8hd_fill_2
XFILLER_22_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__390__A _328_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_269 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _601_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_49_218 vpwr vgnd scs8hd_fill_2
XANTENNA__549__B _548_/X vgnd vpwr scs8hd_diode_2
XFILLER_66_56 vgnd vpwr scs8hd_decap_12
XFILLER_57_273 vpwr vgnd scs8hd_fill_2
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
XFILLER_72_232 vgnd vpwr scs8hd_decap_8
X_522_ _522_/A _523_/B _522_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_148 vpwr vgnd scs8hd_fill_2
XFILLER_82_44 vgnd vpwr scs8hd_decap_12
X_453_ _442_/A _456_/B _453_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_438 vgnd vpwr scs8hd_decap_3
XANTENNA__565__A _591_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_321 vpwr vgnd scs8hd_fill_2
X_384_ _471_/C _409_/C vgnd vpwr scs8hd_buf_1
XFILLER_40_151 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_92 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__459__B _451_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_280 vgnd vpwr scs8hd_decap_12
XFILLER_63_298 vgnd vpwr scs8hd_decap_4
XFILLER_63_287 vpwr vgnd scs8hd_fill_2
XFILLER_51_416 vgnd vpwr scs8hd_decap_4
XFILLER_51_405 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XANTENNA__475__A _442_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_181 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__B _383_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_240 vpwr vgnd scs8hd_fill_2
XFILLER_54_221 vgnd vpwr scs8hd_fill_1
XFILLER_27_435 vgnd vpwr scs8hd_decap_4
XFILLER_27_446 vpwr vgnd scs8hd_fill_2
XFILLER_36_59 vgnd vpwr scs8hd_decap_4
XFILLER_14_107 vgnd vpwr scs8hd_decap_3
XANTENNA__385__A _385_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_427 vgnd vpwr scs8hd_decap_6
XFILLER_14_129 vpwr vgnd scs8hd_fill_2
XFILLER_42_438 vpwr vgnd scs8hd_fill_2
XFILLER_42_449 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_324 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_77_324 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _567_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_77_379 vgnd vpwr scs8hd_decap_12
XANTENNA__279__B _313_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _266_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_468 vgnd vpwr scs8hd_decap_12
XANTENNA__295__A _301_/A vgnd vpwr scs8hd_diode_2
XFILLER_45_287 vpwr vgnd scs8hd_fill_2
X_505_ _504_/X _505_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_449 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_45_298 vgnd vpwr scs8hd_decap_4
XFILLER_13_151 vpwr vgnd scs8hd_fill_2
X_436_ _447_/A _429_/A _436_/Y vgnd vpwr scs8hd_nor2_4
X_367_ _340_/X _367_/B _367_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_471 vpwr vgnd scs8hd_fill_2
XFILLER_41_482 vgnd vpwr scs8hd_decap_6
XFILLER_9_166 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_298_ _301_/A _596_/A _298_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_68_302 vgnd vpwr scs8hd_decap_6
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _653_/HI ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_265 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vpwr vgnd scs8hd_fill_2
XFILLER_24_449 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_313 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_346 vpwr vgnd scs8hd_fill_2
XFILLER_59_357 vpwr vgnd scs8hd_fill_2
XFILLER_70_511 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_63_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_438 vgnd vpwr scs8hd_decap_4
XFILLER_27_287 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_176 vpwr vgnd scs8hd_fill_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_SLEEPB _393_/Y vgnd vpwr scs8hd_diode_2
XFILLER_77_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_338 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_18_254 vpwr vgnd scs8hd_fill_2
XFILLER_18_265 vgnd vpwr scs8hd_decap_3
XFILLER_73_393 vgnd vpwr scs8hd_fill_1
XFILLER_18_298 vgnd vpwr scs8hd_fill_1
X_419_ _522_/A _456_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _609_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_143 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_8
XFILLER_64_382 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_213 vgnd vpwr scs8hd_fill_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_49 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_474 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _541_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_143 vgnd vpwr scs8hd_decap_4
XFILLER_58_79 vpwr vgnd scs8hd_fill_2
XFILLER_58_68 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_327 vgnd vpwr scs8hd_decap_6
XFILLER_74_56 vgnd vpwr scs8hd_decap_12
XFILLER_62_308 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__557__B _561_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XPHY_720 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_753 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_742 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_374 vpwr vgnd scs8hd_fill_2
XPHY_731 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_SLEEPB _354_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__573__A _599_/A vgnd vpwr scs8hd_diode_2
XPHY_786 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_775 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_764 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_797 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_452 vgnd vpwr scs8hd_decap_12
XANTENNA__292__B _594_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _568_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _650_/HI ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_65_146 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_105 vgnd vpwr scs8hd_decap_12
XANTENNA__467__B _467_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_319 vgnd vpwr scs8hd_decap_4
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_61_341 vpwr vgnd scs8hd_fill_2
XFILLER_61_385 vpwr vgnd scs8hd_fill_2
XANTENNA__483__A _482_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_SLEEPB _489_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_327 vpwr vgnd scs8hd_fill_2
XFILLER_56_146 vgnd vpwr scs8hd_fill_1
XFILLER_29_338 vpwr vgnd scs8hd_fill_2
XANTENNA__377__B _376_/B vgnd vpwr scs8hd_diode_2
XFILLER_44_308 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XFILLER_52_352 vpwr vgnd scs8hd_fill_2
XANTENNA__393__A _404_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_503 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q
+ _507_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_260 vpwr vgnd scs8hd_fill_2
XFILLER_60_69 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_459 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q
+ _464_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_75_422 vgnd vpwr scs8hd_decap_4
XANTENNA__568__A _594_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_146 vgnd vpwr scs8hd_decap_3
XFILLER_18_60 vgnd vpwr scs8hd_fill_1
XANTENNA__287__B _327_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_168 vgnd vpwr scs8hd_fill_1
XFILLER_47_179 vpwr vgnd scs8hd_fill_2
XFILLER_43_374 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q
+ _416_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_81 vgnd vpwr scs8hd_decap_8
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_594 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_583 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_572 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_91 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q
+ _364_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_66_444 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__478__A _456_/A vgnd vpwr scs8hd_diode_2
XFILLER_81_403 vgnd vpwr scs8hd_decap_12
XFILLER_26_308 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_SLEEPB _456_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_382 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_341 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_514 vpwr vgnd scs8hd_fill_2
XFILLER_34_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_28 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_69_260 vpwr vgnd scs8hd_fill_2
XFILLER_57_400 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_102 vpwr vgnd scs8hd_fill_2
XFILLER_69_293 vpwr vgnd scs8hd_fill_2
XANTENNA__388__A _314_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_477 vgnd vpwr scs8hd_decap_8
XFILLER_44_127 vpwr vgnd scs8hd_fill_2
XANTENNA__570__B _562_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _647_/HI ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_50 vgnd vpwr scs8hd_decap_8
XFILLER_20_72 vgnd vpwr scs8hd_decap_8
XFILLER_20_83 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_219 vpwr vgnd scs8hd_fill_2
XFILLER_67_208 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_70 vgnd vpwr scs8hd_decap_4
XANTENNA__298__A _301_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_433 vpwr vgnd scs8hd_fill_2
XFILLER_75_241 vgnd vpwr scs8hd_decap_3
XFILLER_75_296 vgnd vpwr scs8hd_decap_8
XFILLER_63_458 vgnd vpwr scs8hd_fill_1
X_598_ _304_/B _581_/A _598_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q
+ _323_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_43_193 vpwr vgnd scs8hd_fill_2
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__480__B _481_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_SLEEPB _420_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_400 vgnd vpwr scs8hd_fill_1
XFILLER_66_285 vgnd vpwr scs8hd_decap_8
XFILLER_54_436 vgnd vpwr scs8hd_decap_3
XFILLER_26_127 vpwr vgnd scs8hd_fill_2
XANTENNA__358__D _409_/D vgnd vpwr scs8hd_diode_2
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_41_108 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _273_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_27 vpwr vgnd scs8hd_fill_2
XFILLER_41_49 vgnd vpwr scs8hd_fill_1
XANTENNA__390__B _387_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_68 vpwr vgnd scs8hd_fill_2
XFILLER_17_105 vgnd vpwr scs8hd_fill_1
XFILLER_45_425 vpwr vgnd scs8hd_fill_2
X_521_ _510_/A _523_/B _521_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_45_469 vgnd vpwr scs8hd_decap_12
XFILLER_82_56 vgnd vpwr scs8hd_decap_6
X_452_ _441_/A _456_/B _452_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__565__B _568_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
X_383_ address[8] _383_/B _471_/C vgnd vpwr scs8hd_nand2_4
XFILLER_13_344 vgnd vpwr scs8hd_fill_1
XANTENNA__581__A _581_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_388 vgnd vpwr scs8hd_decap_8
XFILLER_40_174 vpwr vgnd scs8hd_fill_2
XFILLER_40_185 vgnd vpwr scs8hd_decap_8
XFILLER_40_196 vgnd vpwr scs8hd_decap_4
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_292 vgnd vpwr scs8hd_decap_12
XFILLER_48_241 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_285 vpwr vgnd scs8hd_fill_2
XFILLER_51_428 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_SLEEPB _376_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__475__B _476_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_193 vgnd vpwr scs8hd_fill_1
XFILLER_44_480 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__491__A _423_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__C _358_/C vgnd vpwr scs8hd_diode_2
XFILLER_27_414 vpwr vgnd scs8hd_fill_2
XFILLER_39_263 vpwr vgnd scs8hd_fill_2
XFILLER_39_274 vpwr vgnd scs8hd_fill_2
XFILLER_54_233 vgnd vpwr scs8hd_fill_1
XFILLER_54_266 vgnd vpwr scs8hd_decap_8
XANTENNA__385__B _382_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_406 vgnd vpwr scs8hd_fill_1
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_SLEEPB _510_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_447 vgnd vpwr scs8hd_decap_8
XANTENNA__576__A _270_/B vgnd vpwr scs8hd_diode_2
XFILLER_45_233 vgnd vpwr scs8hd_decap_8
XFILLER_60_203 vgnd vpwr scs8hd_decap_8
X_504_ _409_/A _382_/A _515_/C _482_/D _504_/X vgnd vpwr scs8hd_or4_4
XFILLER_33_428 vpwr vgnd scs8hd_fill_2
XANTENNA__295__B _294_/X vgnd vpwr scs8hd_diode_2
XFILLER_60_247 vgnd vpwr scs8hd_decap_3
XFILLER_26_82 vgnd vpwr scs8hd_decap_6
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_26_491 vgnd vpwr scs8hd_decap_12
XFILLER_13_130 vpwr vgnd scs8hd_fill_2
XFILLER_41_450 vgnd vpwr scs8hd_fill_1
X_435_ _457_/A _429_/X _435_/Y vgnd vpwr scs8hd_nor2_4
X_366_ _404_/A _360_/X _366_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_41_461 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_297_ _297_/A _596_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ _525_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_233 vgnd vpwr scs8hd_decap_4
XANTENNA__486__A _413_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_51_236 vpwr vgnd scs8hd_fill_2
XFILLER_51_225 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_8
XFILLER_74_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_SLEEPB _477_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_233 vpwr vgnd scs8hd_fill_2
XANTENNA__396__A _385_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_247 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y _632_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_133 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_2_398 vgnd vpwr scs8hd_decap_12
XFILLER_65_306 vpwr vgnd scs8hd_fill_2
XFILLER_73_361 vgnd vpwr scs8hd_decap_3
XFILLER_61_501 vgnd vpwr scs8hd_decap_12
XFILLER_37_92 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_418_ _466_/A _422_/B _418_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_483 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_280 vgnd vpwr scs8hd_decap_4
X_349_ _314_/X _348_/X _349_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ _500_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ _457_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_247 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ _405_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_486 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _532_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_166 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ _356_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_306 vpwr vgnd scs8hd_fill_2
XFILLER_74_68 vgnd vpwr scs8hd_decap_12
XFILLER_43_501 vgnd vpwr scs8hd_decap_12
XFILLER_82_180 vgnd vpwr scs8hd_decap_6
XPHY_710 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_236 vgnd vpwr scs8hd_decap_4
XPHY_754 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_743 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_732 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_721 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__573__B _552_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_206 vgnd vpwr scs8hd_decap_8
XPHY_787 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_776 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_765 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_291 vgnd vpwr scs8hd_decap_4
XFILLER_30_239 vpwr vgnd scs8hd_fill_2
XPHY_798 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_464 vgnd vpwr scs8hd_decap_12
XFILLER_65_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_80_117 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_69_420 vpwr vgnd scs8hd_fill_2
XFILLER_69_453 vpwr vgnd scs8hd_fill_2
XFILLER_69_486 vpwr vgnd scs8hd_fill_2
XFILLER_25_501 vgnd vpwr scs8hd_decap_12
XFILLER_64_180 vpwr vgnd scs8hd_fill_2
XFILLER_44_27 vpwr vgnd scs8hd_fill_2
XFILLER_52_386 vgnd vpwr scs8hd_decap_8
XANTENNA__393__B _387_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_515 vgnd vpwr scs8hd_fill_1
XFILLER_12_228 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_272 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__568__B _568_/B vgnd vpwr scs8hd_diode_2
XFILLER_47_114 vpwr vgnd scs8hd_fill_2
XFILLER_75_489 vgnd vpwr scs8hd_decap_12
XFILLER_18_50 vgnd vpwr scs8hd_fill_1
XFILLER_62_106 vgnd vpwr scs8hd_decap_8
XFILLER_18_72 vgnd vpwr scs8hd_decap_8
XANTENNA__584__A _584_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_353 vpwr vgnd scs8hd_fill_2
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_595 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_584 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_573 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_81 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_90 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XANTENNA__478__B _476_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_158 vpwr vgnd scs8hd_fill_2
XFILLER_81_415 vgnd vpwr scs8hd_decap_12
XANTENNA__494__A _494_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_180 vgnd vpwr scs8hd_decap_4
XFILLER_61_161 vpwr vgnd scs8hd_fill_2
XFILLER_61_194 vpwr vgnd scs8hd_fill_2
XFILLER_61_172 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_16 vpwr vgnd scs8hd_fill_2
XFILLER_39_38 vpwr vgnd scs8hd_fill_2
XFILLER_57_445 vpwr vgnd scs8hd_fill_2
XFILLER_57_423 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XANTENNA__388__B _387_/X vgnd vpwr scs8hd_diode_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_6
XFILLER_72_415 vgnd vpwr scs8hd_decap_8
XFILLER_57_489 vgnd vpwr scs8hd_decap_12
XFILLER_72_459 vgnd vpwr scs8hd_decap_12
XFILLER_25_342 vgnd vpwr scs8hd_decap_4
XFILLER_25_397 vgnd vpwr scs8hd_decap_4
XFILLER_40_312 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XANTENNA__579__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_75_220 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__298__B _596_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _652_/HI ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_437 vpwr vgnd scs8hd_fill_2
XFILLER_63_415 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_320 vpwr vgnd scs8hd_fill_2
XFILLER_28_180 vgnd vpwr scs8hd_decap_4
XFILLER_28_191 vgnd vpwr scs8hd_decap_6
XFILLER_71_470 vgnd vpwr scs8hd_decap_12
X_597_ _597_/A _581_/A _597_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_92 vgnd vpwr scs8hd_fill_1
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_367 vpwr vgnd scs8hd_fill_2
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_91 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__489__A _522_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_106 vgnd vpwr scs8hd_decap_8
XFILLER_39_489 vgnd vpwr scs8hd_decap_12
XFILLER_81_245 vgnd vpwr scs8hd_decap_12
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_161 vpwr vgnd scs8hd_fill_2
XFILLER_34_183 vpwr vgnd scs8hd_fill_2
XFILLER_10_507 vgnd vpwr scs8hd_decap_8
XFILLER_22_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__399__A _314_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_286 vpwr vgnd scs8hd_fill_2
X_520_ _509_/A _523_/B _520_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_117 vgnd vpwr scs8hd_decap_3
XFILLER_45_404 vpwr vgnd scs8hd_fill_2
XFILLER_45_415 vgnd vpwr scs8hd_decap_4
XFILLER_57_297 vpwr vgnd scs8hd_fill_2
XFILLER_45_437 vpwr vgnd scs8hd_fill_2
X_451_ _451_/A _456_/B vgnd vpwr scs8hd_buf_1
XFILLER_32_109 vgnd vpwr scs8hd_decap_8
XFILLER_53_481 vgnd vpwr scs8hd_decap_6
X_382_ _382_/A _382_/X vgnd vpwr scs8hd_buf_1
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_367 vgnd vpwr scs8hd_decap_4
XFILLER_13_356 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y _604_/A vgnd vpwr scs8hd_buf_1
XFILLER_31_50 vgnd vpwr scs8hd_decap_4
XFILLER_48_253 vgnd vpwr scs8hd_decap_4
XFILLER_63_212 vgnd vpwr scs8hd_decap_4
XFILLER_36_426 vpwr vgnd scs8hd_fill_2
XFILLER_63_234 vgnd vpwr scs8hd_decap_4
XFILLER_63_223 vpwr vgnd scs8hd_fill_2
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_256 vgnd vpwr scs8hd_decap_3
X_649_ _649_/HI _649_/LO vgnd vpwr scs8hd_conb_1
XFILLER_44_492 vgnd vpwr scs8hd_decap_12
XFILLER_82_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_153 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_197 vpwr vgnd scs8hd_fill_2
XANTENNA__491__B _491_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__D _471_/D vgnd vpwr scs8hd_diode_2
XFILLER_27_426 vgnd vpwr scs8hd_fill_1
XFILLER_54_245 vpwr vgnd scs8hd_fill_2
XFILLER_27_459 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__385__C _409_/C vgnd vpwr scs8hd_diode_2
XFILLER_54_289 vgnd vpwr scs8hd_decap_4
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_50_451 vgnd vpwr scs8hd_decap_6
XFILLER_50_440 vgnd vpwr scs8hd_decap_4
XFILLER_10_304 vpwr vgnd scs8hd_fill_2
XFILLER_10_337 vgnd vpwr scs8hd_decap_12
XFILLER_22_186 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _586_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _649_/HI ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_1_0_clk/X ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XANTENNA__576__B _574_/X vgnd vpwr scs8hd_diode_2
X_503_ _425_/A _495_/A _503_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_256 vgnd vpwr scs8hd_decap_12
XFILLER_60_237 vgnd vpwr scs8hd_decap_8
XFILLER_60_226 vpwr vgnd scs8hd_fill_2
X_434_ _456_/A _429_/X _434_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_259 vgnd vpwr scs8hd_decap_12
XANTENNA__592__A _592_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_164 vgnd vpwr scs8hd_decap_4
X_365_ _392_/A _360_/X _365_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_197 vgnd vpwr scs8hd_decap_3
XFILLER_9_157 vgnd vpwr scs8hd_decap_3
X_296_ _282_/C _241_/B address[3] _259_/A _297_/A vgnd vpwr scs8hd_or4_4
XFILLER_42_60 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_330 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_348 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_76_370 vgnd vpwr scs8hd_decap_12
XFILLER_64_510 vgnd vpwr scs8hd_decap_6
XFILLER_36_201 vgnd vpwr scs8hd_decap_4
XANTENNA__486__B _490_/B vgnd vpwr scs8hd_diode_2
XFILLER_51_204 vgnd vpwr scs8hd_decap_4
XFILLER_36_289 vpwr vgnd scs8hd_fill_2
XFILLER_51_259 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _546_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_326 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_49 vpwr vgnd scs8hd_fill_2
XFILLER_27_223 vpwr vgnd scs8hd_fill_2
XANTENNA__396__B _382_/X vgnd vpwr scs8hd_diode_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_245 vpwr vgnd scs8hd_fill_2
XFILLER_27_267 vgnd vpwr scs8hd_decap_4
XFILLER_82_373 vgnd vpwr scs8hd_decap_12
XFILLER_42_226 vpwr vgnd scs8hd_fill_2
XFILLER_23_473 vpwr vgnd scs8hd_fill_2
XFILLER_23_484 vgnd vpwr scs8hd_decap_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_8
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_2_300 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_123 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__587__A _587_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_510 vgnd vpwr scs8hd_decap_6
XFILLER_61_513 vgnd vpwr scs8hd_decap_3
XFILLER_33_237 vgnd vpwr scs8hd_fill_1
X_417_ _510_/A _466_/A vgnd vpwr scs8hd_buf_1
XFILLER_53_92 vpwr vgnd scs8hd_fill_2
XFILLER_14_495 vgnd vpwr scs8hd_decap_12
X_348_ _356_/B _348_/X vgnd vpwr scs8hd_buf_1
X_279_ _278_/X _313_/A _280_/A vgnd vpwr scs8hd_or2_4
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_123 vgnd vpwr scs8hd_decap_12
XANTENNA__497__A _413_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_8
XFILLER_24_226 vgnd vpwr scs8hd_decap_6
XFILLER_32_281 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_498 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _646_/HI ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_123 vgnd vpwr scs8hd_decap_3
XFILLER_55_340 vpwr vgnd scs8hd_fill_2
XFILLER_70_310 vpwr vgnd scs8hd_fill_2
XFILLER_55_373 vpwr vgnd scs8hd_fill_2
XFILLER_55_362 vpwr vgnd scs8hd_fill_2
XFILLER_15_215 vgnd vpwr scs8hd_fill_1
XFILLER_43_513 vgnd vpwr scs8hd_decap_3
XPHY_711 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_700 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_248 vpwr vgnd scs8hd_fill_2
XPHY_744 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_387 vgnd vpwr scs8hd_decap_8
XPHY_733 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_722 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_218 vpwr vgnd scs8hd_fill_2
XPHY_777 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_766 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_755 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_398 vgnd vpwr scs8hd_decap_4
XFILLER_23_270 vpwr vgnd scs8hd_fill_2
XPHY_799 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_788 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_403 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_476 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_78_410 vgnd vpwr scs8hd_decap_12
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_38_318 vgnd vpwr scs8hd_fill_1
XFILLER_65_126 vpwr vgnd scs8hd_fill_2
XFILLER_48_81 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_80_129 vgnd vpwr scs8hd_decap_12
XFILLER_46_384 vpwr vgnd scs8hd_fill_2
XFILLER_61_321 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_207 vpwr vgnd scs8hd_fill_2
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XFILLER_14_270 vgnd vpwr scs8hd_decap_4
XFILLER_21_229 vpwr vgnd scs8hd_fill_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_69_432 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_104 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _610_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_351 vpwr vgnd scs8hd_fill_2
XFILLER_25_513 vgnd vpwr scs8hd_decap_3
XFILLER_37_362 vpwr vgnd scs8hd_fill_2
XFILLER_52_365 vpwr vgnd scs8hd_fill_2
XFILLER_12_207 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_129 vgnd vpwr scs8hd_decap_6
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XANTENNA__584__B _587_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_365 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _593_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_50 vgnd vpwr scs8hd_fill_1
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XPHY_596 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_585 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_574 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_284 vgnd vpwr scs8hd_decap_12
XFILLER_50_60 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_93 vgnd vpwr scs8hd_fill_1
XFILLER_78_251 vgnd vpwr scs8hd_decap_12
XFILLER_66_413 vpwr vgnd scs8hd_fill_2
XFILLER_38_115 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_332 vgnd vpwr scs8hd_decap_4
XFILLER_46_192 vgnd vpwr scs8hd_decap_4
XFILLER_34_365 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_184 vgnd vpwr scs8hd_decap_3
XFILLER_34_398 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _643_/HI ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_273 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_118 vpwr vgnd scs8hd_fill_2
XFILLER_72_449 vgnd vpwr scs8hd_decap_8
XFILLER_80_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _624_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_376 vpwr vgnd scs8hd_fill_2
XFILLER_71_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_96 vgnd vpwr scs8hd_decap_4
XANTENNA__579__B _578_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_497 vgnd vpwr scs8hd_decap_12
XFILLER_75_254 vpwr vgnd scs8hd_fill_2
XFILLER_63_405 vgnd vpwr scs8hd_fill_1
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XANTENNA__595__A _294_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_596_ _596_/A _581_/A _596_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_365 vgnd vpwr scs8hd_decap_6
XFILLER_71_482 vgnd vpwr scs8hd_decap_6
XFILLER_31_302 vgnd vpwr scs8hd_fill_1
XFILLER_43_162 vgnd vpwr scs8hd_decap_8
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_346 vpwr vgnd scs8hd_fill_2
XFILLER_31_357 vpwr vgnd scs8hd_fill_2
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__489__B _490_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_424 vgnd vpwr scs8hd_fill_1
XFILLER_39_446 vgnd vpwr scs8hd_decap_4
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_81_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _632_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_313 vgnd vpwr scs8hd_decap_12
XFILLER_34_173 vgnd vpwr scs8hd_fill_1
XFILLER_22_346 vgnd vpwr scs8hd_decap_12
XFILLER_22_379 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_390 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_SLEEPB _332_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__399__B _404_/B vgnd vpwr scs8hd_diode_2
XFILLER_66_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_254 vpwr vgnd scs8hd_fill_2
XFILLER_72_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_72_268 vgnd vpwr scs8hd_decap_4
X_450_ _450_/A _451_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_60_408 vgnd vpwr scs8hd_fill_1
XFILLER_25_184 vgnd vpwr scs8hd_decap_3
X_381_ _471_/B _382_/A vgnd vpwr scs8hd_inv_8
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_306 vgnd vpwr scs8hd_decap_12
XFILLER_40_132 vpwr vgnd scs8hd_fill_2
XFILLER_40_143 vpwr vgnd scs8hd_fill_2
XFILLER_15_96 vpwr vgnd scs8hd_fill_2
XFILLER_40_165 vgnd vpwr scs8hd_decap_6
XFILLER_5_501 vgnd vpwr scs8hd_decap_12
XFILLER_31_95 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_449 vgnd vpwr scs8hd_decap_6
XFILLER_48_298 vgnd vpwr scs8hd_decap_8
X_648_ _648_/HI _648_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_80 vgnd vpwr scs8hd_decap_12
X_579_ address[4] _578_/X _579_/X vgnd vpwr scs8hd_or2_4
XFILLER_31_132 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_176 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _556_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_3 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_361 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_39_221 vpwr vgnd scs8hd_fill_2
XFILLER_39_287 vgnd vpwr scs8hd_decap_4
XFILLER_39_298 vgnd vpwr scs8hd_decap_6
XANTENNA__385__D _409_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_110 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_349 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_419 vpwr vgnd scs8hd_fill_2
X_502_ _423_/A _495_/A _502_/Y vgnd vpwr scs8hd_nor2_4
X_433_ _466_/A _429_/X _433_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__592__B _594_/B vgnd vpwr scs8hd_diode_2
X_364_ _391_/A _360_/X _364_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_187 vpwr vgnd scs8hd_fill_2
X_295_ _301_/A _294_/X _295_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_SLEEPB _443_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_342 vgnd vpwr scs8hd_decap_12
XFILLER_68_316 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_382 vgnd vpwr scs8hd_decap_12
XFILLER_36_224 vgnd vpwr scs8hd_decap_3
XFILLER_32_430 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_191 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_39 vgnd vpwr scs8hd_decap_4
XFILLER_27_202 vpwr vgnd scs8hd_fill_2
XANTENNA__396__C _409_/C vgnd vpwr scs8hd_diode_2
XFILLER_82_385 vgnd vpwr scs8hd_decap_12
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_15_419 vpwr vgnd scs8hd_fill_2
XFILLER_23_441 vgnd vpwr scs8hd_decap_4
XFILLER_23_452 vpwr vgnd scs8hd_fill_2
XFILLER_50_293 vgnd vpwr scs8hd_fill_1
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_2_312 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_135 vgnd vpwr scs8hd_decap_12
XANTENNA__587__B _587_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_202 vgnd vpwr scs8hd_fill_1
XFILLER_18_224 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_330 vgnd vpwr scs8hd_decap_4
XFILLER_18_246 vpwr vgnd scs8hd_fill_2
XFILLER_73_385 vgnd vpwr scs8hd_decap_8
XFILLER_73_374 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_SLEEPB _401_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_227 vpwr vgnd scs8hd_fill_2
XFILLER_26_290 vgnd vpwr scs8hd_decap_4
X_416_ _454_/A _422_/B _416_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_71 vpwr vgnd scs8hd_fill_2
X_347_ _346_/X _356_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_278_ address[3] _278_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_113 vgnd vpwr scs8hd_fill_1
XFILLER_38_3 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_135 vgnd vpwr scs8hd_decap_4
XFILLER_68_157 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__497__B _499_/B vgnd vpwr scs8hd_diode_2
XFILLER_49_360 vpwr vgnd scs8hd_fill_2
XFILLER_49_382 vgnd vpwr scs8hd_decap_3
XFILLER_76_190 vgnd vpwr scs8hd_decap_12
XFILLER_24_205 vgnd vpwr scs8hd_decap_8
XFILLER_64_396 vgnd vpwr scs8hd_fill_1
XFILLER_20_433 vgnd vpwr scs8hd_decap_4
XFILLER_32_271 vpwr vgnd scs8hd_fill_2
XFILLER_20_455 vgnd vpwr scs8hd_decap_3
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_74_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _304_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_74_15 vgnd vpwr scs8hd_decap_12
XFILLER_70_333 vgnd vpwr scs8hd_fill_1
XPHY_701 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_745 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_734 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_723 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_712 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_778 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_767 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_756 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_411 vgnd vpwr scs8hd_decap_12
XPHY_789 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_415 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_96 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_SLEEPB _363_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_422 vgnd vpwr scs8hd_decap_12
XANTENNA__598__A _304_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_308 vgnd vpwr scs8hd_decap_3
XFILLER_58_190 vgnd vpwr scs8hd_decap_4
XFILLER_73_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_34_503 vgnd vpwr scs8hd_decap_12
XFILLER_46_363 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_396 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_80_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y _609_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_466 vgnd vpwr scs8hd_decap_12
XFILLER_29_319 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__301__A _301_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_127 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_SLEEPB _497_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_149 vgnd vpwr scs8hd_decap_4
XFILLER_52_311 vpwr vgnd scs8hd_fill_2
XFILLER_37_374 vpwr vgnd scs8hd_fill_2
XFILLER_37_385 vpwr vgnd scs8hd_fill_2
XFILLER_52_322 vpwr vgnd scs8hd_fill_2
XFILLER_37_396 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_208 vgnd vpwr scs8hd_decap_12
XFILLER_69_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_138 vpwr vgnd scs8hd_fill_2
XFILLER_55_193 vgnd vpwr scs8hd_decap_3
XFILLER_55_171 vpwr vgnd scs8hd_fill_2
XFILLER_70_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_62 vgnd vpwr scs8hd_fill_1
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_586 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_575 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_597 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_440 vgnd vpwr scs8hd_decap_12
XFILLER_78_263 vgnd vpwr scs8hd_decap_12
XFILLER_66_436 vgnd vpwr scs8hd_decap_3
XFILLER_81_428 vgnd vpwr scs8hd_decap_12
XFILLER_34_300 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _251_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_388 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_SLEEPB _464_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _598_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q
+ _519_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_29 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _648_/HI ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_69_252 vpwr vgnd scs8hd_fill_2
XFILLER_69_241 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q
+ _476_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_28 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y _627_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_193 vpwr vgnd scs8hd_fill_2
XFILLER_52_141 vgnd vpwr scs8hd_decap_12
XFILLER_80_483 vgnd vpwr scs8hd_decap_12
XFILLER_71_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_303 vgnd vpwr scs8hd_decap_3
XFILLER_40_347 vpwr vgnd scs8hd_fill_2
XFILLER_40_358 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q
+ _433_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _538_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ _376_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__595__B _581_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_595_ _294_/X _581_/A _595_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_50 vpwr vgnd scs8hd_fill_2
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_71 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_281 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_66_244 vpwr vgnd scs8hd_fill_2
XFILLER_39_469 vgnd vpwr scs8hd_decap_4
XFILLER_66_266 vgnd vpwr scs8hd_decap_6
XFILLER_54_428 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_SLEEPB _431_/Y vgnd vpwr scs8hd_diode_2
XFILLER_81_269 vgnd vpwr scs8hd_decap_12
XFILLER_34_152 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q
+ _399_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_491 vgnd vpwr scs8hd_decap_12
XFILLER_45_428 vpwr vgnd scs8hd_fill_2
XFILLER_82_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_450 vpwr vgnd scs8hd_fill_2
XFILLER_53_461 vpwr vgnd scs8hd_fill_2
X_380_ _380_/A _385_/A vgnd vpwr scs8hd_buf_1
XFILLER_13_336 vgnd vpwr scs8hd_decap_8
XFILLER_15_86 vgnd vpwr scs8hd_fill_1
XFILLER_9_318 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q
+ _350_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_513 vgnd vpwr scs8hd_decap_3
XFILLER_0_273 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_56_60 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
X_647_ _647_/HI _647_/LO vgnd vpwr scs8hd_conb_1
XFILLER_51_409 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XFILLER_44_450 vgnd vpwr scs8hd_decap_8
X_578_ address[6] address[7] _578_/C _482_/D _578_/X vgnd vpwr scs8hd_or4_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _572_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _530_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_166 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_373 vgnd vpwr scs8hd_decap_12
XFILLER_68_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _645_/HI ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
.ends

