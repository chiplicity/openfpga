magic
tech EFS8A
magscale 1 2
timestamp 1603297593
<< locali >>
rect 18889 19873 19050 19907
rect 18889 19839 18923 19873
rect 16071 18785 16106 18819
rect 15531 17289 15669 17323
rect 21193 16677 21268 16711
rect 23575 15657 23581 15691
rect 23575 15589 23609 15657
rect 9631 15521 9758 15555
rect 12575 15521 12702 15555
rect 24035 14807 24069 14875
rect 24035 14773 24041 14807
rect 11431 14569 11437 14603
rect 11431 14501 11465 14569
rect 24133 13821 24294 13855
rect 24133 13719 24167 13821
rect 14749 12631 14783 12937
rect 17359 12325 17404 12359
rect 18981 10999 19015 11169
rect 15577 10523 15611 10693
rect 7055 10081 7090 10115
rect 6009 9503 6043 9673
rect 14933 9503 14967 9605
rect 15663 9129 15669 9163
rect 15663 9061 15697 9129
rect 15945 8415 15979 8585
rect 8211 6953 8217 6987
rect 12351 6953 12357 6987
rect 15663 6953 15669 6987
rect 23575 6953 23581 6987
rect 8211 6885 8245 6953
rect 12351 6885 12385 6953
rect 15663 6885 15697 6953
rect 23575 6885 23609 6953
rect 8861 6851 8895 6885
rect 5181 6817 5342 6851
rect 8769 6817 8895 6851
rect 24995 6817 25030 6851
rect 5181 6783 5215 6817
rect 7791 6749 7879 6783
rect 1443 5729 1478 5763
rect 6043 5729 6078 5763
rect 15663 4777 15669 4811
rect 15663 4709 15697 4777
rect 5491 4641 5526 4675
rect 3847 4233 3985 4267
rect 9976 3621 10044 3655
rect 2915 3553 3042 3587
rect 17877 2839 17911 2941
rect 3111 2533 3249 2567
rect 4951 2533 5089 2567
rect 23029 2295 23063 2601
<< viali >>
rect 24501 24905 24535 24939
rect 24317 24701 24351 24735
rect 24869 24701 24903 24735
rect 19901 24361 19935 24395
rect 24777 24361 24811 24395
rect 7424 24225 7458 24259
rect 18372 24225 18406 24259
rect 19717 24225 19751 24259
rect 23121 24225 23155 24259
rect 24593 24225 24627 24259
rect 23305 24089 23339 24123
rect 7527 24021 7561 24055
rect 18475 24021 18509 24055
rect 2881 23817 2915 23851
rect 3893 23817 3927 23851
rect 8125 23817 8159 23851
rect 18429 23817 18463 23851
rect 20085 23817 20119 23851
rect 22661 23817 22695 23851
rect 24777 23817 24811 23851
rect 25145 23817 25179 23851
rect 11437 23749 11471 23783
rect 17049 23749 17083 23783
rect 19165 23749 19199 23783
rect 21189 23749 21223 23783
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 2488 23613 2522 23647
rect 3484 23613 3518 23647
rect 7332 23613 7366 23647
rect 7757 23613 7791 23647
rect 8344 23613 8378 23647
rect 8769 23613 8803 23647
rect 11028 23613 11062 23647
rect 12484 23613 12518 23647
rect 12909 23613 12943 23647
rect 16865 23613 16899 23647
rect 18245 23613 18279 23647
rect 18797 23613 18831 23647
rect 19901 23613 19935 23647
rect 21005 23613 21039 23647
rect 21557 23613 21591 23647
rect 22477 23613 22511 23647
rect 1547 23545 1581 23579
rect 3571 23545 3605 23579
rect 8447 23545 8481 23579
rect 11115 23545 11149 23579
rect 17417 23545 17451 23579
rect 20453 23545 20487 23579
rect 23029 23545 23063 23579
rect 2559 23477 2593 23511
rect 7435 23477 7469 23511
rect 12587 23477 12621 23511
rect 19809 23477 19843 23511
rect 23397 23477 23431 23511
rect 24777 23273 24811 23307
rect 24593 23137 24627 23171
rect 25145 22729 25179 22763
rect 24660 22525 24694 22559
rect 24731 22389 24765 22423
rect 25513 22389 25547 22423
rect 24777 21641 24811 21675
rect 24593 21437 24627 21471
rect 25237 21301 25271 21335
rect 20948 20961 20982 20995
rect 21051 20757 21085 20791
rect 24777 20553 24811 20587
rect 19441 20349 19475 20383
rect 19901 20349 19935 20383
rect 24593 20349 24627 20383
rect 25145 20349 25179 20383
rect 19625 20213 19659 20247
rect 20453 20213 20487 20247
rect 20913 20213 20947 20247
rect 19993 20009 20027 20043
rect 23719 20009 23753 20043
rect 16072 19873 16106 19907
rect 21005 19873 21039 19907
rect 22512 19873 22546 19907
rect 23648 19873 23682 19907
rect 18889 19805 18923 19839
rect 16175 19669 16209 19703
rect 19119 19669 19153 19703
rect 21189 19669 21223 19703
rect 22615 19669 22649 19703
rect 16957 19465 16991 19499
rect 19349 19465 19383 19499
rect 22569 19465 22603 19499
rect 24777 19465 24811 19499
rect 16681 19397 16715 19431
rect 20085 19329 20119 19363
rect 21005 19329 21039 19363
rect 16196 19261 16230 19295
rect 18429 19261 18463 19295
rect 21465 19261 21499 19295
rect 21649 19261 21683 19295
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 20177 19193 20211 19227
rect 20729 19193 20763 19227
rect 21557 19193 21591 19227
rect 16267 19125 16301 19159
rect 18613 19125 18647 19159
rect 19901 19125 19935 19159
rect 23857 19125 23891 19159
rect 19165 18921 19199 18955
rect 17141 18853 17175 18887
rect 17233 18853 17267 18887
rect 19349 18853 19383 18887
rect 19441 18853 19475 18887
rect 21005 18853 21039 18887
rect 21097 18853 21131 18887
rect 16037 18785 16071 18819
rect 23248 18785 23282 18819
rect 24292 18785 24326 18819
rect 17417 18717 17451 18751
rect 19993 18717 20027 18751
rect 21465 18717 21499 18751
rect 21925 18717 21959 18751
rect 16175 18581 16209 18615
rect 18429 18581 18463 18615
rect 23351 18581 23385 18615
rect 24363 18581 24397 18615
rect 21189 18377 21223 18411
rect 21557 18377 21591 18411
rect 25421 18377 25455 18411
rect 16129 18241 16163 18275
rect 18153 18241 18187 18275
rect 18521 18241 18555 18275
rect 20177 18241 20211 18275
rect 20821 18241 20855 18275
rect 21741 18241 21775 18275
rect 22201 18241 22235 18275
rect 23029 18241 23063 18275
rect 12484 18173 12518 18207
rect 12909 18173 12943 18207
rect 14448 18173 14482 18207
rect 14841 18173 14875 18207
rect 15428 18173 15462 18207
rect 17049 18173 17083 18207
rect 23857 18173 23891 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 12587 18105 12621 18139
rect 15209 18105 15243 18139
rect 17141 18105 17175 18139
rect 18245 18105 18279 18139
rect 19349 18105 19383 18139
rect 19993 18105 20027 18139
rect 20269 18105 20303 18139
rect 21833 18105 21867 18139
rect 24409 18105 24443 18139
rect 14519 18037 14553 18071
rect 15531 18037 15565 18071
rect 17417 18037 17451 18071
rect 17877 18037 17911 18071
rect 23489 18037 23523 18071
rect 24685 18037 24719 18071
rect 17877 17833 17911 17867
rect 18245 17833 18279 17867
rect 20177 17833 20211 17867
rect 21097 17833 21131 17867
rect 24133 17833 24167 17867
rect 24777 17833 24811 17867
rect 13093 17765 13127 17799
rect 13185 17765 13219 17799
rect 17049 17765 17083 17799
rect 18613 17765 18647 17799
rect 21649 17765 21683 17799
rect 22201 17765 22235 17799
rect 23213 17765 23247 17799
rect 19165 17697 19199 17731
rect 24593 17697 24627 17731
rect 15853 17629 15887 17663
rect 16957 17629 16991 17663
rect 17601 17629 17635 17663
rect 18521 17629 18555 17663
rect 19809 17629 19843 17663
rect 21557 17629 21591 17663
rect 23121 17629 23155 17663
rect 23581 17629 23615 17663
rect 13645 17561 13679 17595
rect 16497 17493 16531 17527
rect 19441 17493 19475 17527
rect 14013 17289 14047 17323
rect 15669 17289 15703 17323
rect 15853 17289 15887 17323
rect 17417 17289 17451 17323
rect 18337 17289 18371 17323
rect 21833 17289 21867 17323
rect 22109 17289 22143 17323
rect 22477 17289 22511 17323
rect 23121 17289 23155 17323
rect 23397 17289 23431 17323
rect 24961 17289 24995 17323
rect 12909 17221 12943 17255
rect 13645 17221 13679 17255
rect 13093 17153 13127 17187
rect 14381 17153 14415 17187
rect 16497 17153 16531 17187
rect 17141 17153 17175 17187
rect 18521 17153 18555 17187
rect 19165 17153 19199 17187
rect 20729 17153 20763 17187
rect 24041 17153 24075 17187
rect 15301 17085 15335 17119
rect 15460 17085 15494 17119
rect 20453 17085 20487 17119
rect 20913 17085 20947 17119
rect 12265 17017 12299 17051
rect 13185 17017 13219 17051
rect 16313 17017 16347 17051
rect 16589 17017 16623 17051
rect 18613 17017 18647 17051
rect 19533 17017 19567 17051
rect 21275 17017 21309 17051
rect 24133 17017 24167 17051
rect 24685 17017 24719 17051
rect 17877 16949 17911 16983
rect 19901 16949 19935 16983
rect 25513 16949 25547 16983
rect 11161 16745 11195 16779
rect 16957 16745 16991 16779
rect 17969 16745 18003 16779
rect 19717 16745 19751 16779
rect 21833 16745 21867 16779
rect 22201 16745 22235 16779
rect 24041 16745 24075 16779
rect 8125 16677 8159 16711
rect 8217 16677 8251 16711
rect 13185 16677 13219 16711
rect 17411 16677 17445 16711
rect 19118 16677 19152 16711
rect 19993 16677 20027 16711
rect 21159 16677 21193 16711
rect 23029 16677 23063 16711
rect 23581 16677 23615 16711
rect 24501 16677 24535 16711
rect 24593 16677 24627 16711
rect 11345 16609 11379 16643
rect 11621 16609 11655 16643
rect 16129 16609 16163 16643
rect 8769 16541 8803 16575
rect 13093 16541 13127 16575
rect 16221 16541 16255 16575
rect 17049 16541 17083 16575
rect 18797 16541 18831 16575
rect 20913 16541 20947 16575
rect 22937 16541 22971 16575
rect 24777 16541 24811 16575
rect 13645 16473 13679 16507
rect 9873 16405 9907 16439
rect 14013 16405 14047 16439
rect 18245 16405 18279 16439
rect 18705 16405 18739 16439
rect 20729 16405 20763 16439
rect 8953 16201 8987 16235
rect 13737 16201 13771 16235
rect 18475 16201 18509 16235
rect 23029 16201 23063 16235
rect 25145 16201 25179 16235
rect 7849 16133 7883 16167
rect 10149 16133 10183 16167
rect 12587 16133 12621 16167
rect 13461 16133 13495 16167
rect 19165 16133 19199 16167
rect 21097 16133 21131 16167
rect 23397 16133 23431 16167
rect 7113 16065 7147 16099
rect 8033 16065 8067 16099
rect 9597 16065 9631 16099
rect 11161 16065 11195 16099
rect 14013 16065 14047 16099
rect 15577 16065 15611 16099
rect 16497 16065 16531 16099
rect 17877 16065 17911 16099
rect 18797 16065 18831 16099
rect 22109 16065 22143 16099
rect 24225 16065 24259 16099
rect 24501 16065 24535 16099
rect 12484 15997 12518 16031
rect 18404 15997 18438 16031
rect 19625 15997 19659 16031
rect 19993 15997 20027 16031
rect 20177 15997 20211 16031
rect 20545 15997 20579 16031
rect 8125 15929 8159 15963
rect 8677 15929 8711 15963
rect 9413 15929 9447 15963
rect 9689 15929 9723 15963
rect 12173 15929 12207 15963
rect 13093 15929 13127 15963
rect 14105 15929 14139 15963
rect 14657 15929 14691 15963
rect 15669 15929 15703 15963
rect 16221 15929 16255 15963
rect 17509 15929 17543 15963
rect 21925 15929 21959 15963
rect 22201 15929 22235 15963
rect 22753 15929 22787 15963
rect 24317 15929 24351 15963
rect 7481 15861 7515 15895
rect 11345 15861 11379 15895
rect 11805 15861 11839 15895
rect 14933 15861 14967 15895
rect 15393 15861 15427 15895
rect 17141 15861 17175 15895
rect 19441 15861 19475 15895
rect 21465 15861 21499 15895
rect 24041 15861 24075 15895
rect 7849 15657 7883 15691
rect 9827 15657 9861 15691
rect 10425 15657 10459 15691
rect 15393 15657 15427 15691
rect 18613 15657 18647 15691
rect 20361 15657 20395 15691
rect 21005 15657 21039 15691
rect 23581 15657 23615 15691
rect 24133 15657 24167 15691
rect 24777 15657 24811 15691
rect 25145 15657 25179 15691
rect 8125 15589 8159 15623
rect 8217 15589 8251 15623
rect 11069 15589 11103 15623
rect 13829 15589 13863 15623
rect 14381 15589 14415 15623
rect 14841 15589 14875 15623
rect 17141 15589 17175 15623
rect 18061 15589 18095 15623
rect 24501 15589 24535 15623
rect 9597 15521 9631 15555
rect 12541 15521 12575 15555
rect 15301 15521 15335 15555
rect 15761 15521 15795 15555
rect 18797 15521 18831 15555
rect 19257 15521 19291 15555
rect 19533 15521 19567 15555
rect 19717 15521 19751 15555
rect 20913 15521 20947 15555
rect 21465 15521 21499 15555
rect 21741 15521 21775 15555
rect 22109 15521 22143 15555
rect 24961 15521 24995 15555
rect 8769 15453 8803 15487
rect 10977 15453 11011 15487
rect 11253 15453 11287 15487
rect 13737 15453 13771 15487
rect 16865 15453 16899 15487
rect 17049 15453 17083 15487
rect 17693 15453 17727 15487
rect 23213 15453 23247 15487
rect 12771 15385 12805 15419
rect 13461 15385 13495 15419
rect 18429 15385 18463 15419
rect 13093 15317 13127 15351
rect 16497 15317 16531 15351
rect 20729 15317 20763 15351
rect 9965 15113 9999 15147
rect 11437 15113 11471 15147
rect 12725 15113 12759 15147
rect 14749 15113 14783 15147
rect 17877 15113 17911 15147
rect 19257 15113 19291 15147
rect 24593 15113 24627 15147
rect 24961 15113 24995 15147
rect 25559 15113 25593 15147
rect 14013 15045 14047 15079
rect 15945 15045 15979 15079
rect 21097 15045 21131 15079
rect 23029 15045 23063 15079
rect 23397 15045 23431 15079
rect 8033 14977 8067 15011
rect 9229 14977 9263 15011
rect 10517 14977 10551 15011
rect 13093 14977 13127 15011
rect 15209 14977 15243 15011
rect 17141 14977 17175 15011
rect 18797 14977 18831 15011
rect 14289 14909 14323 14943
rect 19993 14909 20027 14943
rect 20177 14909 20211 14943
rect 20545 14909 20579 14943
rect 20913 14909 20947 14943
rect 22017 14909 22051 14943
rect 23673 14909 23707 14943
rect 25456 14909 25490 14943
rect 25881 14909 25915 14943
rect 7389 14841 7423 14875
rect 7481 14841 7515 14875
rect 8769 14841 8803 14875
rect 8953 14841 8987 14875
rect 9045 14841 9079 14875
rect 10609 14841 10643 14875
rect 11161 14841 11195 14875
rect 13455 14841 13489 14875
rect 14933 14841 14967 14875
rect 15025 14841 15059 14875
rect 16497 14841 16531 14875
rect 16589 14841 16623 14875
rect 17509 14841 17543 14875
rect 18153 14841 18187 14875
rect 18245 14841 18279 14875
rect 19533 14841 19567 14875
rect 21465 14841 21499 14875
rect 22569 14841 22603 14875
rect 7205 14773 7239 14807
rect 8401 14773 8435 14807
rect 10333 14773 10367 14807
rect 16313 14773 16347 14807
rect 21833 14773 21867 14807
rect 22201 14773 22235 14807
rect 24041 14773 24075 14807
rect 9689 14569 9723 14603
rect 10977 14569 11011 14603
rect 11437 14569 11471 14603
rect 11989 14569 12023 14603
rect 12633 14569 12667 14603
rect 14933 14569 14967 14603
rect 15439 14569 15473 14603
rect 17601 14569 17635 14603
rect 21097 14569 21131 14603
rect 23673 14569 23707 14603
rect 24133 14569 24167 14603
rect 8401 14501 8435 14535
rect 13093 14501 13127 14535
rect 13690 14501 13724 14535
rect 16681 14501 16715 14535
rect 17233 14501 17267 14535
rect 18245 14501 18279 14535
rect 23029 14501 23063 14535
rect 8636 14433 8670 14467
rect 11069 14433 11103 14467
rect 13369 14433 13403 14467
rect 15368 14433 15402 14467
rect 19625 14433 19659 14467
rect 20085 14433 20119 14467
rect 21741 14433 21775 14467
rect 22017 14433 22051 14467
rect 22385 14433 22419 14467
rect 22753 14433 22787 14467
rect 23949 14433 23983 14467
rect 25421 14433 25455 14467
rect 7389 14365 7423 14399
rect 8723 14365 8757 14399
rect 16589 14365 16623 14399
rect 18153 14365 18187 14399
rect 18429 14365 18463 14399
rect 17969 14297 18003 14331
rect 19349 14297 19383 14331
rect 20545 14297 20579 14331
rect 25605 14297 25639 14331
rect 7941 14229 7975 14263
rect 10149 14229 10183 14263
rect 14289 14229 14323 14263
rect 19809 14229 19843 14263
rect 23305 14229 23339 14263
rect 10425 14025 10459 14059
rect 10793 14025 10827 14059
rect 14289 14025 14323 14059
rect 15853 14025 15887 14059
rect 16221 14025 16255 14059
rect 17785 14025 17819 14059
rect 19165 14025 19199 14059
rect 21189 14025 21223 14059
rect 22937 14025 22971 14059
rect 23949 14025 23983 14059
rect 24363 14025 24397 14059
rect 11529 13957 11563 13991
rect 25697 13957 25731 13991
rect 8677 13889 8711 13923
rect 9505 13889 9539 13923
rect 13185 13889 13219 13923
rect 14473 13889 14507 13923
rect 16497 13889 16531 13923
rect 17141 13889 17175 13923
rect 26065 13889 26099 13923
rect 7941 13821 7975 13855
rect 8401 13821 8435 13855
rect 11345 13821 11379 13855
rect 12725 13821 12759 13855
rect 13001 13821 13035 13855
rect 18188 13821 18222 13855
rect 18613 13821 18647 13855
rect 19533 13821 19567 13855
rect 19717 13821 19751 13855
rect 20085 13821 20119 13855
rect 20453 13821 20487 13855
rect 22144 13821 22178 13855
rect 22569 13821 22603 13855
rect 25288 13821 25322 13855
rect 25375 13821 25409 13855
rect 9867 13753 9901 13787
rect 11161 13753 11195 13787
rect 11897 13753 11931 13787
rect 12265 13753 12299 13787
rect 13645 13753 13679 13787
rect 14565 13753 14599 13787
rect 15117 13753 15151 13787
rect 16589 13753 16623 13787
rect 7849 13685 7883 13719
rect 8953 13685 8987 13719
rect 9413 13685 9447 13719
rect 15393 13685 15427 13719
rect 17417 13685 17451 13719
rect 18291 13685 18325 13719
rect 19349 13685 19383 13719
rect 21557 13685 21591 13719
rect 21925 13685 21959 13719
rect 22247 13685 22281 13719
rect 24133 13685 24167 13719
rect 24685 13685 24719 13719
rect 13829 13481 13863 13515
rect 14657 13481 14691 13515
rect 16957 13481 16991 13515
rect 19349 13481 19383 13515
rect 19901 13481 19935 13515
rect 21281 13481 21315 13515
rect 25467 13481 25501 13515
rect 9873 13413 9907 13447
rect 15761 13413 15795 13447
rect 18331 13413 18365 13447
rect 22937 13413 22971 13447
rect 8309 13345 8343 13379
rect 8493 13345 8527 13379
rect 11304 13345 11338 13379
rect 12725 13345 12759 13379
rect 13001 13345 13035 13379
rect 17969 13345 18003 13379
rect 19717 13345 19751 13379
rect 21741 13345 21775 13379
rect 21925 13345 21959 13379
rect 22293 13345 22327 13379
rect 22661 13345 22695 13379
rect 24133 13345 24167 13379
rect 25396 13345 25430 13379
rect 8769 13277 8803 13311
rect 9781 13277 9815 13311
rect 11391 13277 11425 13311
rect 13185 13277 13219 13311
rect 13461 13277 13495 13311
rect 14197 13277 14231 13311
rect 15669 13277 15703 13311
rect 15945 13277 15979 13311
rect 10333 13209 10367 13243
rect 10885 13141 10919 13175
rect 16681 13141 16715 13175
rect 18889 13141 18923 13175
rect 20269 13141 20303 13175
rect 20637 13141 20671 13175
rect 24041 13141 24075 13175
rect 9321 12937 9355 12971
rect 9965 12937 9999 12971
rect 13829 12937 13863 12971
rect 14749 12937 14783 12971
rect 14841 12937 14875 12971
rect 16037 12937 16071 12971
rect 17509 12937 17543 12971
rect 12173 12869 12207 12903
rect 8309 12801 8343 12835
rect 11253 12801 11287 12835
rect 12909 12801 12943 12835
rect 6837 12733 6871 12767
rect 7389 12733 7423 12767
rect 7573 12733 7607 12767
rect 8401 12733 8435 12767
rect 7941 12665 7975 12699
rect 8723 12665 8757 12699
rect 10885 12665 10919 12699
rect 10977 12665 11011 12699
rect 12817 12665 12851 12699
rect 13271 12665 13305 12699
rect 18429 12869 18463 12903
rect 24777 12869 24811 12903
rect 15117 12801 15151 12835
rect 15485 12801 15519 12835
rect 16405 12801 16439 12835
rect 16589 12801 16623 12835
rect 18797 12801 18831 12835
rect 23857 12801 23891 12835
rect 24225 12801 24259 12835
rect 25329 12801 25363 12835
rect 17877 12733 17911 12767
rect 18245 12733 18279 12767
rect 19257 12733 19291 12767
rect 19717 12733 19751 12767
rect 20269 12733 20303 12767
rect 20453 12733 20487 12767
rect 15209 12665 15243 12699
rect 22109 12665 22143 12699
rect 22201 12665 22235 12699
rect 22753 12665 22787 12699
rect 23949 12665 23983 12699
rect 6653 12597 6687 12631
rect 9689 12597 9723 12631
rect 10701 12597 10735 12631
rect 11897 12597 11931 12631
rect 14749 12597 14783 12631
rect 19073 12597 19107 12631
rect 19349 12597 19383 12631
rect 21005 12597 21039 12631
rect 21465 12597 21499 12631
rect 21925 12597 21959 12631
rect 23029 12597 23063 12631
rect 23489 12597 23523 12631
rect 25789 12597 25823 12631
rect 6929 12393 6963 12427
rect 9045 12393 9079 12427
rect 9965 12393 9999 12427
rect 10241 12393 10275 12427
rect 11437 12393 11471 12427
rect 13921 12393 13955 12427
rect 15117 12393 15151 12427
rect 16221 12393 16255 12427
rect 17969 12393 18003 12427
rect 18797 12393 18831 12427
rect 22937 12393 22971 12427
rect 24041 12393 24075 12427
rect 24317 12393 24351 12427
rect 10838 12325 10872 12359
rect 13363 12325 13397 12359
rect 15663 12325 15697 12359
rect 17325 12325 17359 12359
rect 18429 12325 18463 12359
rect 21735 12325 21769 12359
rect 23442 12325 23476 12359
rect 25053 12325 25087 12359
rect 8033 12257 8067 12291
rect 8493 12257 8527 12291
rect 10517 12257 10551 12291
rect 19257 12257 19291 12291
rect 19533 12257 19567 12291
rect 22293 12257 22327 12291
rect 8585 12189 8619 12223
rect 13001 12189 13035 12223
rect 15301 12189 15335 12223
rect 17049 12189 17083 12223
rect 19717 12189 19751 12223
rect 21097 12189 21131 12223
rect 21373 12189 21407 12223
rect 22569 12189 22603 12223
rect 23121 12189 23155 12223
rect 24961 12189 24995 12223
rect 25237 12189 25271 12223
rect 19349 12121 19383 12155
rect 20729 12121 20763 12155
rect 24777 12121 24811 12155
rect 12541 12053 12575 12087
rect 19073 12053 19107 12087
rect 7665 11849 7699 11883
rect 10149 11849 10183 11883
rect 12817 11849 12851 11883
rect 13921 11849 13955 11883
rect 14749 11849 14783 11883
rect 17785 11849 17819 11883
rect 19763 11849 19797 11883
rect 24869 11849 24903 11883
rect 8309 11781 8343 11815
rect 11161 11781 11195 11815
rect 15577 11781 15611 11815
rect 16037 11781 16071 11815
rect 20637 11781 20671 11815
rect 25697 11781 25731 11815
rect 8493 11713 8527 11747
rect 15025 11713 15059 11747
rect 16313 11713 16347 11747
rect 16635 11713 16669 11747
rect 18061 11713 18095 11747
rect 19349 11713 19383 11747
rect 23765 11713 23799 11747
rect 24225 11713 24259 11747
rect 10241 11645 10275 11679
rect 12265 11645 12299 11679
rect 13001 11645 13035 11679
rect 16548 11645 16582 11679
rect 18153 11645 18187 11679
rect 19660 11645 19694 11679
rect 20085 11645 20119 11679
rect 20913 11645 20947 11679
rect 21189 11645 21223 11679
rect 21741 11645 21775 11679
rect 22017 11645 22051 11679
rect 8814 11577 8848 11611
rect 10562 11577 10596 11611
rect 13322 11577 13356 11611
rect 15117 11577 15151 11611
rect 17417 11577 17451 11611
rect 22201 11577 22235 11611
rect 23857 11577 23891 11611
rect 8033 11509 8067 11543
rect 9413 11509 9447 11543
rect 9689 11509 9723 11543
rect 14473 11509 14507 11543
rect 17049 11509 17083 11543
rect 22477 11509 22511 11543
rect 23121 11509 23155 11543
rect 25237 11509 25271 11543
rect 9045 11305 9079 11339
rect 10701 11305 10735 11339
rect 13093 11305 13127 11339
rect 13737 11305 13771 11339
rect 17601 11305 17635 11339
rect 19073 11305 19107 11339
rect 21189 11305 21223 11339
rect 22661 11305 22695 11339
rect 23029 11305 23063 11339
rect 24225 11305 24259 11339
rect 24915 11305 24949 11339
rect 8769 11237 8803 11271
rect 9873 11237 9907 11271
rect 12173 11237 12207 11271
rect 12265 11237 12299 11271
rect 15485 11237 15519 11271
rect 17877 11237 17911 11271
rect 7021 11169 7055 11203
rect 8033 11169 8067 11203
rect 8585 11169 8619 11203
rect 13737 11169 13771 11203
rect 14105 11169 14139 11203
rect 18981 11169 19015 11203
rect 19257 11169 19291 11203
rect 19717 11169 19751 11203
rect 20729 11169 20763 11203
rect 20913 11169 20947 11203
rect 21373 11169 21407 11203
rect 21741 11169 21775 11203
rect 22109 11169 22143 11203
rect 23305 11169 23339 11203
rect 24844 11169 24878 11203
rect 9781 11101 9815 11135
rect 10241 11101 10275 11135
rect 12817 11101 12851 11135
rect 15393 11101 15427 11135
rect 15669 11101 15703 11135
rect 17785 11101 17819 11135
rect 13461 11033 13495 11067
rect 18337 11033 18371 11067
rect 19809 11101 19843 11135
rect 23949 11101 23983 11135
rect 7205 10965 7239 10999
rect 9413 10965 9447 10999
rect 15025 10965 15059 10999
rect 16313 10965 16347 10999
rect 17233 10965 17267 10999
rect 18705 10965 18739 10999
rect 18981 10965 19015 10999
rect 24685 10965 24719 10999
rect 6653 10761 6687 10795
rect 9413 10761 9447 10795
rect 10609 10761 10643 10795
rect 11161 10761 11195 10795
rect 12265 10761 12299 10795
rect 15761 10761 15795 10795
rect 21005 10761 21039 10795
rect 22293 10761 22327 10795
rect 9045 10693 9079 10727
rect 10241 10693 10275 10727
rect 15577 10693 15611 10727
rect 17509 10693 17543 10727
rect 18981 10693 19015 10727
rect 19901 10693 19935 10727
rect 21649 10693 21683 10727
rect 7849 10625 7883 10659
rect 8769 10625 8803 10659
rect 12541 10625 12575 10659
rect 12817 10625 12851 10659
rect 7056 10557 7090 10591
rect 8033 10557 8067 10591
rect 8585 10557 8619 10591
rect 11380 10557 11414 10591
rect 11805 10557 11839 10591
rect 14105 10557 14139 10591
rect 14657 10557 14691 10591
rect 14749 10557 14783 10591
rect 15209 10557 15243 10591
rect 20269 10625 20303 10659
rect 24317 10625 24351 10659
rect 24961 10625 24995 10659
rect 16313 10557 16347 10591
rect 16773 10557 16807 10591
rect 18061 10557 18095 10591
rect 19809 10557 19843 10591
rect 20085 10557 20119 10591
rect 22661 10557 22695 10591
rect 7159 10489 7193 10523
rect 9689 10489 9723 10523
rect 9781 10489 9815 10523
rect 11483 10489 11517 10523
rect 12633 10489 12667 10523
rect 15577 10489 15611 10523
rect 16221 10489 16255 10523
rect 17877 10489 17911 10523
rect 18423 10489 18457 10523
rect 24409 10489 24443 10523
rect 7573 10421 7607 10455
rect 13645 10421 13679 10455
rect 14841 10421 14875 10455
rect 16405 10421 16439 10455
rect 19257 10421 19291 10455
rect 19625 10421 19659 10455
rect 21281 10421 21315 10455
rect 23213 10421 23247 10455
rect 24133 10421 24167 10455
rect 25237 10421 25271 10455
rect 7159 10217 7193 10251
rect 9505 10217 9539 10251
rect 9873 10217 9907 10251
rect 11529 10217 11563 10251
rect 12633 10217 12667 10251
rect 12909 10217 12943 10251
rect 16405 10217 16439 10251
rect 18337 10217 18371 10251
rect 18889 10217 18923 10251
rect 21373 10217 21407 10251
rect 10885 10149 10919 10183
rect 12075 10149 12109 10183
rect 13553 10149 13587 10183
rect 13645 10149 13679 10183
rect 15847 10149 15881 10183
rect 17417 10149 17451 10183
rect 22937 10149 22971 10183
rect 23489 10149 23523 10183
rect 24501 10149 24535 10183
rect 6076 10081 6110 10115
rect 7021 10081 7055 10115
rect 8033 10081 8067 10115
rect 8585 10081 8619 10115
rect 10149 10081 10183 10115
rect 10609 10081 10643 10115
rect 11713 10081 11747 10115
rect 13277 10081 13311 10115
rect 15485 10081 15519 10115
rect 19073 10081 19107 10115
rect 19257 10081 19291 10115
rect 20913 10081 20947 10115
rect 21189 10081 21223 10115
rect 7941 10013 7975 10047
rect 8769 10013 8803 10047
rect 17325 10013 17359 10047
rect 17969 10013 18003 10047
rect 21925 10013 21959 10047
rect 22845 10013 22879 10047
rect 24409 10013 24443 10047
rect 6147 9945 6181 9979
rect 14105 9945 14139 9979
rect 20637 9945 20671 9979
rect 21005 9945 21039 9979
rect 24961 9945 24995 9979
rect 14749 9877 14783 9911
rect 17049 9877 17083 9911
rect 19901 9877 19935 9911
rect 20269 9877 20303 9911
rect 22293 9877 22327 9911
rect 6009 9673 6043 9707
rect 6285 9673 6319 9707
rect 7113 9673 7147 9707
rect 8125 9673 8159 9707
rect 8493 9673 8527 9707
rect 9873 9673 9907 9707
rect 10149 9673 10183 9707
rect 11805 9673 11839 9707
rect 12265 9673 12299 9707
rect 13369 9673 13403 9707
rect 13645 9673 13679 9707
rect 14795 9673 14829 9707
rect 17233 9673 17267 9707
rect 19073 9673 19107 9707
rect 23489 9673 23523 9707
rect 24225 9673 24259 9707
rect 4859 9537 4893 9571
rect 6653 9605 6687 9639
rect 14013 9605 14047 9639
rect 14933 9605 14967 9639
rect 15209 9605 15243 9639
rect 25421 9605 25455 9639
rect 10425 9537 10459 9571
rect 12449 9537 12483 9571
rect 16037 9537 16071 9571
rect 18153 9537 18187 9571
rect 18797 9537 18831 9571
rect 21833 9537 21867 9571
rect 24501 9537 24535 9571
rect 24961 9537 24995 9571
rect 4772 9469 4806 9503
rect 5800 9469 5834 9503
rect 6009 9469 6043 9503
rect 7624 9469 7658 9503
rect 8585 9469 8619 9503
rect 14724 9469 14758 9503
rect 14933 9469 14967 9503
rect 19441 9469 19475 9503
rect 20269 9469 20303 9503
rect 7711 9401 7745 9435
rect 8947 9401 8981 9435
rect 10517 9401 10551 9435
rect 11069 9401 11103 9435
rect 12770 9401 12804 9435
rect 15761 9401 15795 9435
rect 15853 9401 15887 9435
rect 18245 9401 18279 9435
rect 19625 9401 19659 9435
rect 21005 9401 21039 9435
rect 21741 9401 21775 9435
rect 22195 9401 22229 9435
rect 23949 9401 23983 9435
rect 24593 9401 24627 9435
rect 5181 9333 5215 9367
rect 5871 9333 5905 9367
rect 7481 9333 7515 9367
rect 9505 9333 9539 9367
rect 11345 9333 11379 9367
rect 15577 9333 15611 9367
rect 16681 9333 16715 9367
rect 17877 9333 17911 9367
rect 21373 9333 21407 9367
rect 22753 9333 22787 9367
rect 23121 9333 23155 9367
rect 10701 9129 10735 9163
rect 11069 9129 11103 9163
rect 11345 9129 11379 9163
rect 12449 9129 12483 9163
rect 15117 9129 15151 9163
rect 15669 9129 15703 9163
rect 16221 9129 16255 9163
rect 16497 9129 16531 9163
rect 17969 9129 18003 9163
rect 20361 9129 20395 9163
rect 20637 9129 20671 9163
rect 24685 9129 24719 9163
rect 7205 9061 7239 9095
rect 9045 9061 9079 9095
rect 9781 9061 9815 9095
rect 9873 9061 9907 9095
rect 13553 9061 13587 9095
rect 14105 9061 14139 9095
rect 17370 9061 17404 9095
rect 18797 9061 18831 9095
rect 23718 9061 23752 9095
rect 5457 8993 5491 9027
rect 6561 8993 6595 9027
rect 7021 8993 7055 9027
rect 8033 8993 8067 9027
rect 8493 8993 8527 9027
rect 11437 8993 11471 9027
rect 11805 8993 11839 9027
rect 15301 8993 15335 9027
rect 19165 8993 19199 9027
rect 19441 8993 19475 9027
rect 21097 8993 21131 9027
rect 21557 8993 21591 9027
rect 21925 8993 21959 9027
rect 22293 8993 22327 9027
rect 7481 8925 7515 8959
rect 8585 8925 8619 8959
rect 13461 8925 13495 8959
rect 17049 8925 17083 8959
rect 19625 8925 19659 8959
rect 22569 8925 22603 8959
rect 23397 8925 23431 8959
rect 25145 8925 25179 8959
rect 5641 8857 5675 8891
rect 10333 8857 10367 8891
rect 19257 8857 19291 8891
rect 16865 8789 16899 8823
rect 18245 8789 18279 8823
rect 24317 8789 24351 8823
rect 10057 8585 10091 8619
rect 12817 8585 12851 8619
rect 13185 8585 13219 8619
rect 15117 8585 15151 8619
rect 15945 8585 15979 8619
rect 17233 8585 17267 8619
rect 19717 8585 19751 8619
rect 20361 8585 20395 8619
rect 23121 8585 23155 8619
rect 24685 8585 24719 8619
rect 8493 8449 8527 8483
rect 10885 8449 10919 8483
rect 12173 8449 12207 8483
rect 13461 8449 13495 8483
rect 15347 8449 15381 8483
rect 18199 8517 18233 8551
rect 25421 8517 25455 8551
rect 16313 8449 16347 8483
rect 22293 8449 22327 8483
rect 24041 8449 24075 8483
rect 5181 8381 5215 8415
rect 5733 8381 5767 8415
rect 6929 8381 6963 8415
rect 7481 8381 7515 8415
rect 15244 8381 15278 8415
rect 15945 8381 15979 8415
rect 16037 8381 16071 8415
rect 18128 8381 18162 8415
rect 19165 8381 19199 8415
rect 19901 8381 19935 8415
rect 20821 8381 20855 8415
rect 21281 8381 21315 8415
rect 21649 8381 21683 8415
rect 22017 8381 22051 8415
rect 25237 8381 25271 8415
rect 5549 8313 5583 8347
rect 7665 8313 7699 8347
rect 8401 8313 8435 8347
rect 8855 8313 8889 8347
rect 10977 8313 11011 8347
rect 11529 8313 11563 8347
rect 13553 8313 13587 8347
rect 14105 8313 14139 8347
rect 16405 8313 16439 8347
rect 16957 8313 16991 8347
rect 23765 8313 23799 8347
rect 23857 8313 23891 8347
rect 5917 8245 5951 8279
rect 6561 8245 6595 8279
rect 8033 8245 8067 8279
rect 9413 8245 9447 8279
rect 9689 8245 9723 8279
rect 10701 8245 10735 8279
rect 11897 8245 11931 8279
rect 14381 8245 14415 8279
rect 15669 8245 15703 8279
rect 17693 8245 17727 8279
rect 18521 8245 18555 8279
rect 20637 8245 20671 8279
rect 22569 8245 22603 8279
rect 23489 8245 23523 8279
rect 25697 8245 25731 8279
rect 7113 8041 7147 8075
rect 7481 8041 7515 8075
rect 8953 8041 8987 8075
rect 9781 8041 9815 8075
rect 10793 8041 10827 8075
rect 13185 8041 13219 8075
rect 16773 8041 16807 8075
rect 18613 8041 18647 8075
rect 19533 8041 19567 8075
rect 19993 8041 20027 8075
rect 20269 8041 20303 8075
rect 21097 8041 21131 8075
rect 22109 8041 22143 8075
rect 24501 8041 24535 8075
rect 7757 7973 7791 8007
rect 8677 7973 8711 8007
rect 11621 7973 11655 8007
rect 13553 7973 13587 8007
rect 14105 7973 14139 8007
rect 17141 7973 17175 8007
rect 21373 7973 21407 8007
rect 23305 7973 23339 8007
rect 24225 7973 24259 8007
rect 24685 7973 24719 8007
rect 5549 7905 5583 7939
rect 6561 7905 6595 7939
rect 9689 7905 9723 7939
rect 10241 7905 10275 7939
rect 15669 7905 15703 7939
rect 15945 7905 15979 7939
rect 18797 7905 18831 7939
rect 18981 7905 19015 7939
rect 20913 7905 20947 7939
rect 21741 7905 21775 7939
rect 21925 7905 21959 7939
rect 23857 7905 23891 7939
rect 25237 7905 25271 7939
rect 7665 7837 7699 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 12449 7837 12483 7871
rect 13461 7837 13495 7871
rect 16129 7837 16163 7871
rect 17049 7837 17083 7871
rect 17325 7837 17359 7871
rect 23213 7837 23247 7871
rect 6745 7769 6779 7803
rect 8217 7769 8251 7803
rect 18061 7769 18095 7803
rect 5733 7701 5767 7735
rect 11253 7701 11287 7735
rect 14473 7701 14507 7735
rect 16405 7701 16439 7735
rect 20637 7701 20671 7735
rect 22477 7701 22511 7735
rect 5917 7497 5951 7531
rect 6653 7497 6687 7531
rect 7665 7497 7699 7531
rect 10149 7497 10183 7531
rect 11529 7497 11563 7531
rect 11805 7497 11839 7531
rect 13553 7497 13587 7531
rect 13829 7497 13863 7531
rect 15485 7497 15519 7531
rect 17141 7497 17175 7531
rect 17877 7497 17911 7531
rect 18521 7497 18555 7531
rect 24869 7497 24903 7531
rect 25237 7497 25271 7531
rect 25881 7497 25915 7531
rect 15853 7429 15887 7463
rect 19073 7429 19107 7463
rect 19993 7429 20027 7463
rect 20361 7429 20395 7463
rect 20637 7429 20671 7463
rect 22293 7429 22327 7463
rect 7205 7361 7239 7395
rect 8217 7361 8251 7395
rect 10609 7361 10643 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 16221 7361 16255 7395
rect 19441 7361 19475 7395
rect 21925 7361 21959 7395
rect 23949 7361 23983 7395
rect 5733 7293 5767 7327
rect 14657 7293 14691 7327
rect 14933 7293 14967 7327
rect 18981 7293 19015 7327
rect 19257 7293 19291 7327
rect 20545 7293 20579 7327
rect 20821 7293 20855 7327
rect 22109 7293 22143 7327
rect 25488 7293 25522 7327
rect 8125 7225 8159 7259
rect 8579 7225 8613 7259
rect 10517 7225 10551 7259
rect 10971 7225 11005 7259
rect 12633 7225 12667 7259
rect 14289 7225 14323 7259
rect 16313 7225 16347 7259
rect 16865 7225 16899 7259
rect 18889 7225 18923 7259
rect 21557 7225 21591 7259
rect 24041 7225 24075 7259
rect 24593 7225 24627 7259
rect 5641 7157 5675 7191
rect 6285 7157 6319 7191
rect 9137 7157 9171 7191
rect 9689 7157 9723 7191
rect 12265 7157 12299 7191
rect 14473 7157 14507 7191
rect 21005 7157 21039 7191
rect 22569 7157 22603 7191
rect 22937 7157 22971 7191
rect 23489 7157 23523 7191
rect 25559 7157 25593 7191
rect 7665 6953 7699 6987
rect 8217 6953 8251 6987
rect 9045 6953 9079 6987
rect 12357 6953 12391 6987
rect 12909 6953 12943 6987
rect 14657 6953 14691 6987
rect 15669 6953 15703 6987
rect 16497 6953 16531 6987
rect 18705 6953 18739 6987
rect 20545 6953 20579 6987
rect 23581 6953 23615 6987
rect 6469 6885 6503 6919
rect 8861 6885 8895 6919
rect 10333 6885 10367 6919
rect 17233 6885 17267 6919
rect 19210 6885 19244 6919
rect 14013 6817 14047 6851
rect 20085 6817 20119 6851
rect 20913 6817 20947 6851
rect 21373 6817 21407 6851
rect 21741 6817 21775 6851
rect 22109 6817 22143 6851
rect 24961 6817 24995 6851
rect 5181 6749 5215 6783
rect 6377 6749 6411 6783
rect 7021 6749 7055 6783
rect 7757 6749 7791 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 11989 6749 12023 6783
rect 15301 6749 15335 6783
rect 17141 6749 17175 6783
rect 17417 6749 17451 6783
rect 18889 6749 18923 6783
rect 22385 6749 22419 6783
rect 23213 6749 23247 6783
rect 5411 6681 5445 6715
rect 14197 6681 14231 6715
rect 9873 6613 9907 6647
rect 11437 6613 11471 6647
rect 16221 6613 16255 6647
rect 16957 6613 16991 6647
rect 19809 6613 19843 6647
rect 22661 6613 22695 6647
rect 23029 6613 23063 6647
rect 24133 6613 24167 6647
rect 24409 6613 24443 6647
rect 25099 6613 25133 6647
rect 4905 6409 4939 6443
rect 8309 6409 8343 6443
rect 10885 6409 10919 6443
rect 12081 6409 12115 6443
rect 14013 6409 14047 6443
rect 17785 6409 17819 6443
rect 18981 6409 19015 6443
rect 25053 6409 25087 6443
rect 4629 6341 4663 6375
rect 5871 6341 5905 6375
rect 10517 6341 10551 6375
rect 18199 6341 18233 6375
rect 24317 6341 24351 6375
rect 5365 6273 5399 6307
rect 6561 6273 6595 6307
rect 6929 6273 6963 6307
rect 7573 6273 7607 6307
rect 7941 6273 7975 6307
rect 9689 6273 9723 6307
rect 9965 6273 9999 6307
rect 11713 6273 11747 6307
rect 13737 6273 13771 6307
rect 14381 6273 14415 6307
rect 16129 6273 16163 6307
rect 21281 6273 21315 6307
rect 22477 6273 22511 6307
rect 4721 6205 4755 6239
rect 5800 6205 5834 6239
rect 8896 6205 8930 6239
rect 8999 6205 9033 6239
rect 12449 6205 12483 6239
rect 12909 6205 12943 6239
rect 15301 6205 15335 6239
rect 17325 6205 17359 6239
rect 18128 6205 18162 6239
rect 19809 6205 19843 6239
rect 19993 6205 20027 6239
rect 20361 6205 20395 6239
rect 20729 6205 20763 6239
rect 22017 6205 22051 6239
rect 22109 6205 22143 6239
rect 22293 6205 22327 6239
rect 25272 6205 25306 6239
rect 25697 6205 25731 6239
rect 7021 6137 7055 6171
rect 9413 6137 9447 6171
rect 10057 6137 10091 6171
rect 11345 6137 11379 6171
rect 14743 6137 14777 6171
rect 15669 6137 15703 6171
rect 16037 6137 16071 6171
rect 16491 6137 16525 6171
rect 21925 6137 21959 6171
rect 23765 6137 23799 6171
rect 23857 6137 23891 6171
rect 6285 6069 6319 6103
rect 12541 6069 12575 6103
rect 17049 6069 17083 6103
rect 18613 6069 18647 6103
rect 19349 6069 19383 6103
rect 19625 6069 19659 6103
rect 23305 6069 23339 6103
rect 25375 6069 25409 6103
rect 6929 5865 6963 5899
rect 7159 5865 7193 5899
rect 10701 5865 10735 5899
rect 12725 5865 12759 5899
rect 16405 5865 16439 5899
rect 18429 5865 18463 5899
rect 19993 5865 20027 5899
rect 22661 5865 22695 5899
rect 23305 5865 23339 5899
rect 24041 5865 24075 5899
rect 8217 5797 8251 5831
rect 8769 5797 8803 5831
rect 9873 5797 9907 5831
rect 11897 5797 11931 5831
rect 16773 5797 16807 5831
rect 16865 5797 16899 5831
rect 18705 5797 18739 5831
rect 19533 5797 19567 5831
rect 20637 5797 20671 5831
rect 1409 5729 1443 5763
rect 5064 5729 5098 5763
rect 6009 5729 6043 5763
rect 7056 5729 7090 5763
rect 10425 5729 10459 5763
rect 13921 5729 13955 5763
rect 14105 5729 14139 5763
rect 15301 5729 15335 5763
rect 20269 5729 20303 5763
rect 21373 5729 21407 5763
rect 22477 5729 22511 5763
rect 24225 5729 24259 5763
rect 25212 5729 25246 5763
rect 1547 5661 1581 5695
rect 8125 5661 8159 5695
rect 9413 5661 9447 5695
rect 9781 5661 9815 5695
rect 11805 5661 11839 5695
rect 12449 5661 12483 5695
rect 14197 5661 14231 5695
rect 17049 5661 17083 5695
rect 18613 5661 18647 5695
rect 19257 5661 19291 5695
rect 23029 5661 23063 5695
rect 24593 5661 24627 5695
rect 6147 5593 6181 5627
rect 15853 5593 15887 5627
rect 25283 5593 25317 5627
rect 5135 5525 5169 5559
rect 6469 5525 6503 5559
rect 7481 5525 7515 5559
rect 9137 5525 9171 5559
rect 11437 5525 11471 5559
rect 15485 5525 15519 5559
rect 17969 5525 18003 5559
rect 21373 5525 21407 5559
rect 22109 5525 22143 5559
rect 3295 5321 3329 5355
rect 8309 5321 8343 5355
rect 9689 5321 9723 5355
rect 10057 5321 10091 5355
rect 15577 5321 15611 5355
rect 17417 5321 17451 5355
rect 17877 5321 17911 5355
rect 19809 5321 19843 5355
rect 21373 5321 21407 5355
rect 23029 5321 23063 5355
rect 25053 5321 25087 5355
rect 5273 5253 5307 5287
rect 6285 5253 6319 5287
rect 13645 5253 13679 5287
rect 20453 5253 20487 5287
rect 11529 5185 11563 5219
rect 18889 5185 18923 5219
rect 21925 5185 21959 5219
rect 22569 5185 22603 5219
rect 24133 5185 24167 5219
rect 3224 5117 3258 5151
rect 4788 5117 4822 5151
rect 5784 5117 5818 5151
rect 5871 5117 5905 5151
rect 7021 5117 7055 5151
rect 7389 5117 7423 5151
rect 7941 5117 7975 5151
rect 8493 5117 8527 5151
rect 10701 5117 10735 5151
rect 10977 5117 11011 5151
rect 11253 5117 11287 5151
rect 14473 5117 14507 5151
rect 14565 5117 14599 5151
rect 15025 5117 15059 5151
rect 16313 5117 16347 5151
rect 16497 5117 16531 5151
rect 16865 5117 16899 5151
rect 19533 5117 19567 5151
rect 20361 5117 20395 5151
rect 20637 5117 20671 5151
rect 22017 5117 22051 5151
rect 22109 5117 22143 5151
rect 22293 5117 22327 5151
rect 23673 5117 23707 5151
rect 23765 5117 23799 5151
rect 23949 5117 23983 5151
rect 7665 5049 7699 5083
rect 8814 5049 8848 5083
rect 12173 5049 12207 5083
rect 12541 5049 12575 5083
rect 12633 5049 12667 5083
rect 13185 5049 13219 5083
rect 15301 5049 15335 5083
rect 17141 5049 17175 5083
rect 18981 5049 19015 5083
rect 20269 5049 20303 5083
rect 23489 5049 23523 5083
rect 25237 5049 25271 5083
rect 25789 5049 25823 5083
rect 1593 4981 1627 5015
rect 3709 4981 3743 5015
rect 4859 4981 4893 5015
rect 5549 4981 5583 5015
rect 6653 4981 6687 5015
rect 9413 4981 9447 5015
rect 11897 4981 11931 5015
rect 14013 4981 14047 5015
rect 18521 4981 18555 5015
rect 20821 4981 20855 5015
rect 24685 4981 24719 5015
rect 4583 4777 4617 4811
rect 7849 4777 7883 4811
rect 8309 4777 8343 4811
rect 9045 4777 9079 4811
rect 10885 4777 10919 4811
rect 12909 4777 12943 4811
rect 14657 4777 14691 4811
rect 15669 4777 15703 4811
rect 16957 4777 16991 4811
rect 19533 4777 19567 4811
rect 19993 4777 20027 4811
rect 20453 4777 20487 4811
rect 9505 4709 9539 4743
rect 9965 4709 9999 4743
rect 11707 4709 11741 4743
rect 13277 4709 13311 4743
rect 18521 4709 18555 4743
rect 4512 4641 4546 4675
rect 5457 4641 5491 4675
rect 6009 4641 6043 4675
rect 6745 4641 6779 4675
rect 7021 4641 7055 4675
rect 7481 4641 7515 4675
rect 8217 4641 8251 4675
rect 8493 4641 8527 4675
rect 10517 4641 10551 4675
rect 17049 4641 17083 4675
rect 19165 4641 19199 4675
rect 20913 4641 20947 4675
rect 23029 4641 23063 4675
rect 23765 4641 23799 4675
rect 23949 4641 23983 4675
rect 24593 4641 24627 4675
rect 7205 4573 7239 4607
rect 9873 4573 9907 4607
rect 11345 4573 11379 4607
rect 12541 4573 12575 4607
rect 13185 4573 13219 4607
rect 13553 4573 13587 4607
rect 15301 4573 15335 4607
rect 22109 4573 22143 4607
rect 23121 4573 23155 4607
rect 5595 4505 5629 4539
rect 11161 4505 11195 4539
rect 18153 4505 18187 4539
rect 12265 4437 12299 4471
rect 16221 4437 16255 4471
rect 16589 4437 16623 4471
rect 17233 4437 17267 4471
rect 21097 4437 21131 4471
rect 21557 4437 21591 4471
rect 3617 4233 3651 4267
rect 3985 4233 4019 4267
rect 5549 4233 5583 4267
rect 9781 4233 9815 4267
rect 11897 4233 11931 4267
rect 16221 4233 16255 4267
rect 19165 4233 19199 4267
rect 20913 4233 20947 4267
rect 21281 4233 21315 4267
rect 22845 4233 22879 4267
rect 25421 4233 25455 4267
rect 4629 4165 4663 4199
rect 5871 4165 5905 4199
rect 8401 4165 8435 4199
rect 14105 4165 14139 4199
rect 14381 4165 14415 4199
rect 19809 4165 19843 4199
rect 19993 4165 20027 4199
rect 21557 4165 21591 4199
rect 22569 4165 22603 4199
rect 23765 4165 23799 4199
rect 7665 4097 7699 4131
rect 13185 4097 13219 4131
rect 14565 4097 14599 4131
rect 16405 4097 16439 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 18153 4097 18187 4131
rect 18429 4097 18463 4131
rect 22201 4097 22235 4131
rect 25053 4097 25087 4131
rect 3776 4029 3810 4063
rect 4756 4029 4790 4063
rect 5800 4029 5834 4063
rect 6929 4029 6963 4063
rect 7389 4029 7423 4063
rect 7941 4029 7975 4063
rect 8493 4029 8527 4063
rect 10057 4029 10091 4063
rect 19901 4029 19935 4063
rect 20177 4029 20211 4063
rect 21465 4029 21499 4063
rect 21741 4029 21775 4063
rect 23673 4029 23707 4063
rect 23949 4029 23983 4063
rect 24409 4029 24443 4063
rect 25237 4029 25271 4063
rect 25697 4029 25731 4063
rect 6653 3961 6687 3995
rect 8814 3961 8848 3995
rect 10885 3961 10919 3995
rect 10977 3961 11011 3995
rect 11529 3961 11563 3995
rect 12541 3961 12575 3995
rect 12633 3961 12667 3995
rect 13461 3961 13495 3995
rect 14927 3961 14961 3995
rect 16497 3961 16531 3995
rect 17877 3961 17911 3995
rect 18245 3961 18279 3995
rect 20637 3961 20671 3995
rect 4261 3893 4295 3927
rect 4859 3893 4893 3927
rect 6285 3893 6319 3927
rect 9413 3893 9447 3927
rect 10701 3893 10735 3927
rect 12173 3893 12207 3927
rect 15485 3893 15519 3927
rect 15853 3893 15887 3927
rect 23397 3893 23431 3927
rect 24777 3893 24811 3927
rect 7481 3689 7515 3723
rect 7849 3689 7883 3723
rect 10609 3689 10643 3723
rect 11345 3689 11379 3723
rect 15025 3689 15059 3723
rect 15485 3689 15519 3723
rect 17417 3689 17451 3723
rect 18521 3689 18555 3723
rect 23673 3689 23707 3723
rect 6377 3621 6411 3655
rect 8217 3621 8251 3655
rect 9045 3621 9079 3655
rect 9942 3621 9976 3655
rect 12218 3621 12252 3655
rect 13829 3621 13863 3655
rect 16037 3621 16071 3655
rect 16589 3621 16623 3655
rect 17922 3621 17956 3655
rect 2881 3553 2915 3587
rect 4512 3553 4546 3587
rect 5492 3553 5526 3587
rect 6469 3553 6503 3587
rect 7021 3553 7055 3587
rect 11897 3553 11931 3587
rect 17601 3553 17635 3587
rect 19349 3553 19383 3587
rect 21557 3553 21591 3587
rect 22477 3553 22511 3587
rect 22753 3553 22787 3587
rect 24041 3553 24075 3587
rect 24133 3553 24167 3587
rect 24317 3553 24351 3587
rect 5595 3485 5629 3519
rect 7205 3485 7239 3519
rect 8125 3485 8159 3519
rect 8769 3485 8803 3519
rect 9689 3485 9723 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 15945 3485 15979 3519
rect 22937 3485 22971 3519
rect 24501 3485 24535 3519
rect 11713 3417 11747 3451
rect 13461 3417 13495 3451
rect 19533 3417 19567 3451
rect 22569 3417 22603 3451
rect 3111 3349 3145 3383
rect 4583 3349 4617 3383
rect 5917 3349 5951 3383
rect 9413 3349 9447 3383
rect 10885 3349 10919 3383
rect 12817 3349 12851 3383
rect 13093 3349 13127 3383
rect 14657 3349 14691 3383
rect 18889 3349 18923 3383
rect 19993 3349 20027 3383
rect 21373 3349 21407 3383
rect 22201 3349 22235 3383
rect 4629 3145 4663 3179
rect 5273 3145 5307 3179
rect 6469 3145 6503 3179
rect 7021 3145 7055 3179
rect 8677 3145 8711 3179
rect 10057 3145 10091 3179
rect 11897 3145 11931 3179
rect 13737 3145 13771 3179
rect 15577 3145 15611 3179
rect 15945 3145 15979 3179
rect 17693 3145 17727 3179
rect 19349 3145 19383 3179
rect 20177 3145 20211 3179
rect 21741 3145 21775 3179
rect 24409 3145 24443 3179
rect 19809 3077 19843 3111
rect 22385 3077 22419 3111
rect 24777 3077 24811 3111
rect 3065 3009 3099 3043
rect 5641 3009 5675 3043
rect 8861 3009 8895 3043
rect 11161 3009 11195 3043
rect 12817 3009 12851 3043
rect 16589 3009 16623 3043
rect 18153 3009 18187 3043
rect 21373 3009 21407 3043
rect 22109 3009 22143 3043
rect 24133 3009 24167 3043
rect 2329 2941 2363 2975
rect 2456 2941 2490 2975
rect 3776 2941 3810 2975
rect 4788 2941 4822 2975
rect 5800 2941 5834 2975
rect 7573 2941 7607 2975
rect 7849 2941 7883 2975
rect 8033 2941 8067 2975
rect 17877 2941 17911 2975
rect 19625 2941 19659 2975
rect 21281 2941 21315 2975
rect 22201 2941 22235 2975
rect 24593 2941 24627 2975
rect 9182 2873 9216 2907
rect 10885 2873 10919 2907
rect 10977 2873 11011 2907
rect 12541 2873 12575 2907
rect 12633 2873 12667 2907
rect 14565 2873 14599 2907
rect 14657 2873 14691 2907
rect 15209 2873 15243 2907
rect 16129 2873 16163 2907
rect 16221 2873 16255 2907
rect 17325 2873 17359 2907
rect 18245 2873 18279 2907
rect 18797 2873 18831 2907
rect 20545 2873 20579 2907
rect 22661 2873 22695 2907
rect 23489 2873 23523 2907
rect 2559 2805 2593 2839
rect 3847 2805 3881 2839
rect 4169 2805 4203 2839
rect 4859 2805 4893 2839
rect 5871 2805 5905 2839
rect 8401 2805 8435 2839
rect 9781 2805 9815 2839
rect 10609 2805 10643 2839
rect 14381 2805 14415 2839
rect 17877 2805 17911 2839
rect 23029 2805 23063 2839
rect 25237 2805 25271 2839
rect 6285 2601 6319 2635
rect 6653 2601 6687 2635
rect 7665 2601 7699 2635
rect 8033 2601 8067 2635
rect 9137 2601 9171 2635
rect 10793 2601 10827 2635
rect 11989 2601 12023 2635
rect 12357 2601 12391 2635
rect 17325 2601 17359 2635
rect 23029 2601 23063 2635
rect 3249 2533 3283 2567
rect 5089 2533 5123 2567
rect 5733 2533 5767 2567
rect 8309 2533 8343 2567
rect 9965 2533 9999 2567
rect 11253 2533 11287 2567
rect 12725 2533 12759 2567
rect 12817 2533 12851 2567
rect 13369 2533 13403 2567
rect 15301 2533 15335 2567
rect 15669 2533 15703 2567
rect 17785 2533 17819 2567
rect 18521 2533 18555 2567
rect 19717 2533 19751 2567
rect 21925 2533 21959 2567
rect 1660 2465 1694 2499
rect 3040 2465 3074 2499
rect 4880 2465 4914 2499
rect 7021 2465 7055 2499
rect 11437 2465 11471 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 17141 2465 17175 2499
rect 19901 2465 19935 2499
rect 21005 2465 21039 2499
rect 21189 2465 21223 2499
rect 21465 2465 21499 2499
rect 22293 2465 22327 2499
rect 22753 2465 22787 2499
rect 3433 2397 3467 2431
rect 5825 2397 5859 2431
rect 8217 2397 8251 2431
rect 9505 2397 9539 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 14105 2397 14139 2431
rect 15577 2397 15611 2431
rect 16037 2397 16071 2431
rect 18153 2397 18187 2431
rect 18429 2397 18463 2431
rect 18705 2397 18739 2431
rect 20637 2397 20671 2431
rect 21281 2397 21315 2431
rect 1731 2329 1765 2363
rect 8769 2329 8803 2363
rect 11621 2329 11655 2363
rect 13737 2329 13771 2363
rect 16865 2329 16899 2363
rect 20085 2329 20119 2363
rect 24777 2533 24811 2567
rect 23213 2465 23247 2499
rect 23857 2465 23891 2499
rect 24133 2465 24167 2499
rect 25672 2465 25706 2499
rect 25743 2329 25777 2363
rect 2053 2261 2087 2295
rect 5365 2261 5399 2295
rect 7205 2261 7239 2295
rect 14381 2261 14415 2295
rect 16497 2261 16531 2295
rect 19349 2261 19383 2295
rect 22937 2261 22971 2295
rect 23029 2261 23063 2295
rect 26157 2261 26191 2295
<< metal1 >>
rect 8294 27480 8300 27532
rect 8352 27520 8358 27532
rect 9030 27520 9036 27532
rect 8352 27492 9036 27520
rect 8352 27480 8358 27492
rect 9030 27480 9036 27492
rect 9088 27480 9094 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 24489 24939 24547 24945
rect 24489 24905 24501 24939
rect 24535 24936 24547 24939
rect 26234 24936 26240 24948
rect 24535 24908 26240 24936
rect 24535 24905 24547 24908
rect 24489 24899 24547 24905
rect 26234 24896 26240 24908
rect 26292 24896 26298 24948
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 12342 24800 12348 24812
rect 6972 24772 12348 24800
rect 6972 24760 6978 24772
rect 12342 24760 12348 24772
rect 12400 24760 12406 24812
rect 23474 24692 23480 24744
rect 23532 24732 23538 24744
rect 24305 24735 24363 24741
rect 24305 24732 24317 24735
rect 23532 24704 24317 24732
rect 23532 24692 23538 24704
rect 24305 24701 24317 24704
rect 24351 24732 24363 24735
rect 24857 24735 24915 24741
rect 24857 24732 24869 24735
rect 24351 24704 24869 24732
rect 24351 24701 24363 24704
rect 24305 24695 24363 24701
rect 24857 24701 24869 24704
rect 24903 24701 24915 24735
rect 24857 24695 24915 24701
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 20898 24392 20904 24404
rect 19935 24364 20904 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 20898 24352 20904 24364
rect 20956 24352 20962 24404
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 27338 24392 27344 24404
rect 24811 24364 27344 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 27338 24352 27344 24364
rect 27396 24352 27402 24404
rect 4706 24216 4712 24268
rect 4764 24256 4770 24268
rect 7412 24259 7470 24265
rect 7412 24256 7424 24259
rect 4764 24228 7424 24256
rect 4764 24216 4770 24228
rect 7412 24225 7424 24228
rect 7458 24256 7470 24259
rect 8110 24256 8116 24268
rect 7458 24228 8116 24256
rect 7458 24225 7470 24228
rect 7412 24219 7470 24225
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 17678 24216 17684 24268
rect 17736 24256 17742 24268
rect 18360 24259 18418 24265
rect 18360 24256 18372 24259
rect 17736 24228 18372 24256
rect 17736 24216 17742 24228
rect 18360 24225 18372 24228
rect 18406 24256 18418 24259
rect 19150 24256 19156 24268
rect 18406 24228 19156 24256
rect 18406 24225 18418 24228
rect 18360 24219 18418 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 19978 24256 19984 24268
rect 19751 24228 19984 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 23106 24256 23112 24268
rect 23067 24228 23112 24256
rect 23106 24216 23112 24228
rect 23164 24216 23170 24268
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 25130 24256 25136 24268
rect 24627 24228 25136 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 23293 24123 23351 24129
rect 23293 24089 23305 24123
rect 23339 24120 23351 24123
rect 24854 24120 24860 24132
rect 23339 24092 24860 24120
rect 23339 24089 23351 24092
rect 23293 24083 23351 24089
rect 24854 24080 24860 24092
rect 24912 24080 24918 24132
rect 7515 24055 7573 24061
rect 7515 24021 7527 24055
rect 7561 24052 7573 24055
rect 8018 24052 8024 24064
rect 7561 24024 8024 24052
rect 7561 24021 7573 24024
rect 7515 24015 7573 24021
rect 8018 24012 8024 24024
rect 8076 24012 8082 24064
rect 18463 24055 18521 24061
rect 18463 24021 18475 24055
rect 18509 24052 18521 24055
rect 18874 24052 18880 24064
rect 18509 24024 18880 24052
rect 18509 24021 18521 24024
rect 18463 24015 18521 24021
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2866 23848 2872 23860
rect 2827 23820 2872 23848
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 3878 23848 3884 23860
rect 3839 23820 3884 23848
rect 3878 23808 3884 23820
rect 3936 23808 3942 23860
rect 8110 23848 8116 23860
rect 8071 23820 8116 23848
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 18417 23851 18475 23857
rect 18417 23817 18429 23851
rect 18463 23848 18475 23851
rect 19518 23848 19524 23860
rect 18463 23820 19524 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 20073 23851 20131 23857
rect 20073 23817 20085 23851
rect 20119 23848 20131 23851
rect 21910 23848 21916 23860
rect 20119 23820 21916 23848
rect 20119 23817 20131 23820
rect 20073 23811 20131 23817
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 24118 23848 24124 23860
rect 22695 23820 24124 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 24118 23808 24124 23820
rect 24176 23808 24182 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 1486 23740 1492 23792
rect 1544 23780 1550 23792
rect 1544 23752 4154 23780
rect 1544 23740 1550 23752
rect 474 23604 480 23656
rect 532 23644 538 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 532 23616 1444 23644
rect 532 23604 538 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 2476 23647 2534 23653
rect 2476 23613 2488 23647
rect 2522 23644 2534 23647
rect 2866 23644 2872 23656
rect 2522 23616 2872 23644
rect 2522 23613 2534 23616
rect 2476 23607 2534 23613
rect 2866 23604 2872 23616
rect 2924 23604 2930 23656
rect 3472 23647 3530 23653
rect 3472 23613 3484 23647
rect 3518 23644 3530 23647
rect 3878 23644 3884 23656
rect 3518 23616 3884 23644
rect 3518 23613 3530 23616
rect 3472 23607 3530 23613
rect 3878 23604 3884 23616
rect 3936 23604 3942 23656
rect 4126 23644 4154 23752
rect 6178 23740 6184 23792
rect 6236 23780 6242 23792
rect 11425 23783 11483 23789
rect 11425 23780 11437 23783
rect 6236 23752 11437 23780
rect 6236 23740 6242 23752
rect 7320 23647 7378 23653
rect 7320 23644 7332 23647
rect 4126 23616 7332 23644
rect 7320 23613 7332 23616
rect 7366 23644 7378 23647
rect 7745 23647 7803 23653
rect 7745 23644 7757 23647
rect 7366 23616 7757 23644
rect 7366 23613 7378 23616
rect 7320 23607 7378 23613
rect 7745 23613 7757 23616
rect 7791 23613 7803 23647
rect 7745 23607 7803 23613
rect 7926 23604 7932 23656
rect 7984 23644 7990 23656
rect 11047 23653 11075 23752
rect 11425 23749 11437 23752
rect 11471 23749 11483 23783
rect 11425 23743 11483 23749
rect 17037 23783 17095 23789
rect 17037 23749 17049 23783
rect 17083 23780 17095 23783
rect 18506 23780 18512 23792
rect 17083 23752 18512 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 18506 23740 18512 23752
rect 18564 23740 18570 23792
rect 19150 23780 19156 23792
rect 19111 23752 19156 23780
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 21177 23783 21235 23789
rect 21177 23749 21189 23783
rect 21223 23780 21235 23783
rect 22738 23780 22744 23792
rect 21223 23752 22744 23780
rect 21223 23749 21235 23752
rect 21177 23743 21235 23749
rect 22738 23740 22744 23752
rect 22796 23740 22802 23792
rect 8332 23647 8390 23653
rect 8332 23644 8344 23647
rect 7984 23616 8344 23644
rect 7984 23604 7990 23616
rect 8332 23613 8344 23616
rect 8378 23644 8390 23647
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 8378 23616 8769 23644
rect 8378 23613 8390 23616
rect 8332 23607 8390 23613
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 8757 23607 8815 23613
rect 11016 23647 11075 23653
rect 11016 23613 11028 23647
rect 11062 23616 11075 23647
rect 11062 23613 11074 23616
rect 11016 23607 11074 23613
rect 12342 23604 12348 23656
rect 12400 23644 12406 23656
rect 12472 23647 12530 23653
rect 12472 23644 12484 23647
rect 12400 23616 12484 23644
rect 12400 23604 12406 23616
rect 12472 23613 12484 23616
rect 12518 23644 12530 23647
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12518 23616 12909 23644
rect 12518 23613 12530 23616
rect 12472 23607 12530 23613
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 12897 23607 12955 23613
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 15620 23616 16865 23644
rect 15620 23604 15626 23616
rect 16853 23613 16865 23616
rect 16899 23613 16911 23647
rect 16853 23607 16911 23613
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 3559 23579 3617 23585
rect 1581 23548 2452 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 2424 23520 2452 23548
rect 3559 23545 3571 23579
rect 3605 23576 3617 23579
rect 6730 23576 6736 23588
rect 3605 23548 6736 23576
rect 3605 23545 3617 23548
rect 3559 23539 3617 23545
rect 6730 23536 6736 23548
rect 6788 23536 6794 23588
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 8435 23579 8493 23585
rect 8435 23576 8447 23579
rect 7892 23548 8447 23576
rect 7892 23536 7898 23548
rect 8435 23545 8447 23548
rect 8481 23545 8493 23579
rect 8435 23539 8493 23545
rect 11103 23579 11161 23585
rect 11103 23545 11115 23579
rect 11149 23576 11161 23579
rect 12066 23576 12072 23588
rect 11149 23548 12072 23576
rect 11149 23545 11161 23548
rect 11103 23539 11161 23545
rect 12066 23536 12072 23548
rect 12124 23536 12130 23588
rect 16868 23576 16896 23607
rect 17310 23604 17316 23656
rect 17368 23644 17374 23656
rect 18233 23647 18291 23653
rect 18233 23644 18245 23647
rect 17368 23616 18245 23644
rect 17368 23604 17374 23616
rect 18233 23613 18245 23616
rect 18279 23644 18291 23647
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 18279 23616 18797 23644
rect 18279 23613 18291 23616
rect 18233 23607 18291 23613
rect 18785 23613 18797 23616
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23613 19947 23647
rect 19889 23607 19947 23613
rect 17405 23579 17463 23585
rect 17405 23576 17417 23579
rect 16868 23548 17417 23576
rect 17405 23545 17417 23548
rect 17451 23545 17463 23579
rect 17405 23539 17463 23545
rect 17494 23536 17500 23588
rect 17552 23576 17558 23588
rect 19904 23576 19932 23607
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 20993 23647 21051 23653
rect 20993 23644 21005 23647
rect 20956 23616 21005 23644
rect 20956 23604 20962 23616
rect 20993 23613 21005 23616
rect 21039 23644 21051 23647
rect 21545 23647 21603 23653
rect 21545 23644 21557 23647
rect 21039 23616 21557 23644
rect 21039 23613 21051 23616
rect 20993 23607 21051 23613
rect 21545 23613 21557 23616
rect 21591 23613 21603 23647
rect 21545 23607 21603 23613
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23613 22523 23647
rect 22465 23607 22523 23613
rect 20441 23579 20499 23585
rect 20441 23576 20453 23579
rect 17552 23548 20453 23576
rect 17552 23536 17558 23548
rect 20441 23545 20453 23548
rect 20487 23545 20499 23579
rect 20441 23539 20499 23545
rect 20806 23536 20812 23588
rect 20864 23576 20870 23588
rect 22480 23576 22508 23607
rect 23017 23579 23075 23585
rect 23017 23576 23029 23579
rect 20864 23548 23029 23576
rect 20864 23536 20870 23548
rect 23017 23545 23029 23548
rect 23063 23545 23075 23579
rect 23017 23539 23075 23545
rect 2406 23468 2412 23520
rect 2464 23468 2470 23520
rect 2547 23511 2605 23517
rect 2547 23477 2559 23511
rect 2593 23508 2605 23511
rect 2682 23508 2688 23520
rect 2593 23480 2688 23508
rect 2593 23477 2605 23480
rect 2547 23471 2605 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 6822 23468 6828 23520
rect 6880 23508 6886 23520
rect 7423 23511 7481 23517
rect 7423 23508 7435 23511
rect 6880 23480 7435 23508
rect 6880 23468 6886 23480
rect 7423 23477 7435 23480
rect 7469 23477 7481 23511
rect 7423 23471 7481 23477
rect 12158 23468 12164 23520
rect 12216 23508 12222 23520
rect 12575 23511 12633 23517
rect 12575 23508 12587 23511
rect 12216 23480 12587 23508
rect 12216 23468 12222 23480
rect 12575 23477 12587 23480
rect 12621 23477 12633 23511
rect 12575 23471 12633 23477
rect 19797 23511 19855 23517
rect 19797 23477 19809 23511
rect 19843 23508 19855 23511
rect 19978 23508 19984 23520
rect 19843 23480 19984 23508
rect 19843 23477 19855 23480
rect 19797 23471 19855 23477
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 23106 23508 23112 23520
rect 20772 23480 23112 23508
rect 20772 23468 20778 23480
rect 23106 23468 23112 23480
rect 23164 23508 23170 23520
rect 23385 23511 23443 23517
rect 23385 23508 23397 23511
rect 23164 23480 23397 23508
rect 23164 23468 23170 23480
rect 23385 23477 23397 23480
rect 23431 23477 23443 23511
rect 23385 23471 23443 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 25590 23168 25596 23180
rect 24627 23140 25596 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 25590 23128 25596 23140
rect 25648 23128 25654 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 25133 22763 25191 22769
rect 25133 22729 25145 22763
rect 25179 22760 25191 22763
rect 25222 22760 25228 22772
rect 25179 22732 25228 22760
rect 25179 22729 25191 22732
rect 25133 22723 25191 22729
rect 24648 22559 24706 22565
rect 24648 22525 24660 22559
rect 24694 22556 24706 22559
rect 25148 22556 25176 22723
rect 25222 22720 25228 22732
rect 25280 22720 25286 22772
rect 24694 22528 25176 22556
rect 24694 22525 24706 22528
rect 24648 22519 24706 22525
rect 24118 22380 24124 22432
rect 24176 22420 24182 22432
rect 24719 22423 24777 22429
rect 24719 22420 24731 22423
rect 24176 22392 24731 22420
rect 24176 22380 24182 22392
rect 24719 22389 24731 22392
rect 24765 22389 24777 22423
rect 24719 22383 24777 22389
rect 25501 22423 25559 22429
rect 25501 22389 25513 22423
rect 25547 22420 25559 22423
rect 25590 22420 25596 22432
rect 25547 22392 25596 22420
rect 25547 22389 25559 22392
rect 25501 22383 25559 22389
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21468 24639 21471
rect 24627 21440 25268 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25240 21341 25268 21440
rect 25225 21335 25283 21341
rect 25225 21301 25237 21335
rect 25271 21332 25283 21335
rect 25498 21332 25504 21344
rect 25271 21304 25504 21332
rect 25271 21301 25283 21304
rect 25225 21295 25283 21301
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 22002 21128 22008 21140
rect 20864 21100 22008 21128
rect 20864 21088 20870 21100
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 11146 21020 11152 21072
rect 11204 21060 11210 21072
rect 14826 21060 14832 21072
rect 11204 21032 14832 21060
rect 11204 21020 11210 21032
rect 14826 21020 14832 21032
rect 14884 21020 14890 21072
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 20936 20995 20994 21001
rect 20936 20992 20948 20995
rect 20864 20964 20948 20992
rect 20864 20952 20870 20964
rect 20936 20961 20948 20964
rect 20982 20961 20994 20995
rect 20936 20955 20994 20961
rect 20162 20748 20168 20800
rect 20220 20788 20226 20800
rect 21039 20791 21097 20797
rect 21039 20788 21051 20791
rect 20220 20760 21051 20788
rect 20220 20748 20226 20760
rect 21039 20757 21051 20760
rect 21085 20757 21097 20791
rect 21039 20751 21097 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 24762 20584 24768 20596
rect 24723 20556 24768 20584
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 19429 20383 19487 20389
rect 19429 20380 19441 20383
rect 19392 20352 19441 20380
rect 19392 20340 19398 20352
rect 19429 20349 19441 20352
rect 19475 20380 19487 20383
rect 19889 20383 19947 20389
rect 19889 20380 19901 20383
rect 19475 20352 19901 20380
rect 19475 20349 19487 20352
rect 19429 20343 19487 20349
rect 19889 20349 19901 20352
rect 19935 20349 19947 20383
rect 24578 20380 24584 20392
rect 24491 20352 24584 20380
rect 19889 20343 19947 20349
rect 24578 20340 24584 20352
rect 24636 20380 24642 20392
rect 25133 20383 25191 20389
rect 25133 20380 25145 20383
rect 24636 20352 25145 20380
rect 24636 20340 24642 20352
rect 25133 20349 25145 20352
rect 25179 20349 25191 20383
rect 25133 20343 25191 20349
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19576 20216 19625 20244
rect 19576 20204 19582 20216
rect 19613 20213 19625 20216
rect 19659 20213 19671 20247
rect 20438 20244 20444 20256
rect 20399 20216 20444 20244
rect 19613 20207 19671 20213
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 20806 20204 20812 20256
rect 20864 20244 20870 20256
rect 20901 20247 20959 20253
rect 20901 20244 20913 20247
rect 20864 20216 20913 20244
rect 20864 20204 20870 20216
rect 20901 20213 20913 20216
rect 20947 20213 20959 20247
rect 20901 20207 20959 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 13354 20040 13360 20052
rect 12584 20012 13360 20040
rect 12584 20000 12590 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19981 20043 20039 20049
rect 19981 20040 19993 20043
rect 18932 20012 19993 20040
rect 18932 20000 18938 20012
rect 19981 20009 19993 20012
rect 20027 20040 20039 20043
rect 20070 20040 20076 20052
rect 20027 20012 20076 20040
rect 20027 20009 20039 20012
rect 19981 20003 20039 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 23707 20043 23765 20049
rect 23707 20009 23719 20043
rect 23753 20040 23765 20043
rect 24578 20040 24584 20052
rect 23753 20012 24584 20040
rect 23753 20009 23765 20012
rect 23707 20003 23765 20009
rect 24578 20000 24584 20012
rect 24636 20000 24642 20052
rect 15930 19864 15936 19916
rect 15988 19904 15994 19916
rect 16060 19907 16118 19913
rect 16060 19904 16072 19907
rect 15988 19876 16072 19904
rect 15988 19864 15994 19876
rect 16060 19873 16072 19876
rect 16106 19873 16118 19907
rect 20990 19904 20996 19916
rect 20951 19876 20996 19904
rect 16060 19867 16118 19873
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 22554 19913 22560 19916
rect 22500 19907 22560 19913
rect 22500 19904 22512 19907
rect 21237 19876 22512 19904
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19058 19836 19064 19848
rect 18923 19808 19064 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19978 19796 19984 19848
rect 20036 19836 20042 19848
rect 21237 19836 21265 19876
rect 22500 19873 22512 19876
rect 22546 19873 22560 19907
rect 22500 19867 22560 19873
rect 22554 19864 22560 19867
rect 22612 19864 22618 19916
rect 23636 19907 23694 19913
rect 23636 19873 23648 19907
rect 23682 19904 23694 19907
rect 23842 19904 23848 19916
rect 23682 19876 23848 19904
rect 23682 19873 23694 19876
rect 23636 19867 23694 19873
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 20036 19808 21265 19836
rect 20036 19796 20042 19808
rect 16163 19703 16221 19709
rect 16163 19669 16175 19703
rect 16209 19700 16221 19703
rect 16298 19700 16304 19712
rect 16209 19672 16304 19700
rect 16209 19669 16221 19672
rect 16163 19663 16221 19669
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 19107 19703 19165 19709
rect 19107 19669 19119 19703
rect 19153 19700 19165 19703
rect 19242 19700 19248 19712
rect 19153 19672 19248 19700
rect 19153 19669 19165 19672
rect 19107 19663 19165 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 21174 19700 21180 19712
rect 21135 19672 21180 19700
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 22462 19660 22468 19712
rect 22520 19700 22526 19712
rect 22603 19703 22661 19709
rect 22603 19700 22615 19703
rect 22520 19672 22615 19700
rect 22520 19660 22526 19672
rect 22603 19669 22615 19672
rect 22649 19669 22661 19703
rect 22603 19663 22661 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 16942 19496 16948 19508
rect 16903 19468 16948 19496
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 19058 19456 19064 19508
rect 19116 19496 19122 19508
rect 19337 19499 19395 19505
rect 19337 19496 19349 19499
rect 19116 19468 19349 19496
rect 19116 19456 19122 19468
rect 19337 19465 19349 19468
rect 19383 19465 19395 19499
rect 22554 19496 22560 19508
rect 22515 19468 22560 19496
rect 19337 19459 19395 19465
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 24762 19496 24768 19508
rect 24723 19468 24768 19496
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 16022 19388 16028 19440
rect 16080 19428 16086 19440
rect 16669 19431 16727 19437
rect 16669 19428 16681 19431
rect 16080 19400 16681 19428
rect 16080 19388 16086 19400
rect 16669 19397 16681 19400
rect 16715 19428 16727 19431
rect 17494 19428 17500 19440
rect 16715 19400 17500 19428
rect 16715 19397 16727 19400
rect 16669 19391 16727 19397
rect 17494 19388 17500 19400
rect 17552 19388 17558 19440
rect 20070 19360 20076 19372
rect 20031 19332 20076 19360
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 20990 19360 20996 19372
rect 20312 19332 20996 19360
rect 20312 19320 20318 19332
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 16184 19295 16242 19301
rect 16184 19261 16196 19295
rect 16230 19292 16242 19295
rect 16942 19292 16948 19304
rect 16230 19264 16948 19292
rect 16230 19261 16242 19264
rect 16184 19255 16242 19261
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 21453 19295 21511 19301
rect 21453 19261 21465 19295
rect 21499 19292 21511 19295
rect 21634 19292 21640 19304
rect 21499 19264 21640 19292
rect 21499 19261 21511 19264
rect 21453 19255 21511 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 24581 19295 24639 19301
rect 24581 19261 24593 19295
rect 24627 19292 24639 19295
rect 24854 19292 24860 19304
rect 24627 19264 24860 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 24854 19252 24860 19264
rect 24912 19292 24918 19304
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24912 19264 25145 19292
rect 24912 19252 24918 19264
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 20165 19227 20223 19233
rect 20165 19193 20177 19227
rect 20211 19193 20223 19227
rect 20714 19224 20720 19236
rect 20675 19196 20720 19224
rect 20165 19187 20223 19193
rect 16255 19159 16313 19165
rect 16255 19125 16267 19159
rect 16301 19156 16313 19159
rect 16482 19156 16488 19168
rect 16301 19128 16488 19156
rect 16301 19125 16313 19128
rect 16255 19119 16313 19125
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 18598 19156 18604 19168
rect 18559 19128 18604 19156
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20180 19156 20208 19187
rect 20714 19184 20720 19196
rect 20772 19184 20778 19236
rect 21174 19224 21180 19236
rect 20916 19196 21180 19224
rect 20916 19156 20944 19196
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 21542 19224 21548 19236
rect 21503 19196 21548 19224
rect 21542 19184 21548 19196
rect 21600 19184 21606 19236
rect 23842 19156 23848 19168
rect 19935 19128 20944 19156
rect 23803 19128 23848 19156
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 23842 19116 23848 19128
rect 23900 19116 23906 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 19153 18955 19211 18961
rect 19153 18921 19165 18955
rect 19199 18952 19211 18955
rect 19242 18952 19248 18964
rect 19199 18924 19248 18952
rect 19199 18921 19211 18924
rect 19153 18915 19211 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 17126 18884 17132 18896
rect 16540 18856 17132 18884
rect 16540 18844 16546 18856
rect 17126 18844 17132 18856
rect 17184 18844 17190 18896
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 17402 18884 17408 18896
rect 17267 18856 17408 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 19260 18884 19288 18912
rect 19337 18887 19395 18893
rect 19337 18884 19349 18887
rect 19260 18856 19349 18884
rect 19337 18853 19349 18856
rect 19383 18853 19395 18887
rect 19337 18847 19395 18853
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 19484 18856 19529 18884
rect 19484 18844 19490 18856
rect 20438 18844 20444 18896
rect 20496 18884 20502 18896
rect 20990 18884 20996 18896
rect 20496 18856 20996 18884
rect 20496 18844 20502 18856
rect 20990 18844 20996 18856
rect 21048 18844 21054 18896
rect 21085 18887 21143 18893
rect 21085 18853 21097 18887
rect 21131 18884 21143 18887
rect 21174 18884 21180 18896
rect 21131 18856 21180 18884
rect 21131 18853 21143 18856
rect 21085 18847 21143 18853
rect 21174 18844 21180 18856
rect 21232 18844 21238 18896
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18816 16083 18819
rect 16114 18816 16120 18828
rect 16071 18788 16120 18816
rect 16071 18785 16083 18788
rect 16025 18779 16083 18785
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23236 18819 23294 18825
rect 23236 18816 23248 18819
rect 23072 18788 23248 18816
rect 23072 18776 23078 18788
rect 23236 18785 23248 18788
rect 23282 18785 23294 18819
rect 23236 18779 23294 18785
rect 24280 18819 24338 18825
rect 24280 18785 24292 18819
rect 24326 18816 24338 18819
rect 24762 18816 24768 18828
rect 24326 18788 24768 18816
rect 24326 18785 24338 18788
rect 24280 18779 24338 18785
rect 24762 18776 24768 18788
rect 24820 18776 24826 18828
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 17276 18720 17417 18748
rect 17276 18708 17282 18720
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20714 18748 20720 18760
rect 20027 18720 20720 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21450 18748 21456 18760
rect 21411 18720 21456 18748
rect 21450 18708 21456 18720
rect 21508 18748 21514 18760
rect 21913 18751 21971 18757
rect 21913 18748 21925 18751
rect 21508 18720 21925 18748
rect 21508 18708 21514 18720
rect 21913 18717 21925 18720
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 16163 18615 16221 18621
rect 16163 18581 16175 18615
rect 16209 18612 16221 18615
rect 18138 18612 18144 18624
rect 16209 18584 18144 18612
rect 16209 18581 16221 18584
rect 16163 18575 16221 18581
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 18414 18612 18420 18624
rect 18375 18584 18420 18612
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 23339 18615 23397 18621
rect 23339 18581 23351 18615
rect 23385 18612 23397 18615
rect 24210 18612 24216 18624
rect 23385 18584 24216 18612
rect 23385 18581 23397 18584
rect 23339 18575 23397 18581
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 24351 18615 24409 18621
rect 24351 18581 24363 18615
rect 24397 18612 24409 18615
rect 24670 18612 24676 18624
rect 24397 18584 24676 18612
rect 24397 18581 24409 18584
rect 24351 18575 24409 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 21174 18408 21180 18420
rect 21135 18380 21180 18408
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 21542 18408 21548 18420
rect 21503 18380 21548 18408
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 25406 18408 25412 18420
rect 25367 18380 25412 18408
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 13538 18340 13544 18352
rect 9732 18312 13544 18340
rect 9732 18300 9738 18312
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 12802 18232 12808 18284
rect 12860 18272 12866 18284
rect 16114 18272 16120 18284
rect 12860 18244 16120 18272
rect 12860 18232 12866 18244
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 18138 18272 18144 18284
rect 18099 18244 18144 18272
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 18506 18272 18512 18284
rect 18467 18244 18512 18272
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 20162 18272 20168 18284
rect 20123 18244 20168 18272
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18272 20867 18275
rect 21450 18272 21456 18284
rect 20855 18244 21456 18272
rect 20855 18241 20867 18244
rect 20809 18235 20867 18241
rect 21450 18232 21456 18244
rect 21508 18272 21514 18284
rect 21729 18275 21787 18281
rect 21729 18272 21741 18275
rect 21508 18244 21741 18272
rect 21508 18232 21514 18244
rect 21729 18241 21741 18244
rect 21775 18241 21787 18275
rect 22186 18272 22192 18284
rect 22147 18244 22192 18272
rect 21729 18235 21787 18241
rect 22186 18232 22192 18244
rect 22244 18272 22250 18284
rect 23014 18272 23020 18284
rect 22244 18244 23020 18272
rect 22244 18232 22250 18244
rect 23014 18232 23020 18244
rect 23072 18232 23078 18284
rect 23446 18244 24025 18272
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 14458 18213 14464 18216
rect 12472 18207 12530 18213
rect 12472 18204 12484 18207
rect 12308 18176 12484 18204
rect 12308 18164 12314 18176
rect 12472 18173 12484 18176
rect 12518 18204 12530 18207
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12518 18176 12909 18204
rect 12518 18173 12530 18176
rect 12472 18167 12530 18173
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 14436 18207 14464 18213
rect 14436 18204 14448 18207
rect 14371 18176 14448 18204
rect 12897 18167 12955 18173
rect 14436 18173 14448 18176
rect 14516 18204 14522 18216
rect 14829 18207 14887 18213
rect 14829 18204 14841 18207
rect 14516 18176 14841 18204
rect 14436 18167 14464 18173
rect 14458 18164 14464 18167
rect 14516 18164 14522 18176
rect 14829 18173 14841 18176
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 15416 18207 15474 18213
rect 15416 18173 15428 18207
rect 15462 18173 15474 18207
rect 15416 18167 15474 18173
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18204 17095 18207
rect 17083 18176 17908 18204
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 12575 18139 12633 18145
rect 12575 18105 12587 18139
rect 12621 18136 12633 18139
rect 12621 18108 13486 18136
rect 12621 18105 12633 18108
rect 12575 18099 12633 18105
rect 13458 18068 13486 18108
rect 13538 18096 13544 18148
rect 13596 18136 13602 18148
rect 15197 18139 15255 18145
rect 15197 18136 15209 18139
rect 13596 18108 15209 18136
rect 13596 18096 13602 18108
rect 15197 18105 15209 18108
rect 15243 18136 15255 18139
rect 15431 18136 15459 18167
rect 15243 18108 15459 18136
rect 17129 18139 17187 18145
rect 15243 18105 15255 18108
rect 15197 18099 15255 18105
rect 17129 18105 17141 18139
rect 17175 18105 17187 18139
rect 17129 18099 17187 18105
rect 14366 18068 14372 18080
rect 13458 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14507 18071 14565 18077
rect 14507 18037 14519 18071
rect 14553 18068 14565 18071
rect 15378 18068 15384 18080
rect 14553 18040 15384 18068
rect 14553 18037 14565 18040
rect 14507 18031 14565 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15519 18071 15577 18077
rect 15519 18037 15531 18071
rect 15565 18068 15577 18071
rect 15838 18068 15844 18080
rect 15565 18040 15844 18068
rect 15565 18037 15577 18040
rect 15519 18031 15577 18037
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 17144 18068 17172 18099
rect 17402 18068 17408 18080
rect 17144 18040 17408 18068
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17880 18077 17908 18176
rect 18233 18139 18291 18145
rect 18233 18105 18245 18139
rect 18279 18105 18291 18139
rect 18233 18099 18291 18105
rect 19337 18139 19395 18145
rect 19337 18105 19349 18139
rect 19383 18136 19395 18139
rect 19426 18136 19432 18148
rect 19383 18108 19432 18136
rect 19383 18105 19395 18108
rect 19337 18099 19395 18105
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 17954 18068 17960 18080
rect 17911 18040 17960 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 17954 18028 17960 18040
rect 18012 18068 18018 18080
rect 18248 18068 18276 18099
rect 19426 18096 19432 18108
rect 19484 18136 19490 18148
rect 19981 18139 20039 18145
rect 19981 18136 19993 18139
rect 19484 18108 19993 18136
rect 19484 18096 19490 18108
rect 19981 18105 19993 18108
rect 20027 18136 20039 18139
rect 20254 18136 20260 18148
rect 20027 18108 20260 18136
rect 20027 18105 20039 18108
rect 19981 18099 20039 18105
rect 20254 18096 20260 18108
rect 20312 18096 20318 18148
rect 21821 18139 21879 18145
rect 21821 18105 21833 18139
rect 21867 18105 21879 18139
rect 21821 18099 21879 18105
rect 18012 18040 18276 18068
rect 18012 18028 18018 18040
rect 21542 18028 21548 18080
rect 21600 18068 21606 18080
rect 21836 18068 21864 18099
rect 23106 18096 23112 18148
rect 23164 18136 23170 18148
rect 23446 18136 23474 18244
rect 23845 18207 23903 18213
rect 23845 18173 23857 18207
rect 23891 18173 23903 18207
rect 23845 18167 23903 18173
rect 23164 18108 23474 18136
rect 23164 18096 23170 18108
rect 21600 18040 21864 18068
rect 23477 18071 23535 18077
rect 21600 18028 21606 18040
rect 23477 18037 23489 18071
rect 23523 18068 23535 18071
rect 23860 18068 23888 18167
rect 23997 18136 24025 18244
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 24268 18176 25237 18204
rect 24268 18164 24274 18176
rect 25225 18173 25237 18176
rect 25271 18204 25283 18207
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25271 18176 25789 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 24397 18139 24455 18145
rect 24397 18136 24409 18139
rect 23997 18108 24409 18136
rect 24397 18105 24409 18108
rect 24443 18136 24455 18139
rect 25130 18136 25136 18148
rect 24443 18108 25136 18136
rect 24443 18105 24455 18108
rect 24397 18099 24455 18105
rect 25130 18096 25136 18108
rect 25188 18096 25194 18148
rect 24026 18068 24032 18080
rect 23523 18040 24032 18068
rect 23523 18037 23535 18040
rect 23477 18031 23535 18037
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 24578 18028 24584 18080
rect 24636 18068 24642 18080
rect 24673 18071 24731 18077
rect 24673 18068 24685 18071
rect 24636 18040 24685 18068
rect 24636 18028 24642 18040
rect 24673 18037 24685 18040
rect 24719 18068 24731 18071
rect 24762 18068 24768 18080
rect 24719 18040 24768 18068
rect 24719 18037 24731 18040
rect 24673 18031 24731 18037
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17184 17836 17877 17864
rect 17184 17824 17190 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 18233 17867 18291 17873
rect 18233 17864 18245 17867
rect 18196 17836 18245 17864
rect 18196 17824 18202 17836
rect 18233 17833 18245 17836
rect 18279 17833 18291 17867
rect 20162 17864 20168 17876
rect 20123 17836 20168 17864
rect 18233 17827 18291 17833
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20990 17824 20996 17876
rect 21048 17864 21054 17876
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 21048 17836 21097 17864
rect 21048 17824 21054 17836
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 24118 17864 24124 17876
rect 24079 17836 24124 17864
rect 21085 17827 21143 17833
rect 24118 17824 24124 17836
rect 24176 17824 24182 17876
rect 24765 17867 24823 17873
rect 24765 17833 24777 17867
rect 24811 17864 24823 17867
rect 27522 17864 27528 17876
rect 24811 17836 27528 17864
rect 24811 17833 24823 17836
rect 24765 17827 24823 17833
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 13078 17796 13084 17808
rect 13039 17768 13084 17796
rect 13078 17756 13084 17768
rect 13136 17756 13142 17808
rect 13170 17756 13176 17808
rect 13228 17796 13234 17808
rect 17037 17799 17095 17805
rect 13228 17768 13273 17796
rect 13228 17756 13234 17768
rect 17037 17765 17049 17799
rect 17083 17796 17095 17799
rect 17402 17796 17408 17808
rect 17083 17768 17408 17796
rect 17083 17765 17095 17768
rect 17037 17759 17095 17765
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 18598 17796 18604 17808
rect 18559 17768 18604 17796
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 21634 17796 21640 17808
rect 21595 17768 21640 17796
rect 21634 17756 21640 17768
rect 21692 17756 21698 17808
rect 22186 17796 22192 17808
rect 22147 17768 22192 17796
rect 22186 17756 22192 17768
rect 22244 17756 22250 17808
rect 23106 17756 23112 17808
rect 23164 17796 23170 17808
rect 23201 17799 23259 17805
rect 23201 17796 23213 17799
rect 23164 17768 23213 17796
rect 23164 17756 23170 17768
rect 23201 17765 23213 17768
rect 23247 17765 23259 17799
rect 23201 17759 23259 17765
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 9122 17728 9128 17740
rect 8352 17700 9128 17728
rect 8352 17688 8358 17700
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 19150 17688 19156 17740
rect 19208 17728 19214 17740
rect 24581 17731 24639 17737
rect 19208 17700 19253 17728
rect 19208 17688 19214 17700
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17660 15899 17663
rect 16942 17660 16948 17672
rect 15887 17632 16948 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17660 17647 17663
rect 18506 17660 18512 17672
rect 17635 17632 18512 17660
rect 17635 17629 17647 17632
rect 17589 17623 17647 17629
rect 18506 17620 18512 17632
rect 18564 17660 18570 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 18564 17632 19809 17660
rect 18564 17620 18570 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 20714 17620 20720 17672
rect 20772 17660 20778 17672
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 20772 17632 21557 17660
rect 20772 17620 20778 17632
rect 21545 17629 21557 17632
rect 21591 17660 21603 17663
rect 22186 17660 22192 17672
rect 21591 17632 22192 17660
rect 21591 17629 21603 17632
rect 21545 17623 21603 17629
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23566 17660 23572 17672
rect 23527 17632 23572 17660
rect 23109 17623 23167 17629
rect 13630 17592 13636 17604
rect 13591 17564 13636 17592
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 14366 17552 14372 17604
rect 14424 17592 14430 17604
rect 23124 17592 23152 17623
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 23382 17592 23388 17604
rect 14424 17564 23388 17592
rect 14424 17552 14430 17564
rect 23382 17552 23388 17564
rect 23440 17552 23446 17604
rect 16482 17524 16488 17536
rect 16443 17496 16488 17524
rect 16482 17484 16488 17496
rect 16540 17484 16546 17536
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 19429 17527 19487 17533
rect 19429 17524 19441 17527
rect 18564 17496 19441 17524
rect 18564 17484 18570 17496
rect 19429 17493 19441 17496
rect 19475 17493 19487 17527
rect 19429 17487 19487 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 14001 17323 14059 17329
rect 14001 17320 14013 17323
rect 13136 17292 14013 17320
rect 13136 17280 13142 17292
rect 14001 17289 14013 17292
rect 14047 17289 14059 17323
rect 14001 17283 14059 17289
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 15657 17323 15715 17329
rect 15657 17320 15669 17323
rect 15620 17292 15669 17320
rect 15620 17280 15626 17292
rect 15657 17289 15669 17292
rect 15703 17289 15715 17323
rect 15838 17320 15844 17332
rect 15799 17292 15844 17320
rect 15657 17283 15715 17289
rect 15838 17280 15844 17292
rect 15896 17320 15902 17332
rect 17402 17320 17408 17332
rect 15896 17292 16528 17320
rect 17363 17292 17408 17320
rect 15896 17280 15902 17292
rect 12897 17255 12955 17261
rect 12897 17221 12909 17255
rect 12943 17252 12955 17255
rect 13170 17252 13176 17264
rect 12943 17224 13176 17252
rect 12943 17221 12955 17224
rect 12897 17215 12955 17221
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 13630 17252 13636 17264
rect 13591 17224 13636 17252
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 16500 17193 16528 17292
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 18325 17323 18383 17329
rect 18325 17289 18337 17323
rect 18371 17320 18383 17323
rect 18598 17320 18604 17332
rect 18371 17292 18604 17320
rect 18371 17289 18383 17292
rect 18325 17283 18383 17289
rect 18598 17280 18604 17292
rect 18656 17280 18662 17332
rect 21634 17280 21640 17332
rect 21692 17320 21698 17332
rect 21821 17323 21879 17329
rect 21821 17320 21833 17323
rect 21692 17292 21833 17320
rect 21692 17280 21698 17292
rect 21821 17289 21833 17292
rect 21867 17320 21879 17323
rect 22097 17323 22155 17329
rect 22097 17320 22109 17323
rect 21867 17292 22109 17320
rect 21867 17289 21879 17292
rect 21821 17283 21879 17289
rect 22097 17289 22109 17292
rect 22143 17289 22155 17323
rect 22097 17283 22155 17289
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 22465 17323 22523 17329
rect 22465 17320 22477 17323
rect 22244 17292 22477 17320
rect 22244 17280 22250 17292
rect 22465 17289 22477 17292
rect 22511 17289 22523 17323
rect 23106 17320 23112 17332
rect 23067 17292 23112 17320
rect 22465 17283 22523 17289
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23382 17320 23388 17332
rect 23343 17292 23388 17320
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 24949 17323 25007 17329
rect 24949 17320 24961 17323
rect 24728 17292 24961 17320
rect 24728 17280 24734 17292
rect 24949 17289 24961 17292
rect 24995 17289 25007 17323
rect 24949 17283 25007 17289
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12216 17156 13093 17184
rect 12216 17144 12222 17156
rect 13081 17153 13093 17156
rect 13127 17184 13139 17187
rect 14369 17187 14427 17193
rect 14369 17184 14381 17187
rect 13127 17156 14381 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 14369 17153 14381 17156
rect 14415 17153 14427 17187
rect 14369 17147 14427 17153
rect 16485 17187 16543 17193
rect 16485 17153 16497 17187
rect 16531 17153 16543 17187
rect 16485 17147 16543 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17218 17184 17224 17196
rect 17175 17156 17224 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17218 17144 17224 17156
rect 17276 17184 17282 17196
rect 18506 17184 18512 17196
rect 17276 17156 18512 17184
rect 17276 17144 17282 17156
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 19150 17184 19156 17196
rect 19111 17156 19156 17184
rect 19150 17144 19156 17156
rect 19208 17144 19214 17196
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 19300 17156 20729 17184
rect 19300 17144 19306 17156
rect 20717 17153 20729 17156
rect 20763 17184 20775 17187
rect 24029 17187 24087 17193
rect 20763 17156 21312 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 15448 17119 15506 17125
rect 15448 17116 15460 17119
rect 15335 17088 15460 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 15448 17085 15460 17088
rect 15494 17116 15506 17119
rect 15930 17116 15936 17128
rect 15494 17088 15936 17116
rect 15494 17085 15506 17088
rect 15448 17079 15506 17085
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 20487 17088 20913 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 20901 17085 20913 17088
rect 20947 17116 20959 17119
rect 20990 17116 20996 17128
rect 20947 17088 20996 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 21284 17060 21312 17156
rect 24029 17153 24041 17187
rect 24075 17184 24087 17187
rect 24118 17184 24124 17196
rect 24075 17156 24124 17184
rect 24075 17153 24087 17156
rect 24029 17147 24087 17153
rect 24118 17144 24124 17156
rect 24176 17144 24182 17196
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 13173 17051 13231 17057
rect 12299 17020 13032 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 13004 16980 13032 17020
rect 13173 17017 13185 17051
rect 13219 17017 13231 17051
rect 13173 17011 13231 17017
rect 16301 17051 16359 17057
rect 16301 17017 16313 17051
rect 16347 17048 16359 17051
rect 16482 17048 16488 17060
rect 16347 17020 16488 17048
rect 16347 17017 16359 17020
rect 16301 17011 16359 17017
rect 13188 16980 13216 17011
rect 16482 17008 16488 17020
rect 16540 17048 16546 17060
rect 16577 17051 16635 17057
rect 16577 17048 16589 17051
rect 16540 17020 16589 17048
rect 16540 17008 16546 17020
rect 16577 17017 16589 17020
rect 16623 17048 16635 17051
rect 17954 17048 17960 17060
rect 16623 17020 17960 17048
rect 16623 17017 16635 17020
rect 16577 17011 16635 17017
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 18598 17048 18604 17060
rect 18559 17020 18604 17048
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 19521 17051 19579 17057
rect 19521 17017 19533 17051
rect 19567 17048 19579 17051
rect 20530 17048 20536 17060
rect 19567 17020 20536 17048
rect 19567 17017 19579 17020
rect 19521 17011 19579 17017
rect 20530 17008 20536 17020
rect 20588 17008 20594 17060
rect 21266 17057 21272 17060
rect 21263 17011 21272 17057
rect 21324 17048 21330 17060
rect 21324 17020 21417 17048
rect 21266 17008 21272 17011
rect 21324 17008 21330 17020
rect 23014 17008 23020 17060
rect 23072 17048 23078 17060
rect 24026 17048 24032 17060
rect 23072 17020 24032 17048
rect 23072 17008 23078 17020
rect 24026 17008 24032 17020
rect 24084 17048 24090 17060
rect 24121 17051 24179 17057
rect 24121 17048 24133 17051
rect 24084 17020 24133 17048
rect 24084 17008 24090 17020
rect 24121 17017 24133 17020
rect 24167 17017 24179 17051
rect 24121 17011 24179 17017
rect 24673 17051 24731 17057
rect 24673 17017 24685 17051
rect 24719 17048 24731 17051
rect 24762 17048 24768 17060
rect 24719 17020 24768 17048
rect 24719 17017 24731 17020
rect 24673 17011 24731 17017
rect 24762 17008 24768 17020
rect 24820 17008 24826 17060
rect 14734 16980 14740 16992
rect 13004 16952 14740 16980
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18414 16980 18420 16992
rect 17911 16952 18420 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18414 16940 18420 16952
rect 18472 16980 18478 16992
rect 18616 16980 18644 17008
rect 18472 16952 18644 16980
rect 19889 16983 19947 16989
rect 18472 16940 18478 16952
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20162 16980 20168 16992
rect 19935 16952 20168 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 24486 16940 24492 16992
rect 24544 16980 24550 16992
rect 25501 16983 25559 16989
rect 25501 16980 25513 16983
rect 24544 16952 25513 16980
rect 24544 16940 24550 16952
rect 25501 16949 25513 16952
rect 25547 16949 25559 16983
rect 25501 16943 25559 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 11146 16776 11152 16788
rect 11107 16748 11152 16776
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 16942 16776 16948 16788
rect 16903 16748 16948 16776
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 17954 16776 17960 16788
rect 17915 16748 17960 16776
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 19705 16779 19763 16785
rect 19705 16776 19717 16779
rect 18656 16748 19717 16776
rect 18656 16736 18662 16748
rect 19705 16745 19717 16748
rect 19751 16745 19763 16779
rect 19705 16739 19763 16745
rect 20254 16736 20260 16788
rect 20312 16776 20318 16788
rect 21821 16779 21879 16785
rect 21821 16776 21833 16779
rect 20312 16748 21833 16776
rect 20312 16736 20318 16748
rect 21821 16745 21833 16748
rect 21867 16745 21879 16779
rect 21821 16739 21879 16745
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22189 16779 22247 16785
rect 22189 16776 22201 16779
rect 22152 16748 22201 16776
rect 22152 16736 22158 16748
rect 22189 16745 22201 16748
rect 22235 16776 22247 16779
rect 24026 16776 24032 16788
rect 22235 16748 23474 16776
rect 23987 16748 24032 16776
rect 22235 16745 22247 16748
rect 22189 16739 22247 16745
rect 6822 16668 6828 16720
rect 6880 16708 6886 16720
rect 8110 16708 8116 16720
rect 6880 16680 8116 16708
rect 6880 16668 6886 16680
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 8202 16668 8208 16720
rect 8260 16708 8266 16720
rect 13170 16708 13176 16720
rect 8260 16680 8305 16708
rect 13131 16680 13176 16708
rect 8260 16668 8266 16680
rect 13170 16668 13176 16680
rect 13228 16668 13234 16720
rect 17399 16711 17457 16717
rect 17399 16677 17411 16711
rect 17445 16708 17457 16711
rect 17770 16708 17776 16720
rect 17445 16680 17776 16708
rect 17445 16677 17457 16680
rect 17399 16671 17457 16677
rect 17770 16668 17776 16680
rect 17828 16708 17834 16720
rect 19150 16717 19156 16720
rect 19106 16711 19156 16717
rect 19106 16708 19118 16711
rect 17828 16680 19118 16708
rect 17828 16668 17834 16680
rect 19106 16677 19118 16680
rect 19152 16677 19156 16711
rect 19106 16671 19156 16677
rect 19150 16668 19156 16671
rect 19208 16668 19214 16720
rect 19518 16668 19524 16720
rect 19576 16708 19582 16720
rect 19978 16708 19984 16720
rect 19576 16680 19984 16708
rect 19576 16668 19582 16680
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 21147 16711 21205 16717
rect 21147 16677 21159 16711
rect 21193 16708 21205 16711
rect 21266 16708 21272 16720
rect 21193 16680 21272 16708
rect 21193 16677 21205 16680
rect 21147 16671 21205 16677
rect 21266 16668 21272 16680
rect 21324 16668 21330 16720
rect 23014 16708 23020 16720
rect 22975 16680 23020 16708
rect 23014 16668 23020 16680
rect 23072 16668 23078 16720
rect 23446 16708 23474 16748
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 23566 16708 23572 16720
rect 23446 16680 23572 16708
rect 23566 16668 23572 16680
rect 23624 16668 23630 16720
rect 24486 16708 24492 16720
rect 24447 16680 24492 16708
rect 24486 16668 24492 16680
rect 24544 16668 24550 16720
rect 24581 16711 24639 16717
rect 24581 16677 24593 16711
rect 24627 16708 24639 16711
rect 25130 16708 25136 16720
rect 24627 16680 25136 16708
rect 24627 16677 24639 16680
rect 24581 16671 24639 16677
rect 25130 16668 25136 16680
rect 25188 16668 25194 16720
rect 11330 16640 11336 16652
rect 11291 16612 11336 16640
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16640 11667 16643
rect 11790 16640 11796 16652
rect 11655 16612 11796 16640
rect 11655 16609 11667 16612
rect 11609 16603 11667 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 16114 16640 16120 16652
rect 16075 16612 16120 16640
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 8754 16572 8760 16584
rect 8715 16544 8760 16572
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 16206 16572 16212 16584
rect 16167 16544 16212 16572
rect 13081 16535 13139 16541
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 13096 16504 13124 16535
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16572 17095 16575
rect 17494 16572 17500 16584
rect 17083 16544 17500 16572
rect 17083 16541 17095 16544
rect 17037 16535 17095 16541
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 18785 16575 18843 16581
rect 18785 16572 18797 16575
rect 18656 16544 18797 16572
rect 18656 16532 18662 16544
rect 18785 16541 18797 16544
rect 18831 16541 18843 16575
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 18785 16535 18843 16541
rect 20732 16544 20913 16572
rect 13446 16504 13452 16516
rect 6788 16476 13452 16504
rect 6788 16464 6794 16476
rect 13446 16464 13452 16476
rect 13504 16464 13510 16516
rect 13630 16504 13636 16516
rect 13591 16476 13636 16504
rect 13630 16464 13636 16476
rect 13688 16504 13694 16516
rect 15562 16504 15568 16516
rect 13688 16476 15568 16504
rect 13688 16464 13694 16476
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 20732 16448 20760 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 22186 16532 22192 16584
rect 22244 16572 22250 16584
rect 22925 16575 22983 16581
rect 22925 16572 22937 16575
rect 22244 16544 22937 16572
rect 22244 16532 22250 16544
rect 22925 16541 22937 16544
rect 22971 16541 22983 16575
rect 24762 16572 24768 16584
rect 24723 16544 24768 16572
rect 22925 16535 22983 16541
rect 24762 16532 24768 16544
rect 24820 16532 24826 16584
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 9861 16439 9919 16445
rect 9861 16436 9873 16439
rect 9824 16408 9873 16436
rect 9824 16396 9830 16408
rect 9861 16405 9873 16408
rect 9907 16405 9919 16439
rect 13998 16436 14004 16448
rect 13959 16408 14004 16436
rect 9861 16399 9919 16405
rect 13998 16396 14004 16408
rect 14056 16396 14062 16448
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18233 16439 18291 16445
rect 18233 16436 18245 16439
rect 18196 16408 18245 16436
rect 18196 16396 18202 16408
rect 18233 16405 18245 16408
rect 18279 16405 18291 16439
rect 18690 16436 18696 16448
rect 18651 16408 18696 16436
rect 18233 16399 18291 16405
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 20714 16436 20720 16448
rect 20675 16408 20720 16436
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 8168 16204 8953 16232
rect 8168 16192 8174 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13320 16204 13737 16232
rect 13320 16192 13326 16204
rect 13725 16201 13737 16204
rect 13771 16232 13783 16235
rect 14090 16232 14096 16244
rect 13771 16204 14096 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 18463 16235 18521 16241
rect 18463 16201 18475 16235
rect 18509 16232 18521 16235
rect 22186 16232 22192 16244
rect 18509 16204 22192 16232
rect 18509 16201 18521 16204
rect 18463 16195 18521 16201
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 23014 16232 23020 16244
rect 22975 16204 23020 16232
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 25130 16232 25136 16244
rect 25091 16204 25136 16232
rect 25130 16192 25136 16204
rect 25188 16192 25194 16244
rect 7466 16124 7472 16176
rect 7524 16164 7530 16176
rect 7837 16167 7895 16173
rect 7837 16164 7849 16167
rect 7524 16136 7849 16164
rect 7524 16124 7530 16136
rect 7837 16133 7849 16136
rect 7883 16164 7895 16167
rect 8202 16164 8208 16176
rect 7883 16136 8208 16164
rect 7883 16133 7895 16136
rect 7837 16127 7895 16133
rect 8202 16124 8208 16136
rect 8260 16124 8266 16176
rect 10134 16164 10140 16176
rect 10095 16136 10140 16164
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 12575 16167 12633 16173
rect 12575 16133 12587 16167
rect 12621 16164 12633 16167
rect 13354 16164 13360 16176
rect 12621 16136 13360 16164
rect 12621 16133 12633 16136
rect 12575 16127 12633 16133
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 13446 16124 13452 16176
rect 13504 16164 13510 16176
rect 19150 16164 19156 16176
rect 13504 16136 13549 16164
rect 19111 16136 19156 16164
rect 13504 16124 13510 16136
rect 19150 16124 19156 16136
rect 19208 16164 19214 16176
rect 21085 16167 21143 16173
rect 21085 16164 21097 16167
rect 19208 16136 21097 16164
rect 19208 16124 19214 16136
rect 21085 16133 21097 16136
rect 21131 16164 21143 16167
rect 21910 16164 21916 16176
rect 21131 16136 21916 16164
rect 21131 16133 21143 16136
rect 21085 16127 21143 16133
rect 21910 16124 21916 16136
rect 21968 16124 21974 16176
rect 22204 16164 22232 16192
rect 23385 16167 23443 16173
rect 23385 16164 23397 16167
rect 22204 16136 23397 16164
rect 23385 16133 23397 16136
rect 23431 16133 23443 16167
rect 24762 16164 24768 16176
rect 23385 16127 23443 16133
rect 24228 16136 24768 16164
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16096 7159 16099
rect 8018 16096 8024 16108
rect 7147 16068 8024 16096
rect 7147 16065 7159 16068
rect 7101 16059 7159 16065
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16096 9643 16099
rect 9766 16096 9772 16108
rect 9631 16068 9772 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11330 16096 11336 16108
rect 11195 16068 11336 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11330 16056 11336 16068
rect 11388 16096 11394 16108
rect 12250 16096 12256 16108
rect 11388 16068 12256 16096
rect 11388 16056 11394 16068
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 13998 16096 14004 16108
rect 13911 16068 14004 16096
rect 13998 16056 14004 16068
rect 14056 16096 14062 16108
rect 15286 16096 15292 16108
rect 14056 16068 15292 16096
rect 14056 16056 14062 16068
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15562 16096 15568 16108
rect 15523 16068 15568 16096
rect 15562 16056 15568 16068
rect 15620 16096 15626 16108
rect 16485 16099 16543 16105
rect 16485 16096 16497 16099
rect 15620 16068 16497 16096
rect 15620 16056 15626 16068
rect 16485 16065 16497 16068
rect 16531 16065 16543 16099
rect 16485 16059 16543 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18598 16096 18604 16108
rect 17911 16068 18604 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 22094 16096 22100 16108
rect 22055 16068 22100 16096
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 24228 16105 24256 16136
rect 24762 16124 24768 16136
rect 24820 16124 24826 16176
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16065 24271 16099
rect 24213 16059 24271 16065
rect 24302 16056 24308 16108
rect 24360 16096 24366 16108
rect 24489 16099 24547 16105
rect 24489 16096 24501 16099
rect 24360 16068 24501 16096
rect 24360 16056 24366 16068
rect 24489 16065 24501 16068
rect 24535 16065 24547 16099
rect 24489 16059 24547 16065
rect 12472 16031 12530 16037
rect 12472 16028 12484 16031
rect 12176 16000 12484 16028
rect 8113 15963 8171 15969
rect 8113 15929 8125 15963
rect 8159 15929 8171 15963
rect 8113 15923 8171 15929
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15960 8723 15963
rect 8754 15960 8760 15972
rect 8711 15932 8760 15960
rect 8711 15929 8723 15932
rect 8665 15923 8723 15929
rect 7469 15895 7527 15901
rect 7469 15861 7481 15895
rect 7515 15892 7527 15895
rect 8128 15892 8156 15923
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 9401 15963 9459 15969
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 9677 15963 9735 15969
rect 9677 15960 9689 15963
rect 9447 15932 9689 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 9677 15929 9689 15932
rect 9723 15960 9735 15963
rect 10042 15960 10048 15972
rect 9723 15932 10048 15960
rect 9723 15929 9735 15932
rect 9677 15923 9735 15929
rect 9416 15892 9444 15923
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 11238 15920 11244 15972
rect 11296 15960 11302 15972
rect 12176 15969 12204 16000
rect 12472 15997 12484 16000
rect 12518 15997 12530 16031
rect 12472 15991 12530 15997
rect 18392 16031 18450 16037
rect 18392 15997 18404 16031
rect 18438 16028 18450 16031
rect 18800 16028 18828 16056
rect 18438 16000 18828 16028
rect 19613 16031 19671 16037
rect 18438 15997 18450 16000
rect 18392 15991 18450 15997
rect 19613 15997 19625 16031
rect 19659 15997 19671 16031
rect 19978 16028 19984 16040
rect 19939 16000 19984 16028
rect 19613 15991 19671 15997
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 11296 15932 12173 15960
rect 11296 15920 11302 15932
rect 12161 15929 12173 15932
rect 12207 15929 12219 15963
rect 12161 15923 12219 15929
rect 13081 15963 13139 15969
rect 13081 15929 13093 15963
rect 13127 15960 13139 15963
rect 13170 15960 13176 15972
rect 13127 15932 13176 15960
rect 13127 15929 13139 15932
rect 13081 15923 13139 15929
rect 13170 15920 13176 15932
rect 13228 15960 13234 15972
rect 13814 15960 13820 15972
rect 13228 15932 13820 15960
rect 13228 15920 13234 15932
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 14642 15960 14648 15972
rect 14148 15932 14193 15960
rect 14603 15932 14648 15960
rect 14148 15920 14154 15932
rect 14642 15920 14648 15932
rect 14700 15920 14706 15972
rect 15657 15963 15715 15969
rect 15657 15960 15669 15963
rect 14936 15932 15669 15960
rect 11330 15892 11336 15904
rect 7515 15864 9444 15892
rect 11291 15864 11336 15892
rect 7515 15861 7527 15864
rect 7469 15855 7527 15861
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11790 15892 11796 15904
rect 11751 15864 11796 15892
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 14826 15852 14832 15904
rect 14884 15892 14890 15904
rect 14936 15901 14964 15932
rect 15657 15929 15669 15932
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 15930 15920 15936 15972
rect 15988 15960 15994 15972
rect 16209 15963 16267 15969
rect 16209 15960 16221 15963
rect 15988 15932 16221 15960
rect 15988 15920 15994 15932
rect 16209 15929 16221 15932
rect 16255 15929 16267 15963
rect 17494 15960 17500 15972
rect 17407 15932 17500 15960
rect 16209 15923 16267 15929
rect 17494 15920 17500 15932
rect 17552 15960 17558 15972
rect 17552 15932 19472 15960
rect 17552 15920 17558 15932
rect 14921 15895 14979 15901
rect 14921 15892 14933 15895
rect 14884 15864 14933 15892
rect 14884 15852 14890 15864
rect 14921 15861 14933 15864
rect 14967 15861 14979 15895
rect 14921 15855 14979 15861
rect 15381 15895 15439 15901
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 16114 15892 16120 15904
rect 15427 15864 16120 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 16114 15852 16120 15864
rect 16172 15892 16178 15904
rect 16666 15892 16672 15904
rect 16172 15864 16672 15892
rect 16172 15852 16178 15864
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 17129 15895 17187 15901
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17770 15892 17776 15904
rect 17175 15864 17776 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 19444 15901 19472 15932
rect 19518 15920 19524 15972
rect 19576 15960 19582 15972
rect 19628 15960 19656 15991
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20162 16028 20168 16040
rect 20123 16000 20168 16028
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 20530 16028 20536 16040
rect 20491 16000 20536 16028
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 21913 15963 21971 15969
rect 19576 15932 20852 15960
rect 19576 15920 19582 15932
rect 20824 15904 20852 15932
rect 21913 15929 21925 15963
rect 21959 15960 21971 15963
rect 22186 15960 22192 15972
rect 21959 15932 22192 15960
rect 21959 15929 21971 15932
rect 21913 15923 21971 15929
rect 22186 15920 22192 15932
rect 22244 15920 22250 15972
rect 22741 15963 22799 15969
rect 22741 15929 22753 15963
rect 22787 15960 22799 15963
rect 24210 15960 24216 15972
rect 22787 15932 24216 15960
rect 22787 15929 22799 15932
rect 22741 15923 22799 15929
rect 24210 15920 24216 15932
rect 24268 15920 24274 15972
rect 24305 15963 24363 15969
rect 24305 15929 24317 15963
rect 24351 15929 24363 15963
rect 24305 15923 24363 15929
rect 19429 15895 19487 15901
rect 19429 15861 19441 15895
rect 19475 15861 19487 15895
rect 19429 15855 19487 15861
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 20864 15864 21465 15892
rect 20864 15852 20870 15864
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 24029 15895 24087 15901
rect 24029 15861 24041 15895
rect 24075 15892 24087 15895
rect 24118 15892 24124 15904
rect 24075 15864 24124 15892
rect 24075 15861 24087 15864
rect 24029 15855 24087 15861
rect 24118 15852 24124 15864
rect 24176 15892 24182 15904
rect 24320 15892 24348 15923
rect 24176 15864 24348 15892
rect 24176 15852 24182 15864
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 7834 15688 7840 15700
rect 7795 15660 7840 15688
rect 7834 15648 7840 15660
rect 7892 15688 7898 15700
rect 7892 15660 8156 15688
rect 7892 15648 7898 15660
rect 8128 15629 8156 15660
rect 9766 15648 9772 15700
rect 9824 15697 9830 15700
rect 9824 15691 9873 15697
rect 9824 15657 9827 15691
rect 9861 15657 9873 15691
rect 9824 15651 9873 15657
rect 9824 15648 9830 15651
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10413 15691 10471 15697
rect 10413 15688 10425 15691
rect 10192 15660 10425 15688
rect 10192 15648 10198 15660
rect 10413 15657 10425 15660
rect 10459 15657 10471 15691
rect 10413 15651 10471 15657
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 15381 15691 15439 15697
rect 15381 15688 15393 15691
rect 13412 15660 15393 15688
rect 13412 15648 13418 15660
rect 15381 15657 15393 15660
rect 15427 15657 15439 15691
rect 18598 15688 18604 15700
rect 18559 15660 18604 15688
rect 15381 15651 15439 15657
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 19518 15688 19524 15700
rect 19122 15660 19524 15688
rect 8113 15623 8171 15629
rect 8113 15589 8125 15623
rect 8159 15589 8171 15623
rect 8113 15583 8171 15589
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 11054 15620 11060 15632
rect 8260 15592 8305 15620
rect 11015 15592 11060 15620
rect 8260 15580 8266 15592
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 13998 15620 14004 15632
rect 13872 15592 14004 15620
rect 13872 15580 13878 15592
rect 13998 15580 14004 15592
rect 14056 15580 14062 15632
rect 14369 15623 14427 15629
rect 14369 15589 14381 15623
rect 14415 15620 14427 15623
rect 14642 15620 14648 15632
rect 14415 15592 14648 15620
rect 14415 15589 14427 15592
rect 14369 15583 14427 15589
rect 14642 15580 14648 15592
rect 14700 15580 14706 15632
rect 14734 15580 14740 15632
rect 14792 15620 14798 15632
rect 14829 15623 14887 15629
rect 14829 15620 14841 15623
rect 14792 15592 14841 15620
rect 14792 15580 14798 15592
rect 14829 15589 14841 15592
rect 14875 15589 14887 15623
rect 14829 15583 14887 15589
rect 17129 15623 17187 15629
rect 17129 15589 17141 15623
rect 17175 15620 17187 15623
rect 17494 15620 17500 15632
rect 17175 15592 17500 15620
rect 17175 15589 17187 15592
rect 17129 15583 17187 15589
rect 17494 15580 17500 15592
rect 17552 15580 17558 15632
rect 18049 15623 18107 15629
rect 18049 15589 18061 15623
rect 18095 15620 18107 15623
rect 18690 15620 18696 15632
rect 18095 15592 18696 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 18690 15580 18696 15592
rect 18748 15620 18754 15632
rect 19122 15620 19150 15660
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20530 15688 20536 15700
rect 20395 15660 20536 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 20990 15688 20996 15700
rect 20951 15660 20996 15688
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 23569 15691 23627 15697
rect 23569 15688 23581 15691
rect 23446 15660 23581 15688
rect 23446 15632 23474 15660
rect 23569 15657 23581 15660
rect 23615 15657 23627 15691
rect 23569 15651 23627 15657
rect 24026 15648 24032 15700
rect 24084 15688 24090 15700
rect 24121 15691 24179 15697
rect 24121 15688 24133 15691
rect 24084 15660 24133 15688
rect 24084 15648 24090 15660
rect 24121 15657 24133 15660
rect 24167 15657 24179 15691
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24121 15651 24179 15657
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 25130 15688 25136 15700
rect 25091 15660 25136 15688
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 20162 15620 20168 15632
rect 18748 15592 19150 15620
rect 19536 15592 20168 15620
rect 18748 15580 18754 15592
rect 9582 15552 9588 15564
rect 9543 15524 9588 15552
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 12710 15552 12716 15564
rect 12575 15524 12716 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 8754 15484 8760 15496
rect 8667 15456 8760 15484
rect 8754 15444 8760 15456
rect 8812 15484 8818 15496
rect 10962 15484 10968 15496
rect 8812 15456 10968 15484
rect 8812 15444 8818 15456
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11238 15484 11244 15496
rect 11199 15456 11244 15484
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 15304 15484 15332 15515
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 18800 15561 18828 15592
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 15436 15524 15761 15552
rect 15436 15512 15442 15524
rect 15749 15521 15761 15524
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15552 19303 15555
rect 19426 15552 19432 15564
rect 19291 15524 19432 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 19536 15561 19564 15592
rect 20162 15580 20168 15592
rect 20220 15620 20226 15632
rect 20438 15620 20444 15632
rect 20220 15592 20444 15620
rect 20220 15580 20226 15592
rect 20438 15580 20444 15592
rect 20496 15580 20502 15632
rect 23382 15580 23388 15632
rect 23440 15592 23474 15632
rect 24489 15623 24547 15629
rect 23440 15580 23446 15592
rect 24489 15589 24501 15623
rect 24535 15620 24547 15623
rect 24670 15620 24676 15632
rect 24535 15592 24676 15620
rect 24535 15589 24547 15592
rect 24489 15583 24547 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 15654 15484 15660 15496
rect 15304 15456 15660 15484
rect 13725 15447 13783 15453
rect 12759 15419 12817 15425
rect 12759 15385 12771 15419
rect 12805 15416 12817 15419
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 12805 15388 13461 15416
rect 12805 15385 12817 15388
rect 12759 15379 12817 15385
rect 13449 15385 13461 15388
rect 13495 15416 13507 15419
rect 13740 15416 13768 15447
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15484 16911 15487
rect 17037 15487 17095 15493
rect 17037 15484 17049 15487
rect 16899 15456 17049 15484
rect 16899 15453 16911 15456
rect 16853 15447 16911 15453
rect 17037 15453 17049 15456
rect 17083 15484 17095 15487
rect 17126 15484 17132 15496
rect 17083 15456 17132 15484
rect 17083 15453 17095 15456
rect 17037 15447 17095 15453
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15484 17739 15487
rect 18874 15484 18880 15496
rect 17727 15456 18880 15484
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 19720 15484 19748 15515
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20864 15524 20913 15552
rect 20864 15512 20870 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15521 21511 15555
rect 21726 15552 21732 15564
rect 21687 15524 21732 15552
rect 21453 15515 21511 15521
rect 20346 15484 20352 15496
rect 19162 15456 20352 15484
rect 13495 15388 13768 15416
rect 18417 15419 18475 15425
rect 13495 15385 13507 15388
rect 13449 15379 13507 15385
rect 18417 15385 18429 15419
rect 18463 15416 18475 15419
rect 19162 15416 19190 15456
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 21468 15484 21496 15515
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21876 15524 22109 15552
rect 21876 15512 21882 15524
rect 22097 15521 22109 15524
rect 22143 15521 22155 15555
rect 24946 15552 24952 15564
rect 24907 15524 24952 15552
rect 22097 15515 22155 15521
rect 24946 15512 24952 15524
rect 25004 15512 25010 15564
rect 21237 15456 21496 15484
rect 18463 15388 19190 15416
rect 18463 15385 18475 15388
rect 18417 15379 18475 15385
rect 20162 15376 20168 15428
rect 20220 15416 20226 15428
rect 21082 15416 21088 15428
rect 20220 15388 21088 15416
rect 20220 15376 20226 15388
rect 21082 15376 21088 15388
rect 21140 15416 21146 15428
rect 21237 15416 21265 15456
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23201 15487 23259 15493
rect 23201 15484 23213 15487
rect 22980 15456 23213 15484
rect 22980 15444 22986 15456
rect 23201 15453 23213 15456
rect 23247 15453 23259 15487
rect 23201 15447 23259 15453
rect 21140 15388 21265 15416
rect 21140 15376 21146 15388
rect 13078 15348 13084 15360
rect 13039 15320 13084 15348
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 16482 15348 16488 15360
rect 16443 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 20806 15348 20812 15360
rect 20763 15320 20812 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 9582 15104 9588 15156
rect 9640 15144 9646 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 9640 15116 9965 15144
rect 9640 15104 9646 15116
rect 9953 15113 9965 15116
rect 9999 15144 10011 15147
rect 10870 15144 10876 15156
rect 9999 15116 10876 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11425 15147 11483 15153
rect 11425 15144 11437 15147
rect 11112 15116 11437 15144
rect 11112 15104 11118 15116
rect 11425 15113 11437 15116
rect 11471 15144 11483 15147
rect 11974 15144 11980 15156
rect 11471 15116 11980 15144
rect 11471 15113 11483 15116
rect 11425 15107 11483 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12710 15144 12716 15156
rect 12492 15116 12716 15144
rect 12492 15104 12498 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 13906 15104 13912 15156
rect 13964 15144 13970 15156
rect 14737 15147 14795 15153
rect 14737 15144 14749 15147
rect 13964 15116 14749 15144
rect 13964 15104 13970 15116
rect 14737 15113 14749 15116
rect 14783 15144 14795 15147
rect 15378 15144 15384 15156
rect 14783 15116 15384 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 19245 15147 19303 15153
rect 19245 15144 19257 15147
rect 17911 15116 19257 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 19245 15113 19257 15116
rect 19291 15144 19303 15147
rect 19426 15144 19432 15156
rect 19291 15116 19432 15144
rect 19291 15113 19303 15116
rect 19245 15107 19303 15113
rect 19426 15104 19432 15116
rect 19484 15144 19490 15156
rect 20162 15144 20168 15156
rect 19484 15116 20168 15144
rect 19484 15104 19490 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 23934 15144 23940 15156
rect 22244 15116 23940 15144
rect 22244 15104 22250 15116
rect 23934 15104 23940 15116
rect 23992 15144 23998 15156
rect 24581 15147 24639 15153
rect 24581 15144 24593 15147
rect 23992 15116 24593 15144
rect 23992 15104 23998 15116
rect 24581 15113 24593 15116
rect 24627 15113 24639 15147
rect 24946 15144 24952 15156
rect 24907 15116 24952 15144
rect 24581 15107 24639 15113
rect 24946 15104 24952 15116
rect 25004 15144 25010 15156
rect 25547 15147 25605 15153
rect 25547 15144 25559 15147
rect 25004 15116 25559 15144
rect 25004 15104 25010 15116
rect 25547 15113 25559 15116
rect 25593 15113 25605 15147
rect 25547 15107 25605 15113
rect 14001 15079 14059 15085
rect 14001 15045 14013 15079
rect 14047 15076 14059 15079
rect 14826 15076 14832 15088
rect 14047 15048 14832 15076
rect 14047 15045 14059 15048
rect 14001 15039 14059 15045
rect 14826 15036 14832 15048
rect 14884 15036 14890 15088
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 15933 15079 15991 15085
rect 15933 15076 15945 15079
rect 15712 15048 15945 15076
rect 15712 15036 15718 15048
rect 15933 15045 15945 15048
rect 15979 15076 15991 15079
rect 17678 15076 17684 15088
rect 15979 15048 17684 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 21085 15079 21143 15085
rect 21085 15076 21097 15079
rect 20772 15048 21097 15076
rect 20772 15036 20778 15048
rect 21085 15045 21097 15048
rect 21131 15045 21143 15079
rect 21085 15039 21143 15045
rect 21910 15036 21916 15088
rect 21968 15076 21974 15088
rect 23017 15079 23075 15085
rect 23017 15076 23029 15079
rect 21968 15048 23029 15076
rect 21968 15036 21974 15048
rect 23017 15045 23029 15048
rect 23063 15076 23075 15079
rect 23382 15076 23388 15088
rect 23063 15048 23388 15076
rect 23063 15045 23075 15048
rect 23017 15039 23075 15045
rect 23382 15036 23388 15048
rect 23440 15076 23446 15088
rect 23440 15048 24072 15076
rect 23440 15036 23446 15048
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 9217 15011 9275 15017
rect 9217 15008 9229 15011
rect 8067 14980 9229 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 9217 14977 9229 14980
rect 9263 15008 9275 15011
rect 10134 15008 10140 15020
rect 9263 14980 10140 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 10134 14968 10140 14980
rect 10192 15008 10198 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10192 14980 10517 15008
rect 10192 14968 10198 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 13078 15008 13084 15020
rect 13039 14980 13084 15008
rect 10505 14971 10563 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14700 14980 15209 15008
rect 14700 14968 14706 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 17126 15008 17132 15020
rect 17039 14980 17132 15008
rect 15197 14971 15255 14977
rect 17126 14968 17132 14980
rect 17184 15008 17190 15020
rect 18414 15008 18420 15020
rect 17184 14980 18420 15008
rect 17184 14968 17190 14980
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 15008 18843 15011
rect 18874 15008 18880 15020
rect 18831 14980 18880 15008
rect 18831 14977 18843 14980
rect 18785 14971 18843 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 20806 15008 20812 15020
rect 19996 14980 20812 15008
rect 11330 14900 11336 14952
rect 11388 14940 11394 14952
rect 11388 14912 13814 14940
rect 11388 14900 11394 14912
rect 7374 14872 7380 14884
rect 7335 14844 7380 14872
rect 7374 14832 7380 14844
rect 7432 14832 7438 14884
rect 7466 14832 7472 14884
rect 7524 14872 7530 14884
rect 8757 14875 8815 14881
rect 7524 14844 7569 14872
rect 7524 14832 7530 14844
rect 8757 14841 8769 14875
rect 8803 14872 8815 14875
rect 8938 14872 8944 14884
rect 8803 14844 8944 14872
rect 8803 14841 8815 14844
rect 8757 14835 8815 14841
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 9030 14832 9036 14884
rect 9088 14872 9094 14884
rect 10597 14875 10655 14881
rect 9088 14844 9133 14872
rect 9088 14832 9094 14844
rect 10597 14841 10609 14875
rect 10643 14841 10655 14875
rect 10597 14835 10655 14841
rect 11149 14875 11207 14881
rect 11149 14841 11161 14875
rect 11195 14872 11207 14875
rect 11238 14872 11244 14884
rect 11195 14844 11244 14872
rect 11195 14841 11207 14844
rect 11149 14835 11207 14841
rect 7193 14807 7251 14813
rect 7193 14773 7205 14807
rect 7239 14804 7251 14807
rect 7484 14804 7512 14832
rect 7239 14776 7512 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8260 14776 8401 14804
rect 8260 14764 8266 14776
rect 8389 14773 8401 14776
rect 8435 14804 8447 14807
rect 9048 14804 9076 14832
rect 8435 14776 9076 14804
rect 10321 14807 10379 14813
rect 8435 14773 8447 14776
rect 8389 14767 8447 14773
rect 10321 14773 10333 14807
rect 10367 14804 10379 14807
rect 10612 14804 10640 14835
rect 11238 14832 11244 14844
rect 11296 14832 11302 14884
rect 13443 14875 13501 14881
rect 13443 14841 13455 14875
rect 13489 14872 13501 14875
rect 13630 14872 13636 14884
rect 13489 14844 13636 14872
rect 13489 14841 13501 14844
rect 13443 14835 13501 14841
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 13786 14872 13814 14912
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 19996 14949 20024 14980
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 14056 14912 14289 14940
rect 14056 14900 14062 14912
rect 14277 14909 14289 14912
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14909 20039 14943
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 19981 14903 20039 14909
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 14918 14872 14924 14884
rect 13786 14844 14924 14872
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 15013 14875 15071 14881
rect 15013 14841 15025 14875
rect 15059 14841 15071 14875
rect 16482 14872 16488 14884
rect 16443 14844 16488 14872
rect 15013 14835 15071 14841
rect 10686 14804 10692 14816
rect 10367 14776 10692 14804
rect 10367 14773 10379 14776
rect 10321 14767 10379 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 13906 14804 13912 14816
rect 12768 14776 13912 14804
rect 12768 14764 12774 14776
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15028 14804 15056 14835
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 16577 14875 16635 14881
rect 16577 14841 16589 14875
rect 16623 14872 16635 14875
rect 16666 14872 16672 14884
rect 16623 14844 16672 14872
rect 16623 14841 16635 14844
rect 16577 14835 16635 14841
rect 14792 14776 15056 14804
rect 16301 14807 16359 14813
rect 14792 14764 14798 14776
rect 16301 14773 16313 14807
rect 16347 14804 16359 14807
rect 16592 14804 16620 14835
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 17494 14872 17500 14884
rect 17407 14844 17500 14872
rect 17494 14832 17500 14844
rect 17552 14872 17558 14884
rect 17954 14872 17960 14884
rect 17552 14844 17960 14872
rect 17552 14832 17558 14844
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 18138 14872 18144 14884
rect 18099 14844 18144 14872
rect 18138 14832 18144 14844
rect 18196 14832 18202 14884
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14841 18291 14875
rect 18233 14835 18291 14841
rect 16347 14776 16620 14804
rect 16347 14773 16359 14776
rect 16301 14767 16359 14773
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 18248 14804 18276 14835
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 19521 14875 19579 14881
rect 19521 14872 19533 14875
rect 19116 14844 19533 14872
rect 19116 14832 19122 14844
rect 19521 14841 19533 14844
rect 19567 14872 19579 14875
rect 20548 14872 20576 14903
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20680 14912 20913 14940
rect 20680 14900 20686 14912
rect 20901 14909 20913 14912
rect 20947 14940 20959 14943
rect 20990 14940 20996 14952
rect 20947 14912 20996 14940
rect 20947 14909 20959 14912
rect 20901 14903 20959 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14909 22063 14943
rect 23658 14940 23664 14952
rect 23619 14912 23664 14940
rect 22005 14903 22063 14909
rect 21453 14875 21511 14881
rect 21453 14872 21465 14875
rect 19567 14844 21465 14872
rect 19567 14841 19579 14844
rect 19521 14835 19579 14841
rect 21453 14841 21465 14844
rect 21499 14872 21511 14875
rect 21726 14872 21732 14884
rect 21499 14844 21732 14872
rect 21499 14841 21511 14844
rect 21453 14835 21511 14841
rect 21726 14832 21732 14844
rect 21784 14832 21790 14884
rect 22020 14872 22048 14903
rect 23658 14900 23664 14912
rect 23716 14900 23722 14952
rect 22557 14875 22615 14881
rect 22557 14872 22569 14875
rect 22020 14844 22569 14872
rect 22557 14841 22569 14844
rect 22603 14872 22615 14875
rect 23106 14872 23112 14884
rect 22603 14844 23112 14872
rect 22603 14841 22615 14844
rect 22557 14835 22615 14841
rect 23106 14832 23112 14844
rect 23164 14832 23170 14884
rect 18874 14804 18880 14816
rect 17920 14776 18880 14804
rect 17920 14764 17926 14776
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 21818 14804 21824 14816
rect 20404 14776 21824 14804
rect 20404 14764 20410 14776
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 22186 14804 22192 14816
rect 22147 14776 22192 14804
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 24044 14813 24072 15048
rect 24210 14900 24216 14952
rect 24268 14940 24274 14952
rect 25444 14943 25502 14949
rect 25444 14940 25456 14943
rect 24268 14912 25456 14940
rect 24268 14900 24274 14912
rect 25444 14909 25456 14912
rect 25490 14940 25502 14943
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25490 14912 25881 14940
rect 25490 14909 25502 14912
rect 25444 14903 25502 14909
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 24029 14807 24087 14813
rect 24029 14773 24041 14807
rect 24075 14773 24087 14807
rect 24029 14767 24087 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 8996 14572 9689 14600
rect 8996 14560 9002 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 10962 14600 10968 14612
rect 10923 14572 10968 14600
rect 9677 14563 9735 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11422 14600 11428 14612
rect 11383 14572 11428 14600
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 11974 14600 11980 14612
rect 11935 14572 11980 14600
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 12710 14600 12716 14612
rect 12667 14572 12716 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 14918 14600 14924 14612
rect 14879 14572 14924 14600
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15427 14603 15485 14609
rect 15427 14600 15439 14603
rect 15344 14572 15439 14600
rect 15344 14560 15350 14572
rect 15427 14569 15439 14572
rect 15473 14569 15485 14603
rect 17310 14600 17316 14612
rect 15427 14563 15485 14569
rect 16316 14572 17316 14600
rect 8389 14535 8447 14541
rect 8389 14501 8401 14535
rect 8435 14532 8447 14535
rect 9030 14532 9036 14544
rect 8435 14504 9036 14532
rect 8435 14501 8447 14504
rect 8389 14495 8447 14501
rect 9030 14492 9036 14504
rect 9088 14492 9094 14544
rect 11440 14532 11468 14560
rect 13081 14535 13139 14541
rect 13081 14532 13093 14535
rect 11440 14504 13093 14532
rect 13081 14501 13093 14504
rect 13127 14532 13139 14535
rect 13630 14532 13636 14544
rect 13127 14504 13636 14532
rect 13127 14501 13139 14504
rect 13081 14495 13139 14501
rect 13630 14492 13636 14504
rect 13688 14541 13694 14544
rect 13688 14535 13736 14541
rect 13688 14501 13690 14535
rect 13724 14501 13736 14535
rect 13688 14495 13736 14501
rect 13688 14492 13694 14495
rect 8624 14467 8682 14473
rect 8624 14433 8636 14467
rect 8670 14464 8682 14467
rect 8846 14464 8852 14476
rect 8670 14436 8852 14464
rect 8670 14433 8682 14436
rect 8624 14427 8682 14433
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 11146 14464 11152 14476
rect 11103 14436 11152 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 13354 14464 13360 14476
rect 13315 14436 13360 14464
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 15378 14473 15384 14476
rect 15356 14467 15384 14473
rect 15356 14464 15368 14467
rect 15291 14436 15368 14464
rect 15356 14433 15368 14436
rect 15436 14464 15442 14476
rect 16316 14464 16344 14572
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17589 14603 17647 14609
rect 17589 14569 17601 14603
rect 17635 14600 17647 14603
rect 17862 14600 17868 14612
rect 17635 14572 17868 14600
rect 17635 14569 17647 14572
rect 17589 14563 17647 14569
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 23658 14600 23664 14612
rect 23446 14572 23664 14600
rect 16666 14532 16672 14544
rect 16627 14504 16672 14532
rect 16666 14492 16672 14504
rect 16724 14492 16730 14544
rect 17218 14532 17224 14544
rect 17131 14504 17224 14532
rect 17218 14492 17224 14504
rect 17276 14532 17282 14544
rect 18138 14532 18144 14544
rect 17276 14504 18144 14532
rect 17276 14492 17282 14504
rect 18138 14492 18144 14504
rect 18196 14492 18202 14544
rect 18230 14492 18236 14544
rect 18288 14532 18294 14544
rect 18288 14504 18333 14532
rect 18288 14492 18294 14504
rect 21818 14492 21824 14544
rect 21876 14532 21882 14544
rect 23017 14535 23075 14541
rect 21876 14504 22784 14532
rect 21876 14492 21882 14504
rect 15436 14436 16344 14464
rect 15356 14427 15384 14433
rect 15378 14424 15384 14427
rect 15436 14424 15442 14436
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19484 14436 19625 14464
rect 19484 14424 19490 14436
rect 19613 14433 19625 14436
rect 19659 14464 19671 14467
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19659 14436 20085 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 21726 14464 21732 14476
rect 21687 14436 21732 14464
rect 20073 14427 20131 14433
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 7374 14396 7380 14408
rect 7287 14368 7380 14396
rect 7374 14356 7380 14368
rect 7432 14396 7438 14408
rect 8711 14399 8769 14405
rect 8711 14396 8723 14399
rect 7432 14368 8723 14396
rect 7432 14356 7438 14368
rect 8711 14365 8723 14368
rect 8757 14365 8769 14399
rect 8711 14359 8769 14365
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 16577 14399 16635 14405
rect 16577 14396 16589 14399
rect 15528 14368 16589 14396
rect 15528 14356 15534 14368
rect 16577 14365 16589 14368
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 17460 14368 18153 14396
rect 17460 14356 17466 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18414 14396 18420 14408
rect 18375 14368 18420 14396
rect 18141 14359 18199 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 21082 14356 21088 14408
rect 21140 14396 21146 14408
rect 22020 14396 22048 14427
rect 22186 14424 22192 14476
rect 22244 14464 22250 14476
rect 22370 14464 22376 14476
rect 22244 14436 22376 14464
rect 22244 14424 22250 14436
rect 22370 14424 22376 14436
rect 22428 14424 22434 14476
rect 22756 14473 22784 14504
rect 23017 14501 23029 14535
rect 23063 14532 23075 14535
rect 23446 14532 23474 14572
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 24118 14600 24124 14612
rect 24079 14572 24124 14600
rect 24118 14560 24124 14572
rect 24176 14560 24182 14612
rect 23063 14504 23474 14532
rect 23063 14501 23075 14504
rect 23017 14495 23075 14501
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 22830 14464 22836 14476
rect 22787 14436 22836 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 22830 14424 22836 14436
rect 22888 14424 22894 14476
rect 23934 14464 23940 14476
rect 23895 14436 23940 14464
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 25406 14464 25412 14476
rect 25367 14436 25412 14464
rect 25406 14424 25412 14436
rect 25464 14424 25470 14476
rect 21140 14368 22048 14396
rect 21140 14356 21146 14368
rect 17957 14331 18015 14337
rect 17957 14297 17969 14331
rect 18003 14328 18015 14331
rect 18966 14328 18972 14340
rect 18003 14300 18972 14328
rect 18003 14297 18015 14300
rect 17957 14291 18015 14297
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 19337 14331 19395 14337
rect 19337 14297 19349 14331
rect 19383 14328 19395 14331
rect 20070 14328 20076 14340
rect 19383 14300 20076 14328
rect 19383 14297 19395 14300
rect 19337 14291 19395 14297
rect 20070 14288 20076 14300
rect 20128 14288 20134 14340
rect 20533 14331 20591 14337
rect 20533 14297 20545 14331
rect 20579 14328 20591 14331
rect 20806 14328 20812 14340
rect 20579 14300 20812 14328
rect 20579 14297 20591 14300
rect 20533 14291 20591 14297
rect 20806 14288 20812 14300
rect 20864 14328 20870 14340
rect 25593 14331 25651 14337
rect 25593 14328 25605 14331
rect 20864 14300 25605 14328
rect 20864 14288 20870 14300
rect 25593 14297 25605 14300
rect 25639 14297 25651 14331
rect 25593 14291 25651 14297
rect 7926 14260 7932 14272
rect 7887 14232 7932 14260
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 10137 14263 10195 14269
rect 10137 14260 10149 14263
rect 9548 14232 10149 14260
rect 9548 14220 9554 14232
rect 10137 14229 10149 14232
rect 10183 14229 10195 14263
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 10137 14223 10195 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 18196 14232 19809 14260
rect 18196 14220 18202 14232
rect 19797 14229 19809 14232
rect 19843 14229 19855 14263
rect 19797 14223 19855 14229
rect 22922 14220 22928 14272
rect 22980 14260 22986 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 22980 14232 23305 14260
rect 22980 14220 22986 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10686 14056 10692 14068
rect 10459 14028 10692 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 11146 14056 11152 14068
rect 10827 14028 11152 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 14274 14056 14280 14068
rect 14235 14028 14280 14056
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15528 14028 15853 14056
rect 15528 14016 15534 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 16206 14056 16212 14068
rect 16167 14028 16212 14056
rect 15841 14019 15899 14025
rect 16206 14016 16212 14028
rect 16264 14056 16270 14068
rect 16390 14056 16396 14068
rect 16264 14028 16396 14056
rect 16264 14016 16270 14028
rect 16390 14016 16396 14028
rect 16448 14056 16454 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 16448 14028 17785 14056
rect 16448 14016 16454 14028
rect 17773 14025 17785 14028
rect 17819 14056 17831 14059
rect 18230 14056 18236 14068
rect 17819 14028 18236 14056
rect 17819 14025 17831 14028
rect 17773 14019 17831 14025
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19334 14056 19340 14068
rect 19199 14028 19340 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19334 14016 19340 14028
rect 19392 14056 19398 14068
rect 19518 14056 19524 14068
rect 19392 14028 19524 14056
rect 19392 14016 19398 14028
rect 19518 14016 19524 14028
rect 19576 14016 19582 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 21140 14028 21189 14056
rect 21140 14016 21146 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 22830 14016 22836 14068
rect 22888 14056 22894 14068
rect 22925 14059 22983 14065
rect 22925 14056 22937 14059
rect 22888 14028 22937 14056
rect 22888 14016 22894 14028
rect 22925 14025 22937 14028
rect 22971 14025 22983 14059
rect 23934 14056 23940 14068
rect 23895 14028 23940 14056
rect 22925 14019 22983 14025
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 24351 14059 24409 14065
rect 24351 14025 24363 14059
rect 24397 14056 24409 14059
rect 24854 14056 24860 14068
rect 24397 14028 24860 14056
rect 24397 14025 24409 14028
rect 24351 14019 24409 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 11517 13991 11575 13997
rect 11517 13988 11529 13991
rect 9600 13960 11529 13988
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 9490 13920 9496 13932
rect 8711 13892 9496 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 7926 13852 7932 13864
rect 6788 13824 7932 13852
rect 6788 13812 6794 13824
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8404 13784 8432 13815
rect 9600 13784 9628 13960
rect 11517 13957 11529 13960
rect 11563 13988 11575 13991
rect 11790 13988 11796 14000
rect 11563 13960 11796 13988
rect 11563 13957 11575 13960
rect 11517 13951 11575 13957
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 13136 13960 13216 13988
rect 13136 13948 13142 13960
rect 13188 13929 13216 13960
rect 14366 13948 14372 14000
rect 14424 13948 14430 14000
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 20438 13988 20444 14000
rect 19024 13960 20444 13988
rect 19024 13948 19030 13960
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 20898 13948 20904 14000
rect 20956 13988 20962 14000
rect 25406 13988 25412 14000
rect 20956 13960 25412 13988
rect 20956 13948 20962 13960
rect 25406 13948 25412 13960
rect 25464 13988 25470 14000
rect 25685 13991 25743 13997
rect 25685 13988 25697 13991
rect 25464 13960 25697 13988
rect 25464 13948 25470 13960
rect 25685 13957 25697 13960
rect 25731 13957 25743 13991
rect 25685 13951 25743 13957
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 14384 13920 14412 13948
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 14384 13892 14473 13920
rect 13173 13883 13231 13889
rect 14461 13889 14473 13892
rect 14507 13920 14519 13923
rect 14642 13920 14648 13932
rect 14507 13892 14648 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 16356 13892 16497 13920
rect 16356 13880 16362 13892
rect 16485 13889 16497 13892
rect 16531 13889 16543 13923
rect 16485 13883 16543 13889
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17218 13920 17224 13932
rect 17175 13892 17224 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 20806 13920 20812 13932
rect 19208 13892 20812 13920
rect 19208 13880 19214 13892
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13852 11391 13855
rect 12710 13852 12716 13864
rect 11379 13824 11928 13852
rect 12671 13824 12716 13852
rect 11379 13821 11391 13824
rect 11333 13815 11391 13821
rect 11900 13796 11928 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12912 13824 13001 13852
rect 8404 13756 9628 13784
rect 9855 13787 9913 13793
rect 7837 13719 7895 13725
rect 7837 13685 7849 13719
rect 7883 13716 7895 13719
rect 8404 13716 8432 13756
rect 9855 13753 9867 13787
rect 9901 13784 9913 13787
rect 10134 13784 10140 13796
rect 9901 13756 10140 13784
rect 9901 13753 9913 13756
rect 9855 13747 9913 13753
rect 8478 13716 8484 13728
rect 7883 13688 8484 13716
rect 7883 13685 7895 13688
rect 7837 13679 7895 13685
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8904 13688 8953 13716
rect 8904 13676 8910 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 8941 13679 8999 13685
rect 9401 13719 9459 13725
rect 9401 13685 9413 13719
rect 9447 13716 9459 13719
rect 9870 13716 9898 13747
rect 10134 13744 10140 13756
rect 10192 13784 10198 13796
rect 11149 13787 11207 13793
rect 11149 13784 11161 13787
rect 10192 13756 11161 13784
rect 10192 13744 10198 13756
rect 11149 13753 11161 13756
rect 11195 13784 11207 13787
rect 11422 13784 11428 13796
rect 11195 13756 11428 13784
rect 11195 13753 11207 13756
rect 11149 13747 11207 13753
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 11882 13784 11888 13796
rect 11795 13756 11888 13784
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 12250 13784 12256 13796
rect 12211 13756 12256 13784
rect 12250 13744 12256 13756
rect 12308 13784 12314 13796
rect 12912 13784 12940 13824
rect 12989 13821 13001 13824
rect 13035 13852 13047 13855
rect 13078 13852 13084 13864
rect 13035 13824 13084 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 17310 13812 17316 13864
rect 17368 13852 17374 13864
rect 19536 13861 19564 13892
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 26053 13923 26111 13929
rect 26053 13920 26065 13923
rect 25291 13892 26065 13920
rect 18176 13855 18234 13861
rect 18176 13852 18188 13855
rect 17368 13824 18188 13852
rect 17368 13812 17374 13824
rect 18176 13821 18188 13824
rect 18222 13852 18234 13855
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18222 13824 18613 13852
rect 18222 13821 18234 13824
rect 18176 13815 18234 13821
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19499 13824 19533 13852
rect 18601 13815 18659 13821
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 19521 13815 19579 13821
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19668 13824 19717 13852
rect 19668 13812 19674 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 20070 13852 20076 13864
rect 20031 13824 20076 13852
rect 19705 13815 19763 13821
rect 20070 13812 20076 13824
rect 20128 13852 20134 13864
rect 20128 13824 20300 13852
rect 20128 13812 20134 13824
rect 13630 13784 13636 13796
rect 12308 13756 12940 13784
rect 13591 13756 13636 13784
rect 12308 13744 12314 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 14274 13744 14280 13796
rect 14332 13784 14338 13796
rect 14553 13787 14611 13793
rect 14553 13784 14565 13787
rect 14332 13756 14565 13784
rect 14332 13744 14338 13756
rect 14553 13753 14565 13756
rect 14599 13753 14611 13787
rect 14553 13747 14611 13753
rect 15105 13787 15163 13793
rect 15105 13753 15117 13787
rect 15151 13784 15163 13787
rect 15930 13784 15936 13796
rect 15151 13756 15936 13784
rect 15151 13753 15163 13756
rect 15105 13747 15163 13753
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 16298 13744 16304 13796
rect 16356 13784 16362 13796
rect 16577 13787 16635 13793
rect 16577 13784 16589 13787
rect 16356 13756 16589 13784
rect 16356 13744 16362 13756
rect 16577 13753 16589 13756
rect 16623 13753 16635 13787
rect 16577 13747 16635 13753
rect 15378 13716 15384 13728
rect 9447 13688 9898 13716
rect 15339 13688 15384 13716
rect 9447 13685 9459 13688
rect 9401 13679 9459 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 17402 13716 17408 13728
rect 17363 13688 17408 13716
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 18279 13719 18337 13725
rect 18279 13716 18291 13719
rect 18012 13688 18291 13716
rect 18012 13676 18018 13688
rect 18279 13685 18291 13688
rect 18325 13685 18337 13719
rect 19334 13716 19340 13728
rect 19295 13688 19340 13716
rect 18279 13679 18337 13685
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 20272 13716 20300 13824
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 20404 13824 20453 13852
rect 20404 13812 20410 13824
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 22002 13812 22008 13864
rect 22060 13852 22066 13864
rect 22132 13855 22190 13861
rect 22132 13852 22144 13855
rect 22060 13824 22144 13852
rect 22060 13812 22066 13824
rect 22132 13821 22144 13824
rect 22178 13852 22190 13855
rect 22557 13855 22615 13861
rect 22557 13852 22569 13855
rect 22178 13824 22569 13852
rect 22178 13821 22190 13824
rect 22132 13815 22190 13821
rect 22557 13821 22569 13824
rect 22603 13821 22615 13855
rect 22557 13815 22615 13821
rect 24946 13812 24952 13864
rect 25004 13852 25010 13864
rect 25291 13861 25319 13892
rect 26053 13889 26065 13892
rect 26099 13889 26111 13923
rect 26053 13883 26111 13889
rect 25276 13855 25334 13861
rect 25276 13852 25288 13855
rect 25004 13824 25288 13852
rect 25004 13812 25010 13824
rect 25276 13821 25288 13824
rect 25322 13821 25334 13855
rect 25276 13815 25334 13821
rect 25363 13855 25421 13861
rect 25363 13821 25375 13855
rect 25409 13852 25421 13855
rect 25498 13852 25504 13864
rect 25409 13824 25504 13852
rect 25409 13821 25421 13824
rect 25363 13815 25421 13821
rect 25498 13812 25504 13824
rect 25556 13812 25562 13864
rect 21542 13716 21548 13728
rect 20272 13688 21548 13716
rect 21542 13676 21548 13688
rect 21600 13676 21606 13728
rect 21726 13676 21732 13728
rect 21784 13716 21790 13728
rect 21913 13719 21971 13725
rect 21913 13716 21925 13719
rect 21784 13688 21925 13716
rect 21784 13676 21790 13688
rect 21913 13685 21925 13688
rect 21959 13685 21971 13719
rect 21913 13679 21971 13685
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22235 13719 22293 13725
rect 22235 13716 22247 13719
rect 22152 13688 22247 13716
rect 22152 13676 22158 13688
rect 22235 13685 22247 13688
rect 22281 13685 22293 13719
rect 22235 13679 22293 13685
rect 24121 13719 24179 13725
rect 24121 13685 24133 13719
rect 24167 13716 24179 13719
rect 24210 13716 24216 13728
rect 24167 13688 24216 13716
rect 24167 13685 24179 13688
rect 24121 13679 24179 13685
rect 24210 13676 24216 13688
rect 24268 13716 24274 13728
rect 24673 13719 24731 13725
rect 24673 13716 24685 13719
rect 24268 13688 24685 13716
rect 24268 13676 24274 13688
rect 24673 13685 24685 13688
rect 24719 13685 24731 13719
rect 24673 13679 24731 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 12802 13512 12808 13524
rect 8168 13484 12808 13512
rect 8168 13472 8174 13484
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13412 13484 13829 13512
rect 13412 13472 13418 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14424 13484 14657 13512
rect 14424 13472 14430 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 14645 13475 14703 13481
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16264 13484 16957 13512
rect 16264 13472 16270 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 16945 13475 17003 13481
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19518 13512 19524 13524
rect 19383 13484 19524 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19518 13472 19524 13484
rect 19576 13512 19582 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19576 13484 19901 13512
rect 19576 13472 19582 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21269 13515 21327 13521
rect 21269 13512 21281 13515
rect 21140 13484 21281 13512
rect 21140 13472 21146 13484
rect 21269 13481 21281 13484
rect 21315 13481 21327 13515
rect 21269 13475 21327 13481
rect 25455 13515 25513 13521
rect 25455 13481 25467 13515
rect 25501 13512 25513 13515
rect 25590 13512 25596 13524
rect 25501 13484 25596 13512
rect 25501 13481 25513 13484
rect 25455 13475 25513 13481
rect 9030 13404 9036 13456
rect 9088 13444 9094 13456
rect 9861 13447 9919 13453
rect 9861 13444 9873 13447
rect 9088 13416 9873 13444
rect 9088 13404 9094 13416
rect 9861 13413 9873 13416
rect 9907 13413 9919 13447
rect 15746 13444 15752 13456
rect 15707 13416 15752 13444
rect 9861 13407 9919 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 18319 13447 18377 13453
rect 18319 13413 18331 13447
rect 18365 13444 18377 13447
rect 18782 13444 18788 13456
rect 18365 13416 18788 13444
rect 18365 13413 18377 13416
rect 18319 13407 18377 13413
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 21284 13444 21312 13475
rect 25590 13472 25596 13484
rect 25648 13472 25654 13524
rect 22922 13444 22928 13456
rect 21284 13416 21956 13444
rect 22883 13416 22928 13444
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13345 8355 13379
rect 8478 13376 8484 13388
rect 8439 13348 8484 13376
rect 8297 13339 8355 13345
rect 8312 13308 8340 13339
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 11292 13379 11350 13385
rect 11292 13345 11304 13379
rect 11338 13376 11350 13379
rect 11974 13376 11980 13388
rect 11338 13348 11980 13376
rect 11338 13345 11350 13348
rect 11292 13339 11350 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13376 12771 13379
rect 12802 13376 12808 13388
rect 12759 13348 12808 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 12986 13376 12992 13388
rect 12947 13348 12992 13376
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 17494 13336 17500 13388
rect 17552 13376 17558 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17552 13348 17969 13376
rect 17552 13336 17558 13348
rect 17957 13345 17969 13348
rect 18003 13376 18015 13379
rect 19334 13376 19340 13388
rect 18003 13348 19340 13376
rect 18003 13345 18015 13348
rect 17957 13339 18015 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 21726 13376 21732 13388
rect 21687 13348 21732 13376
rect 19705 13339 19763 13345
rect 8754 13308 8760 13320
rect 8312 13280 8432 13308
rect 8715 13280 8760 13308
rect 8404 13240 8432 13280
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 9950 13308 9956 13320
rect 9815 13280 9956 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9950 13268 9956 13280
rect 10008 13308 10014 13320
rect 11379 13311 11437 13317
rect 11379 13308 11391 13311
rect 10008 13280 11391 13308
rect 10008 13268 10014 13280
rect 11379 13277 11391 13280
rect 11425 13277 11437 13311
rect 13170 13308 13176 13320
rect 13083 13280 13176 13308
rect 11379 13271 11437 13277
rect 13170 13268 13176 13280
rect 13228 13308 13234 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 13228 13280 13461 13308
rect 13228 13268 13234 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 13449 13271 13507 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 15528 13280 15669 13308
rect 15528 13268 15534 13280
rect 15657 13277 15669 13280
rect 15703 13277 15715 13311
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15657 13271 15715 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 18138 13308 18144 13320
rect 16080 13280 18144 13308
rect 16080 13268 16086 13280
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 19720 13308 19748 13339
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 21928 13385 21956 13416
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 21913 13379 21971 13385
rect 21913 13345 21925 13379
rect 21959 13345 21971 13379
rect 21913 13339 21971 13345
rect 22281 13379 22339 13385
rect 22281 13345 22293 13379
rect 22327 13376 22339 13379
rect 22370 13376 22376 13388
rect 22327 13348 22376 13376
rect 22327 13345 22339 13348
rect 22281 13339 22339 13345
rect 19024 13280 19748 13308
rect 19024 13268 19030 13280
rect 21542 13268 21548 13320
rect 21600 13308 21606 13320
rect 22296 13308 22324 13339
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 22480 13348 22661 13376
rect 21600 13280 22324 13308
rect 21600 13268 21606 13280
rect 9674 13240 9680 13252
rect 8404 13212 9680 13240
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 10321 13243 10379 13249
rect 10321 13209 10333 13243
rect 10367 13209 10379 13243
rect 10321 13203 10379 13209
rect 10336 13172 10364 13203
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 16114 13240 16120 13252
rect 11848 13212 16120 13240
rect 11848 13200 11854 13212
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 22480 13240 22508 13348
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 24118 13376 24124 13388
rect 24079 13348 24124 13376
rect 22649 13339 22707 13345
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 25384 13379 25442 13385
rect 25384 13345 25396 13379
rect 25430 13376 25442 13379
rect 25774 13376 25780 13388
rect 25430 13348 25780 13376
rect 25430 13345 25442 13348
rect 25384 13339 25442 13345
rect 25774 13336 25780 13348
rect 25832 13336 25838 13388
rect 21008 13212 22508 13240
rect 21008 13184 21036 13212
rect 10870 13172 10876 13184
rect 10336 13144 10876 13172
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14550 13172 14556 13184
rect 13872 13144 14556 13172
rect 13872 13132 13878 13144
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 16666 13172 16672 13184
rect 16627 13144 16672 13172
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18874 13172 18880 13184
rect 18196 13144 18880 13172
rect 18196 13132 18202 13144
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 20254 13172 20260 13184
rect 20215 13144 20260 13172
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 20625 13175 20683 13181
rect 20625 13172 20637 13175
rect 20404 13144 20637 13172
rect 20404 13132 20410 13144
rect 20625 13141 20637 13144
rect 20671 13172 20683 13175
rect 20990 13172 20996 13184
rect 20671 13144 20996 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 21726 13132 21732 13184
rect 21784 13172 21790 13184
rect 22462 13172 22468 13184
rect 21784 13144 22468 13172
rect 21784 13132 21790 13144
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 24026 13172 24032 13184
rect 23987 13144 24032 13172
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 9088 12940 9321 12968
rect 9088 12928 9094 12940
rect 9309 12937 9321 12940
rect 9355 12968 9367 12971
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9355 12940 9965 12968
rect 9355 12937 9367 12940
rect 9309 12931 9367 12937
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 9953 12931 10011 12937
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 13872 12940 13917 12968
rect 13872 12928 13878 12940
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14148 12940 14749 12968
rect 14148 12928 14154 12940
rect 14737 12937 14749 12940
rect 14783 12968 14795 12971
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 14783 12940 14841 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 14829 12931 14887 12937
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15804 12940 16037 12968
rect 15804 12928 15810 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 16025 12931 16083 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 7892 12872 12173 12900
rect 7892 12860 7898 12872
rect 12161 12869 12173 12872
rect 12207 12900 12219 12903
rect 12986 12900 12992 12912
rect 12207 12872 12992 12900
rect 12207 12869 12219 12872
rect 12161 12863 12219 12869
rect 12986 12860 12992 12872
rect 13044 12900 13050 12912
rect 13262 12900 13268 12912
rect 13044 12872 13268 12900
rect 13044 12860 13050 12872
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 18417 12903 18475 12909
rect 18417 12900 18429 12903
rect 13786 12872 18429 12900
rect 8294 12832 8300 12844
rect 8207 12804 8300 12832
rect 8294 12792 8300 12804
rect 8352 12832 8358 12844
rect 11238 12832 11244 12844
rect 8352 12804 8753 12832
rect 11199 12804 11244 12832
rect 8352 12792 8358 12804
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 8386 12764 8392 12776
rect 7607 12736 8392 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 6641 12631 6699 12637
rect 6641 12597 6653 12631
rect 6687 12628 6699 12631
rect 6840 12628 6868 12727
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 7392 12696 7420 12727
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 8725 12764 8753 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12832 12955 12835
rect 13170 12832 13176 12844
rect 12943 12804 13176 12832
rect 12943 12801 12955 12804
rect 12897 12795 12955 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 8725 12736 8754 12764
rect 7929 12699 7987 12705
rect 7929 12696 7941 12699
rect 6972 12668 7941 12696
rect 6972 12656 6978 12668
rect 7929 12665 7941 12668
rect 7975 12696 7987 12699
rect 8478 12696 8484 12708
rect 7975 12668 8484 12696
rect 7975 12665 7987 12668
rect 7929 12659 7987 12665
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 8726 12705 8754 12736
rect 8711 12699 8769 12705
rect 8711 12665 8723 12699
rect 8757 12665 8769 12699
rect 10870 12696 10876 12708
rect 10831 12668 10876 12696
rect 8711 12659 8769 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 10965 12699 11023 12705
rect 10965 12665 10977 12699
rect 11011 12665 11023 12699
rect 12802 12696 12808 12708
rect 12715 12668 12808 12696
rect 10965 12659 11023 12665
rect 7834 12628 7840 12640
rect 6687 12600 7840 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 9674 12628 9680 12640
rect 9635 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10689 12631 10747 12637
rect 10689 12597 10701 12631
rect 10735 12628 10747 12631
rect 10980 12628 11008 12659
rect 12802 12656 12808 12668
rect 12860 12696 12866 12708
rect 13259 12699 13317 12705
rect 13259 12696 13271 12699
rect 12860 12668 13271 12696
rect 12860 12656 12866 12668
rect 13259 12665 13271 12668
rect 13305 12696 13317 12699
rect 13630 12696 13636 12708
rect 13305 12668 13636 12696
rect 13305 12665 13317 12668
rect 13259 12659 13317 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 11422 12628 11428 12640
rect 10735 12600 11428 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 11885 12631 11943 12637
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 11974 12628 11980 12640
rect 11931 12600 11980 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 13786 12628 13814 12872
rect 18417 12869 18429 12872
rect 18463 12869 18475 12903
rect 24765 12903 24823 12909
rect 24765 12900 24777 12903
rect 18417 12863 18475 12869
rect 24044 12872 24777 12900
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 15194 12832 15200 12844
rect 15151 12804 15200 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15470 12832 15476 12844
rect 15431 12804 15476 12832
rect 15470 12792 15476 12804
rect 15528 12832 15534 12844
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 15528 12804 16405 12832
rect 15528 12792 15534 12804
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16393 12795 16451 12801
rect 16577 12835 16635 12841
rect 16577 12801 16589 12835
rect 16623 12832 16635 12835
rect 17402 12832 17408 12844
rect 16623 12804 17408 12832
rect 16623 12801 16635 12804
rect 16577 12795 16635 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 18782 12832 18788 12844
rect 18695 12804 18788 12832
rect 18782 12792 18788 12804
rect 18840 12832 18846 12844
rect 20622 12832 20628 12844
rect 18840 12804 20628 12832
rect 18840 12792 18846 12804
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 23845 12835 23903 12841
rect 23845 12801 23857 12835
rect 23891 12832 23903 12835
rect 24044 12832 24072 12872
rect 24765 12869 24777 12872
rect 24811 12900 24823 12903
rect 24811 12872 25360 12900
rect 24811 12869 24823 12872
rect 24765 12863 24823 12869
rect 24210 12832 24216 12844
rect 23891 12804 24072 12832
rect 24171 12804 24216 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 24210 12792 24216 12804
rect 24268 12792 24274 12844
rect 25332 12841 25360 12872
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 17911 12736 18245 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18233 12733 18245 12736
rect 18279 12764 18291 12767
rect 18966 12764 18972 12776
rect 18279 12736 18972 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 19150 12724 19156 12776
rect 19208 12764 19214 12776
rect 19245 12767 19303 12773
rect 19245 12764 19257 12767
rect 19208 12736 19257 12764
rect 19208 12724 19214 12736
rect 19245 12733 19257 12736
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19576 12736 19717 12764
rect 19576 12724 19582 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 20257 12767 20315 12773
rect 20257 12733 20269 12767
rect 20303 12733 20315 12767
rect 20257 12727 20315 12733
rect 15197 12699 15255 12705
rect 15197 12665 15209 12699
rect 15243 12665 15255 12699
rect 15197 12659 15255 12665
rect 12952 12600 13814 12628
rect 14737 12631 14795 12637
rect 12952 12588 12958 12600
rect 14737 12597 14749 12631
rect 14783 12628 14795 12631
rect 15212 12628 15240 12659
rect 14783 12600 15240 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 18932 12600 19073 12628
rect 18932 12588 18938 12600
rect 19061 12597 19073 12600
rect 19107 12597 19119 12631
rect 19334 12628 19340 12640
rect 19295 12600 19340 12628
rect 19061 12591 19119 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 20272 12628 20300 12727
rect 20346 12724 20352 12776
rect 20404 12764 20410 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20404 12736 20453 12764
rect 20404 12724 20410 12736
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 20441 12727 20499 12733
rect 22094 12696 22100 12708
rect 22055 12668 22100 12696
rect 22094 12656 22100 12668
rect 22152 12656 22158 12708
rect 22189 12699 22247 12705
rect 22189 12665 22201 12699
rect 22235 12696 22247 12699
rect 22278 12696 22284 12708
rect 22235 12668 22284 12696
rect 22235 12665 22247 12668
rect 22189 12659 22247 12665
rect 20530 12628 20536 12640
rect 20272 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12628 20594 12640
rect 20993 12631 21051 12637
rect 20993 12628 21005 12631
rect 20588 12600 21005 12628
rect 20588 12588 20594 12600
rect 20993 12597 21005 12600
rect 21039 12628 21051 12631
rect 21453 12631 21511 12637
rect 21453 12628 21465 12631
rect 21039 12600 21465 12628
rect 21039 12597 21051 12600
rect 20993 12591 21051 12597
rect 21453 12597 21465 12600
rect 21499 12628 21511 12631
rect 21542 12628 21548 12640
rect 21499 12600 21548 12628
rect 21499 12597 21511 12600
rect 21453 12591 21511 12597
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 21913 12631 21971 12637
rect 21913 12597 21925 12631
rect 21959 12628 21971 12631
rect 22204 12628 22232 12659
rect 22278 12656 22284 12668
rect 22336 12656 22342 12708
rect 22738 12696 22744 12708
rect 22699 12668 22744 12696
rect 22738 12656 22744 12668
rect 22796 12656 22802 12708
rect 23937 12699 23995 12705
rect 23937 12665 23949 12699
rect 23983 12696 23995 12699
rect 24026 12696 24032 12708
rect 23983 12668 24032 12696
rect 23983 12665 23995 12668
rect 23937 12659 23995 12665
rect 21959 12600 22232 12628
rect 21959 12597 21971 12600
rect 21913 12591 21971 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 22520 12600 23029 12628
rect 22520 12588 22526 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 23017 12591 23075 12597
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 23952 12628 23980 12659
rect 24026 12656 24032 12668
rect 24084 12656 24090 12708
rect 25774 12628 25780 12640
rect 23523 12600 23980 12628
rect 25735 12600 25780 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 25774 12588 25780 12600
rect 25832 12588 25838 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 6914 12424 6920 12436
rect 6875 12396 6920 12424
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8444 12396 9045 12424
rect 8444 12384 8450 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9950 12424 9956 12436
rect 9911 12396 9956 12424
rect 9033 12387 9091 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10192 12396 10241 12424
rect 10192 12384 10198 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 11422 12424 11428 12436
rect 11383 12396 11428 12424
rect 10229 12387 10287 12393
rect 10244 12356 10272 12387
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 13906 12424 13912 12436
rect 13867 12396 13912 12424
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 15194 12424 15200 12436
rect 15151 12396 15200 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 16209 12427 16267 12433
rect 16209 12424 16221 12427
rect 15804 12396 16221 12424
rect 15804 12384 15810 12396
rect 16209 12393 16221 12396
rect 16255 12393 16267 12427
rect 16209 12387 16267 12393
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 17957 12427 18015 12433
rect 17957 12424 17969 12427
rect 16724 12396 17969 12424
rect 16724 12384 16730 12396
rect 17957 12393 17969 12396
rect 18003 12393 18015 12427
rect 17957 12387 18015 12393
rect 18785 12427 18843 12433
rect 18785 12393 18797 12427
rect 18831 12424 18843 12427
rect 19150 12424 19156 12436
rect 18831 12396 19156 12424
rect 18831 12393 18843 12396
rect 18785 12387 18843 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22925 12427 22983 12433
rect 22925 12424 22937 12427
rect 22152 12396 22937 12424
rect 22152 12384 22158 12396
rect 22925 12393 22937 12396
rect 22971 12393 22983 12427
rect 22925 12387 22983 12393
rect 24029 12427 24087 12433
rect 24029 12393 24041 12427
rect 24075 12424 24087 12427
rect 24118 12424 24124 12436
rect 24075 12396 24124 12424
rect 24075 12393 24087 12396
rect 24029 12387 24087 12393
rect 24118 12384 24124 12396
rect 24176 12424 24182 12436
rect 24305 12427 24363 12433
rect 24305 12424 24317 12427
rect 24176 12396 24317 12424
rect 24176 12384 24182 12396
rect 24305 12393 24317 12396
rect 24351 12393 24363 12427
rect 24305 12387 24363 12393
rect 10826 12359 10884 12365
rect 10826 12356 10838 12359
rect 10244 12328 10838 12356
rect 10826 12325 10838 12328
rect 10872 12325 10884 12359
rect 10826 12319 10884 12325
rect 13351 12359 13409 12365
rect 13351 12325 13363 12359
rect 13397 12356 13409 12359
rect 13630 12356 13636 12368
rect 13397 12328 13636 12356
rect 13397 12325 13409 12328
rect 13351 12319 13409 12325
rect 13630 12316 13636 12328
rect 13688 12356 13694 12368
rect 15651 12359 15709 12365
rect 15651 12356 15663 12359
rect 13688 12328 15663 12356
rect 13688 12316 13694 12328
rect 15651 12325 15663 12328
rect 15697 12356 15709 12359
rect 15930 12356 15936 12368
rect 15697 12328 15936 12356
rect 15697 12325 15709 12328
rect 15651 12319 15709 12325
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 17310 12356 17316 12368
rect 17271 12328 17316 12356
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 18417 12359 18475 12365
rect 18417 12325 18429 12359
rect 18463 12356 18475 12359
rect 18463 12328 19564 12356
rect 18463 12325 18475 12328
rect 18417 12319 18475 12325
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8478 12288 8484 12300
rect 8439 12260 8484 12288
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 8812 12260 10517 12288
rect 8812 12248 8818 12260
rect 10505 12257 10517 12260
rect 10551 12288 10563 12291
rect 10686 12288 10692 12300
rect 10551 12260 10692 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 11940 12260 17442 12288
rect 11940 12248 11946 12260
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 14516 12192 15301 12220
rect 14516 12180 14522 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 17034 12220 17040 12232
rect 16995 12192 17040 12220
rect 15289 12183 15347 12189
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 17414 12220 17442 12260
rect 19058 12248 19064 12300
rect 19116 12288 19122 12300
rect 19536 12297 19564 12328
rect 20622 12316 20628 12368
rect 20680 12356 20686 12368
rect 21723 12359 21781 12365
rect 21723 12356 21735 12359
rect 20680 12328 21735 12356
rect 20680 12316 20686 12328
rect 21723 12325 21735 12328
rect 21769 12356 21781 12359
rect 21910 12356 21916 12368
rect 21769 12328 21916 12356
rect 21769 12325 21781 12328
rect 21723 12319 21781 12325
rect 21910 12316 21916 12328
rect 21968 12356 21974 12368
rect 23014 12356 23020 12368
rect 21968 12328 23020 12356
rect 21968 12316 21974 12328
rect 23014 12316 23020 12328
rect 23072 12356 23078 12368
rect 23430 12359 23488 12365
rect 23430 12356 23442 12359
rect 23072 12328 23442 12356
rect 23072 12316 23078 12328
rect 23430 12325 23442 12328
rect 23476 12325 23488 12359
rect 24762 12356 24768 12368
rect 23430 12319 23488 12325
rect 24596 12328 24768 12356
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19116 12260 19257 12288
rect 19116 12248 19122 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19521 12291 19579 12297
rect 19521 12257 19533 12291
rect 19567 12288 19579 12291
rect 20162 12288 20168 12300
rect 19567 12260 20168 12288
rect 19567 12257 19579 12260
rect 19521 12251 19579 12257
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12288 22339 12291
rect 22646 12288 22652 12300
rect 22327 12260 22652 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 22646 12248 22652 12260
rect 22704 12288 22710 12300
rect 24596 12288 24624 12328
rect 24762 12316 24768 12328
rect 24820 12356 24826 12368
rect 25041 12359 25099 12365
rect 25041 12356 25053 12359
rect 24820 12328 25053 12356
rect 24820 12316 24826 12328
rect 25041 12325 25053 12328
rect 25087 12325 25099 12359
rect 25041 12319 25099 12325
rect 22704 12260 24624 12288
rect 22704 12248 22710 12260
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 17414 12192 19717 12220
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 19705 12183 19763 12189
rect 20088 12192 21097 12220
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15838 12152 15844 12164
rect 15252 12124 15844 12152
rect 15252 12112 15258 12124
rect 15838 12112 15844 12124
rect 15896 12112 15902 12164
rect 19337 12155 19395 12161
rect 19337 12121 19349 12155
rect 19383 12152 19395 12155
rect 19518 12152 19524 12164
rect 19383 12124 19524 12152
rect 19383 12121 19395 12124
rect 19337 12115 19395 12121
rect 19518 12112 19524 12124
rect 19576 12152 19582 12164
rect 20088 12152 20116 12192
rect 21085 12189 21097 12192
rect 21131 12220 21143 12223
rect 21174 12220 21180 12232
rect 21131 12192 21180 12220
rect 21131 12189 21143 12192
rect 21085 12183 21143 12189
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 21358 12220 21364 12232
rect 21319 12192 21364 12220
rect 21358 12180 21364 12192
rect 21416 12220 21422 12232
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 21416 12192 22569 12220
rect 21416 12180 21422 12192
rect 22557 12189 22569 12192
rect 22603 12189 22615 12223
rect 22557 12183 22615 12189
rect 23014 12180 23020 12232
rect 23072 12220 23078 12232
rect 23109 12223 23167 12229
rect 23109 12220 23121 12223
rect 23072 12192 23121 12220
rect 23072 12180 23078 12192
rect 23109 12189 23121 12192
rect 23155 12189 23167 12223
rect 23109 12183 23167 12189
rect 24670 12180 24676 12232
rect 24728 12220 24734 12232
rect 24949 12223 25007 12229
rect 24949 12220 24961 12223
rect 24728 12192 24961 12220
rect 24728 12180 24734 12192
rect 24949 12189 24961 12192
rect 24995 12189 25007 12223
rect 25225 12223 25283 12229
rect 25225 12220 25237 12223
rect 24949 12183 25007 12189
rect 25056 12192 25237 12220
rect 19576 12124 20116 12152
rect 19576 12112 19582 12124
rect 20254 12112 20260 12164
rect 20312 12152 20318 12164
rect 20717 12155 20775 12161
rect 20717 12152 20729 12155
rect 20312 12124 20729 12152
rect 20312 12112 20318 12124
rect 20717 12121 20729 12124
rect 20763 12152 20775 12155
rect 22002 12152 22008 12164
rect 20763 12124 22008 12152
rect 20763 12121 20775 12124
rect 20717 12115 20775 12121
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 23750 12112 23756 12164
rect 23808 12152 23814 12164
rect 24765 12155 24823 12161
rect 24765 12152 24777 12155
rect 23808 12124 24777 12152
rect 23808 12112 23814 12124
rect 24765 12121 24777 12124
rect 24811 12152 24823 12155
rect 25056 12152 25084 12192
rect 25225 12189 25237 12192
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 24811 12124 25084 12152
rect 24811 12121 24823 12124
rect 24765 12115 24823 12121
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12894 12084 12900 12096
rect 12575 12056 12900 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 19061 12087 19119 12093
rect 19061 12084 19073 12087
rect 18748 12056 19073 12084
rect 18748 12044 18754 12056
rect 19061 12053 19073 12056
rect 19107 12084 19119 12087
rect 20346 12084 20352 12096
rect 19107 12056 20352 12084
rect 19107 12053 19119 12056
rect 19061 12047 19119 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 7653 11883 7711 11889
rect 7653 11849 7665 11883
rect 7699 11880 7711 11883
rect 8478 11880 8484 11892
rect 7699 11852 8484 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 10134 11880 10140 11892
rect 8817 11852 10140 11880
rect 8294 11812 8300 11824
rect 8255 11784 8300 11812
rect 8294 11772 8300 11784
rect 8352 11772 8358 11824
rect 8312 11676 8340 11772
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8570 11744 8576 11756
rect 8527 11716 8576 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 8817 11676 8845 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 12802 11880 12808 11892
rect 12763 11852 12808 11880
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13909 11883 13967 11889
rect 13909 11849 13921 11883
rect 13955 11880 13967 11883
rect 14090 11880 14096 11892
rect 13955 11852 14096 11880
rect 13955 11849 13967 11852
rect 13909 11843 13967 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 14608 11852 14749 11880
rect 14608 11840 14614 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 14737 11843 14795 11849
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 10100 11784 11161 11812
rect 10100 11772 10106 11784
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11149 11775 11207 11781
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 8312 11648 8845 11676
rect 7466 11568 7472 11620
rect 7524 11608 7530 11620
rect 8817 11617 8845 11648
rect 9692 11648 10241 11676
rect 8802 11611 8860 11617
rect 7524 11580 8569 11608
rect 7524 11568 7530 11580
rect 8018 11540 8024 11552
rect 7979 11512 8024 11540
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 8541 11540 8569 11580
rect 8802 11577 8814 11611
rect 8848 11577 8860 11611
rect 8802 11571 8860 11577
rect 9214 11540 9220 11552
rect 8541 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11540 9278 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9272 11512 9413 11540
rect 9272 11500 9278 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9692 11549 9720 11648
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12989 11679 13047 11685
rect 12989 11676 13001 11679
rect 12299 11648 13001 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 12989 11645 13001 11648
rect 13035 11676 13047 11679
rect 13722 11676 13728 11688
rect 13035 11648 13728 11676
rect 13035 11645 13047 11648
rect 12989 11639 13047 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 10134 11568 10140 11620
rect 10192 11608 10198 11620
rect 10550 11611 10608 11617
rect 10550 11608 10562 11611
rect 10192 11580 10562 11608
rect 10192 11568 10198 11580
rect 10550 11577 10562 11580
rect 10596 11577 10608 11611
rect 10550 11571 10608 11577
rect 12802 11568 12808 11620
rect 12860 11608 12866 11620
rect 13310 11611 13368 11617
rect 13310 11608 13322 11611
rect 12860 11580 13322 11608
rect 12860 11568 12866 11580
rect 13310 11577 13322 11580
rect 13356 11577 13368 11611
rect 14752 11608 14780 11843
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17092 11852 17785 11880
rect 17092 11840 17098 11852
rect 17773 11849 17785 11852
rect 17819 11880 17831 11883
rect 19334 11880 19340 11892
rect 17819 11852 19340 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19751 11883 19809 11889
rect 19751 11849 19763 11883
rect 19797 11880 19809 11883
rect 19797 11852 23474 11880
rect 19797 11849 19809 11852
rect 19751 11843 19809 11849
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 15565 11815 15623 11821
rect 15565 11812 15577 11815
rect 15528 11784 15577 11812
rect 15528 11772 15534 11784
rect 15565 11781 15577 11784
rect 15611 11781 15623 11815
rect 15565 11775 15623 11781
rect 15930 11772 15936 11824
rect 15988 11812 15994 11824
rect 16025 11815 16083 11821
rect 16025 11812 16037 11815
rect 15988 11784 16037 11812
rect 15988 11772 15994 11784
rect 16025 11781 16037 11784
rect 16071 11812 16083 11815
rect 17310 11812 17316 11824
rect 16071 11784 17316 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 17310 11772 17316 11784
rect 17368 11812 17374 11824
rect 20622 11812 20628 11824
rect 17368 11784 17448 11812
rect 20583 11784 20628 11812
rect 17368 11772 17374 11784
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 15059 11716 16313 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 16301 11713 16313 11716
rect 16347 11744 16359 11747
rect 16623 11747 16681 11753
rect 16623 11744 16635 11747
rect 16347 11716 16635 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16623 11713 16635 11716
rect 16669 11713 16681 11747
rect 16623 11707 16681 11713
rect 16536 11679 16594 11685
rect 16536 11645 16548 11679
rect 16582 11676 16594 11679
rect 16582 11648 17080 11676
rect 16582 11645 16594 11648
rect 16536 11639 16594 11645
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 14752 11580 15117 11608
rect 13310 11571 13368 11577
rect 15105 11577 15117 11580
rect 15151 11577 15163 11611
rect 15105 11571 15163 11577
rect 17052 11552 17080 11648
rect 17420 11617 17448 11784
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 23446 11812 23474 11852
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 24857 11883 24915 11889
rect 24857 11880 24869 11883
rect 24820 11852 24869 11880
rect 24820 11840 24826 11852
rect 24857 11849 24869 11852
rect 24903 11849 24915 11883
rect 24857 11843 24915 11849
rect 24670 11812 24676 11824
rect 23446 11784 24676 11812
rect 24670 11772 24676 11784
rect 24728 11812 24734 11824
rect 25685 11815 25743 11821
rect 25685 11812 25697 11815
rect 24728 11784 25697 11812
rect 24728 11772 24734 11784
rect 25685 11781 25697 11784
rect 25731 11781 25743 11815
rect 25685 11775 25743 11781
rect 18046 11744 18052 11756
rect 18007 11716 18052 11744
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19518 11744 19524 11756
rect 19383 11716 19524 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 22738 11704 22744 11756
rect 22796 11744 22802 11756
rect 23750 11744 23756 11756
rect 22796 11716 23756 11744
rect 22796 11704 22802 11716
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 24210 11744 24216 11756
rect 24171 11716 24216 11744
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 18138 11676 18144 11688
rect 18099 11648 18144 11676
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 19648 11679 19706 11685
rect 19648 11676 19660 11679
rect 18656 11648 19660 11676
rect 18656 11636 18662 11648
rect 19648 11645 19660 11648
rect 19694 11676 19706 11679
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19694 11648 20085 11676
rect 19694 11645 19706 11648
rect 19648 11639 19706 11645
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20898 11676 20904 11688
rect 20859 11648 20904 11676
rect 20073 11639 20131 11645
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 21174 11676 21180 11688
rect 21135 11648 21180 11676
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 21729 11679 21787 11685
rect 21729 11645 21741 11679
rect 21775 11645 21787 11679
rect 22002 11676 22008 11688
rect 21963 11648 22008 11676
rect 21729 11639 21787 11645
rect 17405 11611 17463 11617
rect 17405 11577 17417 11611
rect 17451 11608 17463 11611
rect 18782 11608 18788 11620
rect 17451 11580 18788 11608
rect 17451 11577 17463 11580
rect 17405 11571 17463 11577
rect 18782 11568 18788 11580
rect 18840 11568 18846 11620
rect 21744 11552 21772 11639
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 22189 11611 22247 11617
rect 22189 11577 22201 11611
rect 22235 11608 22247 11611
rect 23014 11608 23020 11620
rect 22235 11580 23020 11608
rect 22235 11577 22247 11580
rect 22189 11571 22247 11577
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 23845 11611 23903 11617
rect 23845 11577 23857 11611
rect 23891 11608 23903 11611
rect 24118 11608 24124 11620
rect 23891 11580 24124 11608
rect 23891 11577 23903 11580
rect 23845 11571 23903 11577
rect 24118 11568 24124 11580
rect 24176 11568 24182 11620
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9640 11512 9689 11540
rect 9640 11500 9646 11512
rect 9677 11509 9689 11512
rect 9723 11509 9735 11543
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 9677 11503 9735 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 17034 11540 17040 11552
rect 16995 11512 17040 11540
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 22465 11543 22523 11549
rect 22465 11540 22477 11543
rect 21784 11512 22477 11540
rect 21784 11500 21790 11512
rect 22465 11509 22477 11512
rect 22511 11509 22523 11543
rect 22465 11503 22523 11509
rect 22922 11500 22928 11552
rect 22980 11540 22986 11552
rect 23109 11543 23167 11549
rect 23109 11540 23121 11543
rect 22980 11512 23121 11540
rect 22980 11500 22986 11512
rect 23109 11509 23121 11512
rect 23155 11509 23167 11543
rect 25222 11540 25228 11552
rect 25183 11512 25228 11540
rect 23109 11503 23167 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 9033 11339 9091 11345
rect 9033 11336 9045 11339
rect 8628 11308 9045 11336
rect 8628 11296 8634 11308
rect 9033 11305 9045 11308
rect 9079 11305 9091 11339
rect 10686 11336 10692 11348
rect 10647 11308 10692 11336
rect 9033 11299 9091 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12802 11336 12808 11348
rect 12400 11308 12808 11336
rect 12400 11296 12406 11308
rect 12802 11296 12808 11308
rect 12860 11336 12866 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12860 11308 13093 11336
rect 12860 11296 12866 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13722 11336 13728 11348
rect 13683 11308 13728 11336
rect 13081 11299 13139 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 17589 11339 17647 11345
rect 13964 11308 15516 11336
rect 13964 11296 13970 11308
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 9582 11268 9588 11280
rect 8803 11240 9588 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 9861 11271 9919 11277
rect 9861 11237 9873 11271
rect 9907 11268 9919 11271
rect 10042 11268 10048 11280
rect 9907 11240 10048 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 12161 11271 12219 11277
rect 12161 11268 12173 11271
rect 10836 11240 12173 11268
rect 10836 11228 10842 11240
rect 12161 11237 12173 11240
rect 12207 11237 12219 11271
rect 12161 11231 12219 11237
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 15488 11277 15516 11308
rect 17589 11305 17601 11339
rect 17635 11336 17647 11339
rect 18138 11336 18144 11348
rect 17635 11308 18144 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 19058 11336 19064 11348
rect 19019 11308 19064 11336
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21358 11336 21364 11348
rect 21223 11308 21364 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 22646 11336 22652 11348
rect 22607 11308 22652 11336
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 23014 11336 23020 11348
rect 22975 11308 23020 11336
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 24213 11339 24271 11345
rect 24213 11336 24225 11339
rect 24176 11308 24225 11336
rect 24176 11296 24182 11308
rect 24213 11305 24225 11308
rect 24259 11305 24271 11339
rect 24213 11299 24271 11305
rect 24903 11339 24961 11345
rect 24903 11305 24915 11339
rect 24949 11336 24961 11339
rect 25038 11336 25044 11348
rect 24949 11308 25044 11336
rect 24949 11305 24961 11308
rect 24903 11299 24961 11305
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 15473 11271 15531 11277
rect 12308 11240 12353 11268
rect 12308 11228 12314 11240
rect 15473 11237 15485 11271
rect 15519 11268 15531 11271
rect 15746 11268 15752 11280
rect 15519 11240 15752 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 17862 11268 17868 11280
rect 17823 11240 17868 11268
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 20346 11228 20352 11280
rect 20404 11268 20410 11280
rect 20404 11240 22140 11268
rect 20404 11228 20410 11240
rect 7006 11200 7012 11212
rect 6967 11172 7012 11200
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7984 11172 8033 11200
rect 7984 11160 7990 11172
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 8536 11172 8585 11200
rect 8536 11160 8542 11172
rect 8573 11169 8585 11172
rect 8619 11200 8631 11203
rect 9398 11200 9404 11212
rect 8619 11172 9404 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13964 11172 14105 11200
rect 13964 11160 13970 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 18969 11203 19027 11209
rect 18969 11169 18981 11203
rect 19015 11200 19027 11203
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 19015 11172 19257 11200
rect 19015 11169 19027 11172
rect 18969 11163 19027 11169
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 19392 11172 19717 11200
rect 19392 11160 19398 11172
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 20898 11200 20904 11212
rect 20763 11172 20904 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 21174 11160 21180 11212
rect 21232 11200 21238 11212
rect 21361 11203 21419 11209
rect 21361 11200 21373 11203
rect 21232 11172 21373 11200
rect 21232 11160 21238 11172
rect 21361 11169 21373 11172
rect 21407 11169 21419 11203
rect 21726 11200 21732 11212
rect 21687 11172 21732 11200
rect 21361 11163 21419 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 22112 11209 22140 11240
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11169 22155 11203
rect 22097 11163 22155 11169
rect 23198 11160 23204 11212
rect 23256 11200 23262 11212
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 23256 11172 23305 11200
rect 23256 11160 23262 11172
rect 23293 11169 23305 11172
rect 23339 11169 23351 11203
rect 23293 11163 23351 11169
rect 24832 11203 24890 11209
rect 24832 11169 24844 11203
rect 24878 11200 24890 11203
rect 25130 11200 25136 11212
rect 24878 11172 25136 11200
rect 24878 11169 24890 11172
rect 24832 11163 24890 11169
rect 25130 11160 25136 11172
rect 25188 11160 25194 11212
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9416 11104 9781 11132
rect 7193 10999 7251 11005
rect 7193 10965 7205 10999
rect 7239 10996 7251 10999
rect 8570 10996 8576 11008
rect 7239 10968 8576 10996
rect 7239 10965 7251 10968
rect 7193 10959 7251 10965
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9416 11005 9444 11104
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 10226 11132 10232 11144
rect 10187 11104 10232 11132
rect 9769 11095 9827 11101
rect 10226 11092 10232 11104
rect 10284 11132 10290 11144
rect 10870 11132 10876 11144
rect 10284 11104 10876 11132
rect 10284 11092 10290 11104
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 12802 11132 12808 11144
rect 12763 11104 12808 11132
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 15028 11104 15393 11132
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 12986 11064 12992 11076
rect 11480 11036 12992 11064
rect 11480 11024 11486 11036
rect 12986 11024 12992 11036
rect 13044 11064 13050 11076
rect 13449 11067 13507 11073
rect 13449 11064 13461 11067
rect 13044 11036 13461 11064
rect 13044 11024 13050 11036
rect 13449 11033 13461 11036
rect 13495 11033 13507 11067
rect 13449 11027 13507 11033
rect 9401 10999 9459 11005
rect 9401 10996 9413 10999
rect 9364 10968 9413 10996
rect 9364 10956 9370 10968
rect 9401 10965 9413 10968
rect 9447 10965 9459 10999
rect 9401 10959 9459 10965
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 15028 11005 15056 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 15528 11104 15669 11132
rect 15528 11092 15534 11104
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 17368 11104 17785 11132
rect 17368 11092 17374 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 19797 11135 19855 11141
rect 19797 11132 19809 11135
rect 17773 11095 17831 11101
rect 17972 11104 19809 11132
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 17972 11064 18000 11104
rect 19797 11101 19809 11104
rect 19843 11101 19855 11135
rect 19797 11095 19855 11101
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11132 23995 11135
rect 24210 11132 24216 11144
rect 23983 11104 24216 11132
rect 23983 11101 23995 11104
rect 23937 11095 23995 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 18322 11064 18328 11076
rect 15620 11036 18000 11064
rect 18283 11036 18328 11064
rect 15620 11024 15626 11036
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 15013 10999 15071 11005
rect 15013 10996 15025 10999
rect 14700 10968 15025 10996
rect 14700 10956 14706 10968
rect 15013 10965 15025 10968
rect 15059 10965 15071 10999
rect 15013 10959 15071 10965
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 16264 10968 16313 10996
rect 16264 10956 16270 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 16301 10959 16359 10965
rect 17221 10999 17279 11005
rect 17221 10965 17233 10999
rect 17267 10996 17279 10999
rect 17310 10996 17316 11008
rect 17267 10968 17316 10996
rect 17267 10965 17279 10968
rect 17221 10959 17279 10965
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 17494 10956 17500 11008
rect 17552 10996 17558 11008
rect 17678 10996 17684 11008
rect 17552 10968 17684 10996
rect 17552 10956 17558 10968
rect 17678 10956 17684 10968
rect 17736 10996 17742 11008
rect 18693 10999 18751 11005
rect 18693 10996 18705 10999
rect 17736 10968 18705 10996
rect 17736 10956 17742 10968
rect 18693 10965 18705 10968
rect 18739 10996 18751 10999
rect 18969 10999 19027 11005
rect 18969 10996 18981 10999
rect 18739 10968 18981 10996
rect 18739 10965 18751 10968
rect 18693 10959 18751 10965
rect 18969 10965 18981 10968
rect 19015 10965 19027 10999
rect 24670 10996 24676 11008
rect 24631 10968 24676 10996
rect 18969 10959 19027 10965
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 7006 10792 7012 10804
rect 6687 10764 7012 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 9398 10792 9404 10804
rect 9359 10764 9404 10792
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10100 10764 10609 10792
rect 10100 10752 10106 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 10836 10764 11161 10792
rect 10836 10752 10842 10764
rect 11149 10761 11161 10764
rect 11195 10761 11207 10795
rect 12250 10792 12256 10804
rect 12211 10764 12256 10792
rect 11149 10755 11207 10761
rect 12250 10752 12256 10764
rect 12308 10792 12314 10804
rect 13630 10792 13636 10804
rect 12308 10764 13636 10792
rect 12308 10752 12314 10764
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 15746 10792 15752 10804
rect 15707 10764 15752 10792
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 20993 10795 21051 10801
rect 18932 10764 19564 10792
rect 18932 10752 18938 10764
rect 19536 10736 19564 10764
rect 20993 10761 21005 10795
rect 21039 10792 21051 10795
rect 21174 10792 21180 10804
rect 21039 10764 21180 10792
rect 21039 10761 21051 10764
rect 20993 10755 21051 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 22278 10792 22284 10804
rect 22239 10764 22284 10792
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 8036 10696 9045 10724
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 6604 10628 7849 10656
rect 6604 10616 6610 10628
rect 7837 10625 7849 10628
rect 7883 10656 7895 10659
rect 7926 10656 7932 10668
rect 7883 10628 7932 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 7926 10616 7932 10628
rect 7984 10656 7990 10668
rect 8036 10656 8064 10696
rect 9033 10693 9045 10696
rect 9079 10724 9091 10727
rect 9950 10724 9956 10736
rect 9079 10696 9956 10724
rect 9079 10693 9091 10696
rect 9033 10687 9091 10693
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 10226 10724 10232 10736
rect 10187 10696 10232 10724
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 12434 10724 12440 10736
rect 10744 10696 12440 10724
rect 10744 10684 10750 10696
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 13262 10684 13268 10736
rect 13320 10724 13326 10736
rect 15565 10727 15623 10733
rect 15565 10724 15577 10727
rect 13320 10696 15577 10724
rect 13320 10684 13326 10696
rect 15565 10693 15577 10696
rect 15611 10693 15623 10727
rect 15565 10687 15623 10693
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 17862 10724 17868 10736
rect 17543 10696 17868 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 17862 10684 17868 10696
rect 17920 10724 17926 10736
rect 18969 10727 19027 10733
rect 18969 10724 18981 10727
rect 17920 10696 18981 10724
rect 17920 10684 17926 10696
rect 18969 10693 18981 10696
rect 19015 10693 19027 10727
rect 18969 10687 19027 10693
rect 19518 10684 19524 10736
rect 19576 10724 19582 10736
rect 19889 10727 19947 10733
rect 19889 10724 19901 10727
rect 19576 10696 19901 10724
rect 19576 10684 19582 10696
rect 19889 10693 19901 10696
rect 19935 10693 19947 10727
rect 19889 10687 19947 10693
rect 20898 10684 20904 10736
rect 20956 10724 20962 10736
rect 21637 10727 21695 10733
rect 21637 10724 21649 10727
rect 20956 10696 21649 10724
rect 20956 10684 20962 10696
rect 21637 10693 21649 10696
rect 21683 10693 21695 10727
rect 21637 10687 21695 10693
rect 7984 10628 8064 10656
rect 7984 10616 7990 10628
rect 8036 10597 8064 10628
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10656 8815 10659
rect 11514 10656 11520 10668
rect 8803 10628 11520 10656
rect 8803 10625 8815 10628
rect 8757 10619 8815 10625
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12526 10656 12532 10668
rect 12124 10628 12532 10656
rect 12124 10616 12130 10628
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 13906 10656 13912 10668
rect 13412 10628 13912 10656
rect 13412 10616 13418 10628
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 20257 10659 20315 10665
rect 20257 10656 20269 10659
rect 14608 10628 20269 10656
rect 14608 10616 14614 10628
rect 20257 10625 20269 10628
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 24305 10659 24363 10665
rect 24305 10656 24317 10659
rect 23532 10628 24317 10656
rect 23532 10616 23538 10628
rect 24305 10625 24317 10628
rect 24351 10656 24363 10659
rect 24670 10656 24676 10668
rect 24351 10628 24676 10656
rect 24351 10625 24363 10628
rect 24305 10619 24363 10625
rect 24670 10616 24676 10628
rect 24728 10616 24734 10668
rect 24946 10656 24952 10668
rect 24907 10628 24952 10656
rect 24946 10616 24952 10628
rect 25004 10616 25010 10668
rect 7044 10591 7102 10597
rect 7044 10557 7056 10591
rect 7090 10557 7102 10591
rect 7044 10551 7102 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10557 8079 10591
rect 8570 10588 8576 10600
rect 8531 10560 8576 10588
rect 8021 10551 8079 10557
rect 7059 10452 7087 10551
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11368 10591 11426 10597
rect 11368 10588 11380 10591
rect 11296 10560 11380 10588
rect 11296 10548 11302 10560
rect 11368 10557 11380 10560
rect 11414 10588 11426 10591
rect 11790 10588 11796 10600
rect 11414 10560 11796 10588
rect 11414 10557 11426 10560
rect 11368 10551 11426 10557
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14139 10560 14657 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14645 10557 14657 10560
rect 14691 10588 14703 10591
rect 14737 10591 14795 10597
rect 14737 10588 14749 10591
rect 14691 10560 14749 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 14737 10557 14749 10560
rect 14783 10557 14795 10591
rect 14737 10551 14795 10557
rect 7147 10523 7205 10529
rect 7147 10489 7159 10523
rect 7193 10520 7205 10523
rect 9490 10520 9496 10532
rect 7193 10492 9496 10520
rect 7193 10489 7205 10492
rect 7147 10483 7205 10489
rect 9490 10480 9496 10492
rect 9548 10520 9554 10532
rect 9677 10523 9735 10529
rect 9677 10520 9689 10523
rect 9548 10492 9689 10520
rect 9548 10480 9554 10492
rect 9677 10489 9689 10492
rect 9723 10489 9735 10523
rect 9677 10483 9735 10489
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10489 9827 10523
rect 9769 10483 9827 10489
rect 11471 10523 11529 10529
rect 11471 10489 11483 10523
rect 11517 10520 11529 10523
rect 12342 10520 12348 10532
rect 11517 10492 12348 10520
rect 11517 10489 11529 10492
rect 11471 10483 11529 10489
rect 7558 10452 7564 10464
rect 7059 10424 7564 10452
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9784 10452 9812 10483
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 12676 10492 12721 10520
rect 12676 10480 12682 10492
rect 12894 10480 12900 10532
rect 12952 10520 12958 10532
rect 13722 10520 13728 10532
rect 12952 10492 13728 10520
rect 12952 10480 12958 10492
rect 13722 10480 13728 10492
rect 13780 10520 13786 10532
rect 14108 10520 14136 10551
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 14884 10560 15209 10588
rect 14884 10548 14890 10560
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 13780 10492 14136 10520
rect 15565 10523 15623 10529
rect 13780 10480 13786 10492
rect 15565 10489 15577 10523
rect 15611 10520 15623 10523
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 15611 10492 16221 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 16209 10489 16221 10492
rect 16255 10520 16267 10523
rect 16316 10520 16344 10551
rect 16390 10548 16396 10600
rect 16448 10588 16454 10600
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 16448 10560 16773 10588
rect 16448 10548 16454 10560
rect 16761 10557 16773 10560
rect 16807 10588 16819 10591
rect 17770 10588 17776 10600
rect 16807 10560 17776 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 20073 10591 20131 10597
rect 20073 10557 20085 10591
rect 20119 10588 20131 10591
rect 20162 10588 20168 10600
rect 20119 10560 20168 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 16482 10520 16488 10532
rect 16255 10492 16488 10520
rect 16255 10489 16267 10492
rect 16209 10483 16267 10489
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 17865 10523 17923 10529
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18411 10523 18469 10529
rect 18411 10520 18423 10523
rect 17911 10492 18423 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 18411 10489 18423 10492
rect 18457 10520 18469 10523
rect 18782 10520 18788 10532
rect 18457 10492 18788 10520
rect 18457 10489 18469 10492
rect 18411 10483 18469 10489
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 19812 10520 19840 10551
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 22646 10588 22652 10600
rect 22607 10560 22652 10588
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 24397 10523 24455 10529
rect 19812 10492 20116 10520
rect 20088 10464 20116 10492
rect 24397 10489 24409 10523
rect 24443 10489 24455 10523
rect 24397 10483 24455 10489
rect 9858 10452 9864 10464
rect 9272 10424 9864 10452
rect 9272 10412 9278 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 13412 10424 13645 10452
rect 13412 10412 13418 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 13633 10415 13691 10421
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14516 10424 14841 10452
rect 14516 10412 14522 10424
rect 14829 10421 14841 10424
rect 14875 10421 14887 10455
rect 14829 10415 14887 10421
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 16393 10455 16451 10461
rect 16393 10452 16405 10455
rect 16356 10424 16405 10452
rect 16356 10412 16362 10424
rect 16393 10421 16405 10424
rect 16439 10421 16451 10455
rect 16393 10415 16451 10421
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 19242 10452 19248 10464
rect 17828 10424 19248 10452
rect 17828 10412 17834 10424
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19576 10424 19625 10452
rect 19576 10412 19582 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 19613 10415 19671 10421
rect 20070 10412 20076 10464
rect 20128 10452 20134 10464
rect 21269 10455 21327 10461
rect 21269 10452 21281 10455
rect 20128 10424 21281 10452
rect 20128 10412 20134 10424
rect 21269 10421 21281 10424
rect 21315 10452 21327 10455
rect 21726 10452 21732 10464
rect 21315 10424 21732 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 23198 10452 23204 10464
rect 23159 10424 23204 10452
rect 23198 10412 23204 10424
rect 23256 10412 23262 10464
rect 24121 10455 24179 10461
rect 24121 10421 24133 10455
rect 24167 10452 24179 10455
rect 24412 10452 24440 10483
rect 24854 10452 24860 10464
rect 24167 10424 24860 10452
rect 24167 10421 24179 10424
rect 24121 10415 24179 10421
rect 24854 10412 24860 10424
rect 24912 10412 24918 10464
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 25225 10455 25283 10461
rect 25225 10452 25237 10455
rect 25188 10424 25237 10452
rect 25188 10412 25194 10424
rect 25225 10421 25237 10424
rect 25271 10421 25283 10455
rect 25225 10415 25283 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 7147 10251 7205 10257
rect 7147 10217 7159 10251
rect 7193 10248 7205 10251
rect 9306 10248 9312 10260
rect 7193 10220 9312 10248
rect 7193 10217 7205 10220
rect 7147 10211 7205 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9858 10248 9864 10260
rect 9819 10220 9864 10248
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 11514 10248 11520 10260
rect 11475 10220 11520 10248
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10248 12682 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12676 10220 12909 10248
rect 12676 10208 12682 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 12897 10211 12955 10217
rect 16393 10251 16451 10257
rect 16393 10217 16405 10251
rect 16439 10248 16451 10251
rect 17218 10248 17224 10260
rect 16439 10220 17224 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 17218 10208 17224 10220
rect 17276 10248 17282 10260
rect 17276 10220 17448 10248
rect 17276 10208 17282 10220
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 10873 10183 10931 10189
rect 10008 10152 10640 10180
rect 10008 10140 10014 10152
rect 6064 10115 6122 10121
rect 6064 10081 6076 10115
rect 6110 10112 6122 10115
rect 6638 10112 6644 10124
rect 6110 10084 6644 10112
rect 6110 10081 6122 10084
rect 6064 10075 6122 10081
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7098 10112 7104 10124
rect 7055 10084 7104 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 8018 10112 8024 10124
rect 7979 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8570 10112 8576 10124
rect 8483 10084 8576 10112
rect 8570 10072 8576 10084
rect 8628 10112 8634 10124
rect 9858 10112 9864 10124
rect 8628 10084 9864 10112
rect 8628 10072 8634 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10612 10121 10640 10152
rect 10873 10149 10885 10183
rect 10919 10180 10931 10183
rect 11422 10180 11428 10192
rect 10919 10152 11428 10180
rect 10919 10149 10931 10152
rect 10873 10143 10931 10149
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10112 10655 10115
rect 11146 10112 11152 10124
rect 10643 10084 11152 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 11532 10112 11560 10208
rect 12063 10183 12121 10189
rect 12063 10149 12075 10183
rect 12109 10180 12121 10183
rect 12250 10180 12256 10192
rect 12109 10152 12256 10180
rect 12109 10149 12121 10152
rect 12063 10143 12121 10149
rect 12250 10140 12256 10152
rect 12308 10140 12314 10192
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 13538 10180 13544 10192
rect 12400 10152 13544 10180
rect 12400 10140 12406 10152
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 15835 10183 15893 10189
rect 13688 10152 13733 10180
rect 13688 10140 13694 10152
rect 15835 10149 15847 10183
rect 15881 10180 15893 10183
rect 15930 10180 15936 10192
rect 15881 10152 15936 10180
rect 15881 10149 15893 10152
rect 15835 10143 15893 10149
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 17310 10180 17316 10192
rect 16132 10152 17316 10180
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 11532 10084 11713 10112
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12584 10084 13277 10112
rect 12584 10072 12590 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 15473 10115 15531 10121
rect 15473 10081 15485 10115
rect 15519 10112 15531 10115
rect 15562 10112 15568 10124
rect 15519 10084 15568 10112
rect 15519 10081 15531 10084
rect 15473 10075 15531 10081
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8588 10044 8616 10072
rect 7975 10016 8616 10044
rect 8757 10047 8815 10053
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 12434 10044 12440 10056
rect 8803 10016 12440 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 16132 10044 16160 10152
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 17420 10189 17448 10220
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18104 10220 18337 10248
rect 18104 10208 18110 10220
rect 18325 10217 18337 10220
rect 18371 10248 18383 10251
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18371 10220 18889 10248
rect 18371 10217 18383 10220
rect 18325 10211 18383 10217
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 18877 10211 18935 10217
rect 18966 10208 18972 10260
rect 19024 10248 19030 10260
rect 21361 10251 21419 10257
rect 21361 10248 21373 10251
rect 19024 10220 21373 10248
rect 19024 10208 19030 10220
rect 21361 10217 21373 10220
rect 21407 10217 21419 10251
rect 21361 10211 21419 10217
rect 17405 10183 17463 10189
rect 17405 10149 17417 10183
rect 17451 10149 17463 10183
rect 17405 10143 17463 10149
rect 22925 10183 22983 10189
rect 22925 10149 22937 10183
rect 22971 10180 22983 10183
rect 23198 10180 23204 10192
rect 22971 10152 23204 10180
rect 22971 10149 22983 10152
rect 22925 10143 22983 10149
rect 23198 10140 23204 10152
rect 23256 10140 23262 10192
rect 23474 10140 23480 10192
rect 23532 10180 23538 10192
rect 23532 10152 23577 10180
rect 23532 10140 23538 10152
rect 24210 10140 24216 10192
rect 24268 10180 24274 10192
rect 24489 10183 24547 10189
rect 24489 10180 24501 10183
rect 24268 10152 24501 10180
rect 24268 10140 24274 10152
rect 24489 10149 24501 10152
rect 24535 10149 24547 10183
rect 24489 10143 24547 10149
rect 19058 10112 19064 10124
rect 19019 10084 19064 10112
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 19242 10112 19248 10124
rect 19203 10084 19248 10112
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 20438 10072 20444 10124
rect 20496 10112 20502 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20496 10084 20913 10112
rect 20496 10072 20502 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 21177 10115 21235 10121
rect 21177 10081 21189 10115
rect 21223 10112 21235 10115
rect 21358 10112 21364 10124
rect 21223 10084 21364 10112
rect 21223 10081 21235 10084
rect 21177 10075 21235 10081
rect 12860 10016 16160 10044
rect 17313 10047 17371 10053
rect 12860 10004 12866 10016
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10044 18015 10047
rect 18322 10044 18328 10056
rect 18003 10016 18328 10044
rect 18003 10013 18015 10016
rect 17957 10007 18015 10013
rect 6135 9979 6193 9985
rect 6135 9945 6147 9979
rect 6181 9976 6193 9979
rect 10410 9976 10416 9988
rect 6181 9948 10416 9976
rect 6181 9945 6193 9948
rect 6135 9939 6193 9945
rect 10410 9936 10416 9948
rect 10468 9936 10474 9988
rect 14090 9976 14096 9988
rect 14051 9948 14096 9976
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 12894 9908 12900 9920
rect 10192 9880 12900 9908
rect 10192 9868 10198 9880
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 14274 9868 14280 9920
rect 14332 9908 14338 9920
rect 14737 9911 14795 9917
rect 14737 9908 14749 9911
rect 14332 9880 14749 9908
rect 14332 9868 14338 9880
rect 14737 9877 14749 9880
rect 14783 9908 14795 9911
rect 14826 9908 14832 9920
rect 14783 9880 14832 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 17034 9908 17040 9920
rect 16995 9880 17040 9908
rect 17034 9868 17040 9880
rect 17092 9908 17098 9920
rect 17328 9908 17356 10007
rect 18322 10004 18328 10016
rect 18380 10044 18386 10056
rect 18782 10044 18788 10056
rect 18380 10016 18788 10044
rect 18380 10004 18386 10016
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 20916 10044 20944 10075
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 20916 10016 21925 10044
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 22830 10044 22836 10056
rect 22791 10016 22836 10044
rect 21913 10007 21971 10013
rect 22830 10004 22836 10016
rect 22888 10044 22894 10056
rect 24397 10047 24455 10053
rect 22888 10016 23474 10044
rect 22888 10004 22894 10016
rect 18690 9936 18696 9988
rect 18748 9976 18754 9988
rect 20622 9976 20628 9988
rect 18748 9948 20628 9976
rect 18748 9936 18754 9948
rect 20622 9936 20628 9948
rect 20680 9936 20686 9988
rect 20990 9976 20996 9988
rect 20951 9948 20996 9976
rect 20990 9936 20996 9948
rect 21048 9936 21054 9988
rect 23446 9976 23474 10016
rect 24397 10013 24409 10047
rect 24443 10044 24455 10047
rect 24762 10044 24768 10056
rect 24443 10016 24768 10044
rect 24443 10013 24455 10016
rect 24397 10007 24455 10013
rect 24762 10004 24768 10016
rect 24820 10044 24826 10056
rect 25222 10044 25228 10056
rect 24820 10016 25228 10044
rect 24820 10004 24826 10016
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 23566 9976 23572 9988
rect 23446 9948 23572 9976
rect 23566 9936 23572 9948
rect 23624 9936 23630 9988
rect 24118 9936 24124 9988
rect 24176 9976 24182 9988
rect 24949 9979 25007 9985
rect 24949 9976 24961 9979
rect 24176 9948 24961 9976
rect 24176 9936 24182 9948
rect 24949 9945 24961 9948
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 17092 9880 17356 9908
rect 19889 9911 19947 9917
rect 17092 9868 17098 9880
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20070 9908 20076 9920
rect 19935 9880 20076 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 20162 9868 20168 9920
rect 20220 9908 20226 9920
rect 20257 9911 20315 9917
rect 20257 9908 20269 9911
rect 20220 9880 20269 9908
rect 20220 9868 20226 9880
rect 20257 9877 20269 9880
rect 20303 9908 20315 9911
rect 21358 9908 21364 9920
rect 20303 9880 21364 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 22278 9908 22284 9920
rect 22239 9880 22284 9908
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 24210 9908 24216 9920
rect 23348 9880 24216 9908
rect 23348 9868 23354 9880
rect 24210 9868 24216 9880
rect 24268 9868 24274 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 5997 9707 6055 9713
rect 5997 9673 6009 9707
rect 6043 9704 6055 9707
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 6043 9676 6285 9704
rect 6043 9673 6055 9676
rect 5997 9667 6055 9673
rect 6273 9673 6285 9676
rect 6319 9704 6331 9707
rect 7098 9704 7104 9716
rect 6319 9676 7104 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8481 9707 8539 9713
rect 8481 9673 8493 9707
rect 8527 9704 8539 9707
rect 9214 9704 9220 9716
rect 8527 9676 9220 9704
rect 8527 9673 8539 9676
rect 8481 9667 8539 9673
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 9858 9704 9864 9716
rect 9819 9676 9864 9704
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 10008 9676 10149 9704
rect 10008 9664 10014 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 10284 9676 11805 9704
rect 10284 9664 10290 9676
rect 11793 9673 11805 9676
rect 11839 9704 11851 9707
rect 12250 9704 12256 9716
rect 11839 9676 12256 9704
rect 11839 9673 11851 9676
rect 11793 9667 11851 9673
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 13357 9707 13415 9713
rect 13357 9673 13369 9707
rect 13403 9704 13415 9707
rect 13630 9704 13636 9716
rect 13403 9676 13636 9704
rect 13403 9673 13415 9676
rect 13357 9667 13415 9673
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 14783 9707 14841 9713
rect 14783 9704 14795 9707
rect 14700 9676 14795 9704
rect 14700 9664 14706 9676
rect 14783 9673 14795 9676
rect 14829 9673 14841 9707
rect 14783 9667 14841 9673
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15930 9704 15936 9716
rect 15712 9676 15936 9704
rect 15712 9664 15718 9676
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 17218 9704 17224 9716
rect 17179 9676 17224 9704
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 19058 9704 19064 9716
rect 19019 9676 19064 9704
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 23477 9707 23535 9713
rect 23477 9673 23489 9707
rect 23523 9704 23535 9707
rect 23566 9704 23572 9716
rect 23523 9676 23572 9704
rect 23523 9673 23535 9676
rect 23477 9667 23535 9673
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 24210 9704 24216 9716
rect 24171 9676 24216 9704
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 6638 9636 6644 9648
rect 6551 9608 6644 9636
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 11974 9636 11980 9648
rect 6696 9608 11980 9636
rect 6696 9596 6702 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 13538 9596 13544 9648
rect 13596 9636 13602 9648
rect 14001 9639 14059 9645
rect 14001 9636 14013 9639
rect 13596 9608 14013 9636
rect 13596 9596 13602 9608
rect 14001 9605 14013 9608
rect 14047 9605 14059 9639
rect 14001 9599 14059 9605
rect 14921 9639 14979 9645
rect 14921 9605 14933 9639
rect 14967 9636 14979 9639
rect 15197 9639 15255 9645
rect 15197 9636 15209 9639
rect 14967 9608 15209 9636
rect 14967 9605 14979 9608
rect 14921 9599 14979 9605
rect 15197 9605 15209 9608
rect 15243 9636 15255 9639
rect 22186 9636 22192 9648
rect 15243 9608 22192 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 22186 9596 22192 9608
rect 22244 9596 22250 9648
rect 25409 9639 25467 9645
rect 25409 9636 25421 9639
rect 24504 9608 25421 9636
rect 4847 9571 4905 9577
rect 4847 9537 4859 9571
rect 4893 9568 4905 9571
rect 9306 9568 9312 9580
rect 4893 9540 9312 9568
rect 4893 9537 4905 9540
rect 4847 9531 4905 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 10410 9568 10416 9580
rect 10371 9540 10416 9568
rect 10410 9528 10416 9540
rect 10468 9568 10474 9580
rect 11054 9568 11060 9580
rect 10468 9540 11060 9568
rect 10468 9528 10474 9540
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 12434 9568 12440 9580
rect 12395 9540 12440 9568
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 14148 9540 16037 9568
rect 14148 9528 14154 9540
rect 16025 9537 16037 9540
rect 16071 9568 16083 9571
rect 17034 9568 17040 9580
rect 16071 9540 17040 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18230 9568 18236 9580
rect 18187 9540 18236 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 18782 9568 18788 9580
rect 18743 9540 18788 9568
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9568 21879 9571
rect 22278 9568 22284 9580
rect 21867 9540 22284 9568
rect 21867 9537 21879 9540
rect 21821 9531 21879 9537
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 24118 9528 24124 9580
rect 24176 9568 24182 9580
rect 24504 9577 24532 9608
rect 25409 9605 25421 9608
rect 25455 9605 25467 9639
rect 25409 9599 25467 9605
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 24176 9540 24501 9568
rect 24176 9528 24182 9540
rect 24489 9537 24501 9540
rect 24535 9537 24547 9571
rect 24946 9568 24952 9580
rect 24907 9540 24952 9568
rect 24489 9531 24547 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 4760 9503 4818 9509
rect 4760 9469 4772 9503
rect 4806 9500 4818 9503
rect 5788 9503 5846 9509
rect 4806 9472 5212 9500
rect 4806 9469 4818 9472
rect 4760 9463 4818 9469
rect 5184 9376 5212 9472
rect 5788 9469 5800 9503
rect 5834 9500 5846 9503
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5834 9472 6009 9500
rect 5834 9469 5846 9472
rect 5788 9463 5846 9469
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 7612 9503 7670 9509
rect 7612 9469 7624 9503
rect 7658 9500 7670 9503
rect 8110 9500 8116 9512
rect 7658 9472 8116 9500
rect 7658 9469 7670 9472
rect 7612 9463 7670 9469
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9214 9500 9220 9512
rect 8956 9472 9220 9500
rect 7699 9435 7757 9441
rect 7699 9401 7711 9435
rect 7745 9432 7757 9435
rect 8754 9432 8760 9444
rect 7745 9404 8760 9432
rect 7745 9401 7757 9404
rect 7699 9395 7757 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 8956 9441 8984 9472
rect 9214 9460 9220 9472
rect 9272 9500 9278 9512
rect 10226 9500 10232 9512
rect 9272 9472 10232 9500
rect 9272 9460 9278 9472
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 14712 9503 14770 9509
rect 14712 9469 14724 9503
rect 14758 9500 14770 9503
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 14758 9472 14933 9500
rect 14758 9469 14770 9472
rect 14712 9463 14770 9469
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19536 9500 19564 9528
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 19475 9472 20269 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 8935 9435 8993 9441
rect 8935 9401 8947 9435
rect 8981 9401 8993 9435
rect 10505 9435 10563 9441
rect 10505 9432 10517 9435
rect 8935 9395 8993 9401
rect 9508 9404 10517 9432
rect 5166 9364 5172 9376
rect 5127 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5859 9367 5917 9373
rect 5859 9333 5871 9367
rect 5905 9364 5917 9367
rect 6086 9364 6092 9376
rect 5905 9336 6092 9364
rect 5905 9333 5917 9336
rect 5859 9327 5917 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 7469 9367 7527 9373
rect 7469 9333 7481 9367
rect 7515 9364 7527 9367
rect 8018 9364 8024 9376
rect 7515 9336 8024 9364
rect 7515 9333 7527 9336
rect 7469 9327 7527 9333
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 9508 9373 9536 9404
rect 10505 9401 10517 9404
rect 10551 9401 10563 9435
rect 10505 9395 10563 9401
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 8720 9336 9505 9364
rect 8720 9324 8726 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 10520 9364 10548 9395
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 10836 9404 11069 9432
rect 10836 9392 10842 9404
rect 11057 9401 11069 9404
rect 11103 9401 11115 9435
rect 11057 9395 11115 9401
rect 12250 9392 12256 9444
rect 12308 9432 12314 9444
rect 12758 9435 12816 9441
rect 12758 9432 12770 9435
rect 12308 9404 12770 9432
rect 12308 9392 12314 9404
rect 12758 9401 12770 9404
rect 12804 9401 12816 9435
rect 12758 9395 12816 9401
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 15749 9435 15807 9441
rect 15749 9432 15761 9435
rect 14240 9404 15761 9432
rect 14240 9392 14246 9404
rect 15749 9401 15761 9404
rect 15795 9401 15807 9435
rect 15749 9395 15807 9401
rect 15841 9435 15899 9441
rect 15841 9401 15853 9435
rect 15887 9432 15899 9435
rect 16206 9432 16212 9444
rect 15887 9404 16212 9432
rect 15887 9401 15899 9404
rect 15841 9395 15899 9401
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 10520 9336 11345 9364
rect 9493 9327 9551 9333
rect 11333 9333 11345 9336
rect 11379 9364 11391 9367
rect 11606 9364 11612 9376
rect 11379 9336 11612 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 15565 9367 15623 9373
rect 15565 9333 15577 9367
rect 15611 9364 15623 9367
rect 15654 9364 15660 9376
rect 15611 9336 15660 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 15764 9364 15792 9395
rect 16206 9392 16212 9404
rect 16264 9392 16270 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 15764 9336 16681 9364
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 16669 9327 16727 9333
rect 17865 9367 17923 9373
rect 17865 9333 17877 9367
rect 17911 9364 17923 9367
rect 17954 9364 17960 9376
rect 17911 9336 17960 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 17954 9324 17960 9336
rect 18012 9364 18018 9376
rect 18248 9364 18276 9395
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19613 9435 19671 9441
rect 19613 9432 19625 9435
rect 19576 9404 19625 9432
rect 19576 9392 19582 9404
rect 19613 9401 19625 9404
rect 19659 9401 19671 9435
rect 20272 9432 20300 9463
rect 20990 9432 20996 9444
rect 20272 9404 20996 9432
rect 19613 9395 19671 9401
rect 20990 9392 20996 9404
rect 21048 9432 21054 9444
rect 21450 9432 21456 9444
rect 21048 9404 21456 9432
rect 21048 9392 21054 9404
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 21729 9435 21787 9441
rect 21729 9401 21741 9435
rect 21775 9432 21787 9435
rect 22183 9435 22241 9441
rect 22183 9432 22195 9435
rect 21775 9404 22195 9432
rect 21775 9401 21787 9404
rect 21729 9395 21787 9401
rect 22183 9401 22195 9404
rect 22229 9432 22241 9435
rect 22922 9432 22928 9444
rect 22229 9404 22928 9432
rect 22229 9401 22241 9404
rect 22183 9395 22241 9401
rect 22922 9392 22928 9404
rect 22980 9432 22986 9444
rect 23566 9432 23572 9444
rect 22980 9404 23572 9432
rect 22980 9392 22986 9404
rect 23566 9392 23572 9404
rect 23624 9392 23630 9444
rect 23937 9435 23995 9441
rect 23937 9401 23949 9435
rect 23983 9432 23995 9435
rect 24581 9435 24639 9441
rect 23983 9404 24440 9432
rect 23983 9401 23995 9404
rect 23937 9395 23995 9401
rect 21358 9364 21364 9376
rect 18012 9336 18276 9364
rect 21319 9336 21364 9364
rect 18012 9324 18018 9336
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 22741 9367 22799 9373
rect 22741 9333 22753 9367
rect 22787 9364 22799 9367
rect 23109 9367 23167 9373
rect 23109 9364 23121 9367
rect 22787 9336 23121 9364
rect 22787 9333 22799 9336
rect 22741 9327 22799 9333
rect 23109 9333 23121 9336
rect 23155 9364 23167 9367
rect 23198 9364 23204 9376
rect 23155 9336 23204 9364
rect 23155 9333 23167 9336
rect 23109 9327 23167 9333
rect 23198 9324 23204 9336
rect 23256 9324 23262 9376
rect 24412 9364 24440 9404
rect 24581 9401 24593 9435
rect 24627 9432 24639 9435
rect 24670 9432 24676 9444
rect 24627 9404 24676 9432
rect 24627 9401 24639 9404
rect 24581 9395 24639 9401
rect 24596 9364 24624 9395
rect 24670 9392 24676 9404
rect 24728 9392 24734 9444
rect 24412 9336 24624 9364
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6144 9132 9812 9160
rect 6144 9120 6150 9132
rect 9784 9104 9812 9132
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10192 9132 10701 9160
rect 10192 9120 10198 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 10689 9123 10747 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11330 9160 11336 9172
rect 11291 9132 11336 9160
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12434 9160 12440 9172
rect 12395 9132 12440 9160
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 15470 9160 15476 9172
rect 15151 9132 15476 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 16206 9160 16212 9172
rect 16167 9132 16212 9160
rect 16206 9120 16212 9132
rect 16264 9160 16270 9172
rect 16390 9160 16396 9172
rect 16264 9132 16396 9160
rect 16264 9120 16270 9132
rect 16390 9120 16396 9132
rect 16448 9160 16454 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16448 9132 16497 9160
rect 16448 9120 16454 9132
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 17954 9160 17960 9172
rect 17915 9132 17960 9160
rect 16485 9123 16543 9129
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 20349 9163 20407 9169
rect 20349 9129 20361 9163
rect 20395 9160 20407 9163
rect 20438 9160 20444 9172
rect 20395 9132 20444 9160
rect 20395 9129 20407 9132
rect 20349 9123 20407 9129
rect 7193 9095 7251 9101
rect 7193 9061 7205 9095
rect 7239 9092 7251 9095
rect 8570 9092 8576 9104
rect 7239 9064 8576 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 8570 9052 8576 9064
rect 8628 9092 8634 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8628 9064 9045 9092
rect 8628 9052 8634 9064
rect 9033 9061 9045 9064
rect 9079 9061 9091 9095
rect 9766 9092 9772 9104
rect 9679 9064 9772 9092
rect 9033 9055 9091 9061
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 9916 9064 9961 9092
rect 9916 9052 9922 9064
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 13541 9095 13599 9101
rect 13541 9092 13553 9095
rect 12676 9064 13553 9092
rect 12676 9052 12682 9064
rect 13541 9061 13553 9064
rect 13587 9061 13599 9095
rect 14090 9092 14096 9104
rect 14051 9064 14096 9092
rect 13541 9055 13599 9061
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 17358 9095 17416 9101
rect 17358 9092 17370 9095
rect 17276 9064 17370 9092
rect 17276 9052 17282 9064
rect 17358 9061 17370 9064
rect 17404 9061 17416 9095
rect 17358 9055 17416 9061
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 18785 9095 18843 9101
rect 18785 9092 18797 9095
rect 17828 9064 18797 9092
rect 17828 9052 17834 9064
rect 18785 9061 18797 9064
rect 18831 9092 18843 9095
rect 18966 9092 18972 9104
rect 18831 9064 18972 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 19978 9092 19984 9104
rect 19168 9064 19984 9092
rect 5442 9024 5448 9036
rect 5403 8996 5448 9024
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 6546 9024 6552 9036
rect 6507 8996 6552 9024
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6656 8996 7021 9024
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 6656 8888 6684 8996
rect 7009 8993 7021 8996
rect 7055 9024 7067 9027
rect 7374 9024 7380 9036
rect 7055 8996 7380 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8478 9024 8484 9036
rect 8439 8996 8484 9024
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 11422 9024 11428 9036
rect 11383 8996 11428 9024
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 11882 9024 11888 9036
rect 11839 8996 11888 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 15286 9024 15292 9036
rect 15199 8996 15292 9024
rect 15286 8984 15292 8996
rect 15344 9024 15350 9036
rect 16298 9024 16304 9036
rect 15344 8996 16304 9024
rect 15344 8984 15350 8996
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 19168 9033 19196 9064
rect 19978 9052 19984 9064
rect 20036 9092 20042 9104
rect 20364 9092 20392 9123
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 20622 9160 20628 9172
rect 20583 9132 20628 9160
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 24673 9163 24731 9169
rect 24673 9129 24685 9163
rect 24719 9160 24731 9163
rect 24762 9160 24768 9172
rect 24719 9132 24768 9160
rect 24719 9129 24731 9132
rect 24673 9123 24731 9129
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 20036 9064 20392 9092
rect 20036 9052 20042 9064
rect 23566 9052 23572 9104
rect 23624 9092 23630 9104
rect 23706 9095 23764 9101
rect 23706 9092 23718 9095
rect 23624 9064 23718 9092
rect 23624 9052 23630 9064
rect 23706 9061 23718 9064
rect 23752 9061 23764 9095
rect 23706 9055 23764 9061
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 9024 19487 9027
rect 19702 9024 19708 9036
rect 19475 8996 19708 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 21085 9027 21143 9033
rect 21085 9024 21097 9027
rect 20864 8996 21097 9024
rect 20864 8984 20870 8996
rect 21085 8993 21097 8996
rect 21131 8993 21143 9027
rect 21085 8987 21143 8993
rect 21266 8984 21272 9036
rect 21324 9024 21330 9036
rect 21545 9027 21603 9033
rect 21545 9024 21557 9027
rect 21324 8996 21557 9024
rect 21324 8984 21330 8996
rect 21545 8993 21557 8996
rect 21591 8993 21603 9027
rect 21910 9024 21916 9036
rect 21871 8996 21916 9024
rect 21545 8987 21603 8993
rect 21910 8984 21916 8996
rect 21968 8984 21974 9036
rect 22281 9027 22339 9033
rect 22281 8993 22293 9027
rect 22327 8993 22339 9027
rect 22281 8987 22339 8993
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 6788 8928 7481 8956
rect 6788 8916 6794 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 7469 8919 7527 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 13170 8956 13176 8968
rect 8812 8928 13176 8956
rect 8812 8916 8818 8928
rect 13170 8916 13176 8928
rect 13228 8956 13234 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13228 8928 13461 8956
rect 13228 8916 13234 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8956 17095 8959
rect 17678 8956 17684 8968
rect 17083 8928 17684 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 19613 8959 19671 8965
rect 19613 8956 19625 8959
rect 17828 8928 19625 8956
rect 17828 8916 17834 8928
rect 19613 8925 19625 8928
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 22002 8956 22008 8968
rect 21692 8928 22008 8956
rect 21692 8916 21698 8928
rect 22002 8916 22008 8928
rect 22060 8956 22066 8968
rect 22296 8956 22324 8987
rect 22060 8928 22324 8956
rect 22557 8959 22615 8965
rect 22060 8916 22066 8928
rect 22557 8925 22569 8959
rect 22603 8956 22615 8959
rect 23385 8959 23443 8965
rect 23385 8956 23397 8959
rect 22603 8928 23397 8956
rect 22603 8925 22615 8928
rect 22557 8919 22615 8925
rect 23385 8925 23397 8928
rect 23431 8956 23443 8959
rect 24026 8956 24032 8968
rect 23431 8928 24032 8956
rect 23431 8925 23443 8928
rect 23385 8919 23443 8925
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 24210 8916 24216 8968
rect 24268 8956 24274 8968
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 24268 8928 25145 8956
rect 24268 8916 24274 8928
rect 25133 8925 25145 8928
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 5675 8860 6684 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 10318 8888 10324 8900
rect 8996 8860 10324 8888
rect 8996 8848 9002 8860
rect 10318 8848 10324 8860
rect 10376 8888 10382 8900
rect 10778 8888 10784 8900
rect 10376 8860 10784 8888
rect 10376 8848 10382 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 14182 8888 14188 8900
rect 11204 8860 14188 8888
rect 11204 8848 11210 8860
rect 14182 8848 14188 8860
rect 14240 8848 14246 8900
rect 19245 8891 19303 8897
rect 19245 8857 19257 8891
rect 19291 8888 19303 8891
rect 19518 8888 19524 8900
rect 19291 8860 19524 8888
rect 19291 8857 19303 8860
rect 19245 8851 19303 8857
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 11054 8820 11060 8832
rect 8168 8792 11060 8820
rect 8168 8780 8174 8792
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16853 8823 16911 8829
rect 16853 8820 16865 8823
rect 16632 8792 16865 8820
rect 16632 8780 16638 8792
rect 16853 8789 16865 8792
rect 16899 8789 16911 8823
rect 18230 8820 18236 8832
rect 18191 8792 18236 8820
rect 16853 8783 16911 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 24305 8823 24363 8829
rect 24305 8789 24317 8823
rect 24351 8820 24363 8823
rect 24854 8820 24860 8832
rect 24351 8792 24860 8820
rect 24351 8789 24363 8792
rect 24305 8783 24363 8789
rect 24854 8780 24860 8792
rect 24912 8820 24918 8832
rect 25222 8820 25228 8832
rect 24912 8792 25228 8820
rect 24912 8780 24918 8792
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9824 8588 10057 8616
rect 9824 8576 9830 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12676 8588 12817 8616
rect 12676 8576 12682 8588
rect 12805 8585 12817 8588
rect 12851 8616 12863 8619
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12851 8588 13185 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 13173 8585 13185 8588
rect 13219 8616 13231 8619
rect 13538 8616 13544 8628
rect 13219 8588 13544 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 15105 8619 15163 8625
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15286 8616 15292 8628
rect 15151 8588 15292 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 17218 8616 17224 8628
rect 15979 8588 17224 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 19702 8616 19708 8628
rect 19615 8588 19708 8616
rect 19702 8576 19708 8588
rect 19760 8616 19766 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 19760 8588 20361 8616
rect 19760 8576 19766 8588
rect 20349 8585 20361 8588
rect 20395 8616 20407 8619
rect 20898 8616 20904 8628
rect 20395 8588 20904 8616
rect 20395 8585 20407 8588
rect 20349 8579 20407 8585
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 23109 8619 23167 8625
rect 23109 8585 23121 8619
rect 23155 8616 23167 8619
rect 23290 8616 23296 8628
rect 23155 8588 23296 8616
rect 23155 8585 23167 8588
rect 23109 8579 23167 8585
rect 23290 8576 23296 8588
rect 23348 8616 23354 8628
rect 23842 8616 23848 8628
rect 23348 8588 23848 8616
rect 23348 8576 23354 8588
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 24026 8576 24032 8628
rect 24084 8616 24090 8628
rect 24673 8619 24731 8625
rect 24673 8616 24685 8619
rect 24084 8588 24685 8616
rect 24084 8576 24090 8588
rect 24673 8585 24685 8588
rect 24719 8585 24731 8619
rect 24673 8579 24731 8585
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 9640 8520 13492 8548
rect 9640 8508 9646 8520
rect 13464 8492 13492 8520
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 18187 8551 18245 8557
rect 18187 8548 18199 8551
rect 13780 8520 18199 8548
rect 13780 8508 13786 8520
rect 18187 8517 18199 8520
rect 18233 8517 18245 8551
rect 18187 8511 18245 8517
rect 21358 8508 21364 8560
rect 21416 8548 21422 8560
rect 25409 8551 25467 8557
rect 25409 8548 25421 8551
rect 21416 8520 25421 8548
rect 21416 8508 21422 8520
rect 25409 8517 25421 8520
rect 25455 8517 25467 8551
rect 25409 8511 25467 8517
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8570 8480 8576 8492
rect 8527 8452 8576 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10376 8452 10885 8480
rect 10376 8440 10382 8452
rect 10873 8449 10885 8452
rect 10919 8480 10931 8483
rect 12161 8483 12219 8489
rect 12161 8480 12173 8483
rect 10919 8452 12173 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 12161 8449 12173 8452
rect 12207 8449 12219 8483
rect 13446 8480 13452 8492
rect 13359 8452 13452 8480
rect 12161 8443 12219 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 15335 8483 15393 8489
rect 15335 8449 15347 8483
rect 15381 8480 15393 8483
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 15381 8452 16313 8480
rect 15381 8449 15393 8452
rect 15335 8443 15393 8449
rect 16301 8449 16313 8452
rect 16347 8480 16359 8483
rect 16574 8480 16580 8492
rect 16347 8452 16580 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 22278 8480 22284 8492
rect 20680 8452 22048 8480
rect 22239 8452 22284 8480
rect 20680 8440 20686 8452
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8412 5227 8415
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5215 8384 5733 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 5721 8381 5733 8384
rect 5767 8412 5779 8415
rect 5994 8412 6000 8424
rect 5767 8384 6000 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6788 8384 6929 8412
rect 6788 8372 6794 8384
rect 6917 8381 6929 8384
rect 6963 8412 6975 8415
rect 7282 8412 7288 8424
rect 6963 8384 7288 8412
rect 6963 8381 6975 8384
rect 6917 8375 6975 8381
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7466 8412 7472 8424
rect 7427 8384 7472 8412
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 15232 8415 15290 8421
rect 15232 8412 15244 8415
rect 15068 8384 15244 8412
rect 15068 8372 15074 8384
rect 15232 8381 15244 8384
rect 15278 8381 15290 8415
rect 15232 8375 15290 8381
rect 15654 8372 15660 8424
rect 15712 8412 15718 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15712 8384 15945 8412
rect 15712 8372 15718 8384
rect 15933 8381 15945 8384
rect 15979 8412 15991 8415
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15979 8384 16037 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 18116 8415 18174 8421
rect 18116 8381 18128 8415
rect 18162 8412 18174 8415
rect 19153 8415 19211 8421
rect 18162 8384 18460 8412
rect 18162 8381 18174 8384
rect 18116 8375 18174 8381
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5537 8347 5595 8353
rect 5537 8344 5549 8347
rect 5500 8316 5549 8344
rect 5500 8304 5506 8316
rect 5537 8313 5549 8316
rect 5583 8344 5595 8347
rect 6086 8344 6092 8356
rect 5583 8316 6092 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 7653 8347 7711 8353
rect 7653 8313 7665 8347
rect 7699 8344 7711 8347
rect 8202 8344 8208 8356
rect 7699 8316 8208 8344
rect 7699 8313 7711 8316
rect 7653 8307 7711 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8389 8347 8447 8353
rect 8389 8313 8401 8347
rect 8435 8344 8447 8347
rect 8843 8347 8901 8353
rect 8843 8344 8855 8347
rect 8435 8316 8855 8344
rect 8435 8313 8447 8316
rect 8389 8307 8447 8313
rect 8843 8313 8855 8316
rect 8889 8344 8901 8347
rect 9214 8344 9220 8356
rect 8889 8316 9220 8344
rect 8889 8313 8901 8316
rect 8843 8307 8901 8313
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11020 8316 11065 8344
rect 11020 8304 11026 8316
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11204 8316 11529 8344
rect 11204 8304 11210 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 14090 8344 14096 8356
rect 13596 8316 13641 8344
rect 14051 8316 14096 8344
rect 13596 8304 13602 8316
rect 14090 8304 14096 8316
rect 14148 8344 14154 8356
rect 16390 8344 16396 8356
rect 14148 8316 16252 8344
rect 16351 8316 16396 8344
rect 14148 8304 14154 8316
rect 5905 8279 5963 8285
rect 5905 8245 5917 8279
rect 5951 8276 5963 8279
rect 6362 8276 6368 8288
rect 5951 8248 6368 8276
rect 5951 8245 5963 8248
rect 5905 8239 5963 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 6822 8276 6828 8288
rect 6604 8248 6828 8276
rect 6604 8236 6610 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 8018 8276 8024 8288
rect 7979 8248 8024 8276
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 9398 8276 9404 8288
rect 9359 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8276 9462 8288
rect 9677 8279 9735 8285
rect 9677 8276 9689 8279
rect 9456 8248 9689 8276
rect 9456 8236 9462 8248
rect 9677 8245 9689 8248
rect 9723 8276 9735 8279
rect 9858 8276 9864 8288
rect 9723 8248 9864 8276
rect 9723 8245 9735 8248
rect 9677 8239 9735 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 10980 8276 11008 8304
rect 11882 8276 11888 8288
rect 10735 8248 11008 8276
rect 11843 8248 11888 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14369 8279 14427 8285
rect 14369 8276 14381 8279
rect 13504 8248 14381 8276
rect 13504 8236 13510 8248
rect 14369 8245 14381 8248
rect 14415 8245 14427 8279
rect 14369 8239 14427 8245
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 15657 8279 15715 8285
rect 15657 8276 15669 8279
rect 15068 8248 15669 8276
rect 15068 8236 15074 8248
rect 15657 8245 15669 8248
rect 15703 8276 15715 8279
rect 16114 8276 16120 8288
rect 15703 8248 16120 8276
rect 15703 8245 15715 8248
rect 15657 8239 15715 8245
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 16224 8276 16252 8316
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 16945 8347 17003 8353
rect 16945 8313 16957 8347
rect 16991 8344 17003 8347
rect 18230 8344 18236 8356
rect 16991 8316 18236 8344
rect 16991 8313 17003 8316
rect 16945 8307 17003 8313
rect 16960 8276 16988 8307
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 18432 8288 18460 8384
rect 19153 8381 19165 8415
rect 19199 8412 19211 8415
rect 19886 8412 19892 8424
rect 19199 8384 19892 8412
rect 19199 8381 19211 8384
rect 19153 8375 19211 8381
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 20806 8412 20812 8424
rect 20767 8384 20812 8412
rect 20806 8372 20812 8384
rect 20864 8372 20870 8424
rect 21266 8412 21272 8424
rect 21227 8384 21272 8412
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21637 8415 21695 8421
rect 21637 8381 21649 8415
rect 21683 8412 21695 8415
rect 21910 8412 21916 8424
rect 21683 8384 21916 8412
rect 21683 8381 21695 8384
rect 21637 8375 21695 8381
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 21652 8344 21680 8375
rect 21910 8372 21916 8384
rect 21968 8372 21974 8424
rect 22020 8421 22048 8452
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 24029 8483 24087 8489
rect 24029 8480 24041 8483
rect 23440 8452 24041 8480
rect 23440 8440 23446 8452
rect 24029 8449 24041 8452
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8381 22063 8415
rect 22005 8375 22063 8381
rect 22554 8372 22560 8424
rect 22612 8372 22618 8424
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 25096 8384 25237 8412
rect 25096 8372 25102 8384
rect 25225 8381 25237 8384
rect 25271 8412 25283 8415
rect 25271 8384 25728 8412
rect 25271 8381 25283 8384
rect 25225 8375 25283 8381
rect 20036 8316 21680 8344
rect 22572 8344 22600 8372
rect 23750 8344 23756 8356
rect 22572 8316 23756 8344
rect 20036 8304 20042 8316
rect 23750 8304 23756 8316
rect 23808 8304 23814 8356
rect 23842 8304 23848 8356
rect 23900 8344 23906 8356
rect 23900 8316 23945 8344
rect 23900 8304 23906 8316
rect 25700 8288 25728 8384
rect 17678 8276 17684 8288
rect 16224 8248 16988 8276
rect 17639 8248 17684 8276
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 18509 8279 18567 8285
rect 18509 8276 18521 8279
rect 18472 8248 18521 8276
rect 18472 8236 18478 8248
rect 18509 8245 18521 8248
rect 18555 8245 18567 8279
rect 20622 8276 20628 8288
rect 20583 8248 20628 8276
rect 18509 8239 18567 8245
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 21726 8236 21732 8288
rect 21784 8276 21790 8288
rect 22462 8276 22468 8288
rect 21784 8248 22468 8276
rect 21784 8236 21790 8248
rect 22462 8236 22468 8248
rect 22520 8276 22526 8288
rect 22557 8279 22615 8285
rect 22557 8276 22569 8279
rect 22520 8248 22569 8276
rect 22520 8236 22526 8248
rect 22557 8245 22569 8248
rect 22603 8245 22615 8279
rect 22557 8239 22615 8245
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23566 8276 23572 8288
rect 23523 8248 23572 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23566 8236 23572 8248
rect 23624 8236 23630 8288
rect 25682 8276 25688 8288
rect 25643 8248 25688 8276
rect 25682 8236 25688 8248
rect 25740 8236 25746 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7466 8072 7472 8084
rect 7147 8044 7472 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7466 8032 7472 8044
rect 7524 8072 7530 8084
rect 7524 8044 8524 8072
rect 7524 8032 7530 8044
rect 8496 8016 8524 8044
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8628 8044 8953 8072
rect 8628 8032 8634 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 9766 8072 9772 8084
rect 9727 8044 9772 8072
rect 8941 8035 8999 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 10778 8072 10784 8084
rect 10691 8044 10784 8072
rect 10778 8032 10784 8044
rect 10836 8072 10842 8084
rect 11330 8072 11336 8084
rect 10836 8044 11336 8072
rect 10836 8032 10842 8044
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 13170 8072 13176 8084
rect 11480 8044 12801 8072
rect 13131 8044 13176 8072
rect 11480 8032 11486 8044
rect 7742 8004 7748 8016
rect 7703 7976 7748 8004
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 7892 7976 8340 8004
rect 7892 7964 7898 7976
rect 5534 7936 5540 7948
rect 5495 7908 5540 7936
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 8312 7936 8340 7976
rect 8478 7964 8484 8016
rect 8536 8004 8542 8016
rect 8665 8007 8723 8013
rect 8665 8004 8677 8007
rect 8536 7976 8677 8004
rect 8536 7964 8542 7976
rect 8665 7973 8677 7976
rect 8711 8004 8723 8007
rect 11606 8004 11612 8016
rect 8711 7976 10180 8004
rect 11567 7976 11612 8004
rect 8711 7973 8723 7976
rect 8665 7967 8723 7973
rect 10152 7948 10180 7976
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 12773 8004 12801 8044
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 14274 8072 14280 8084
rect 13274 8044 14280 8072
rect 13274 8004 13302 8044
rect 14274 8032 14280 8044
rect 14332 8072 14338 8084
rect 14332 8044 15700 8072
rect 14332 8032 14338 8044
rect 12773 7976 13302 8004
rect 13541 8007 13599 8013
rect 13541 7973 13553 8007
rect 13587 8004 13599 8007
rect 13630 8004 13636 8016
rect 13587 7976 13636 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 14090 8004 14096 8016
rect 14051 7976 14096 8004
rect 14090 7964 14096 7976
rect 14148 7964 14154 8016
rect 9490 7936 9496 7948
rect 6595 7908 7052 7936
rect 8312 7908 9496 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 7024 7880 7052 7908
rect 9490 7896 9496 7908
rect 9548 7936 9554 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9548 7908 9689 7936
rect 9548 7896 9554 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 15672 7945 15700 8044
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 16761 8075 16819 8081
rect 16761 8072 16773 8075
rect 16448 8044 16773 8072
rect 16448 8032 16454 8044
rect 16761 8041 16773 8044
rect 16807 8072 16819 8075
rect 16807 8044 17172 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17144 8016 17172 8044
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 17736 8044 18613 8072
rect 17736 8032 17742 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 19518 8072 19524 8084
rect 19479 8044 19524 8072
rect 18601 8035 18659 8041
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 19978 8072 19984 8084
rect 19939 8044 19984 8072
rect 19978 8032 19984 8044
rect 20036 8072 20042 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 20036 8044 20269 8072
rect 20036 8032 20042 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 21085 8075 21143 8081
rect 21085 8072 21097 8075
rect 20257 8035 20315 8041
rect 20364 8044 21097 8072
rect 17126 8004 17132 8016
rect 17039 7976 17132 8004
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 20364 8004 20392 8044
rect 21085 8041 21097 8044
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22097 8075 22155 8081
rect 22097 8072 22109 8075
rect 21968 8044 22109 8072
rect 21968 8032 21974 8044
rect 22097 8041 22109 8044
rect 22143 8041 22155 8075
rect 22097 8035 22155 8041
rect 23750 8032 23756 8084
rect 23808 8072 23814 8084
rect 24489 8075 24547 8081
rect 24489 8072 24501 8075
rect 23808 8044 24501 8072
rect 23808 8032 23814 8044
rect 24489 8041 24501 8044
rect 24535 8041 24547 8075
rect 24489 8035 24547 8041
rect 18800 7976 20392 8004
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10192 7908 10241 7936
rect 10192 7896 10198 7908
rect 10229 7905 10241 7908
rect 10275 7936 10287 7939
rect 15657 7939 15715 7945
rect 10275 7908 11002 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 7650 7868 7656 7880
rect 7611 7840 7656 7868
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 6733 7803 6791 7809
rect 6733 7769 6745 7803
rect 6779 7800 6791 7803
rect 8110 7800 8116 7812
rect 6779 7772 8116 7800
rect 6779 7769 6791 7772
rect 6733 7763 6791 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8205 7803 8263 7809
rect 8205 7769 8217 7803
rect 8251 7769 8263 7803
rect 10974 7800 11002 7908
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 15746 7936 15752 7948
rect 15703 7908 15752 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 15933 7939 15991 7945
rect 15933 7905 15945 7939
rect 15979 7936 15991 7939
rect 16022 7936 16028 7948
rect 15979 7908 16028 7936
rect 15979 7905 15991 7908
rect 15933 7899 15991 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18800 7945 18828 7976
rect 20622 7964 20628 8016
rect 20680 8004 20686 8016
rect 21266 8004 21272 8016
rect 20680 7976 21272 8004
rect 20680 7964 20686 7976
rect 21266 7964 21272 7976
rect 21324 8004 21330 8016
rect 21361 8007 21419 8013
rect 21361 8004 21373 8007
rect 21324 7976 21373 8004
rect 21324 7964 21330 7976
rect 21361 7973 21373 7976
rect 21407 7973 21419 8007
rect 23290 8004 23296 8016
rect 23251 7976 23296 8004
rect 21361 7967 21419 7973
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 24210 8004 24216 8016
rect 24171 7976 24216 8004
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 24670 8004 24676 8016
rect 24631 7976 24676 8004
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 18785 7939 18843 7945
rect 18785 7936 18797 7939
rect 18012 7908 18797 7936
rect 18012 7896 18018 7908
rect 18785 7905 18797 7908
rect 18831 7905 18843 7939
rect 18966 7936 18972 7948
rect 18927 7908 18972 7936
rect 18785 7899 18843 7905
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 20901 7939 20959 7945
rect 20901 7905 20913 7939
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 11790 7828 11796 7840
rect 11848 7868 11854 7880
rect 12437 7871 12495 7877
rect 12437 7868 12449 7871
rect 11848 7840 12449 7868
rect 11848 7828 11854 7840
rect 12437 7837 12449 7840
rect 12483 7837 12495 7871
rect 12437 7831 12495 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13722 7868 13728 7880
rect 13495 7840 13728 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 16114 7868 16120 7880
rect 16075 7840 16120 7868
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17310 7868 17316 7880
rect 17271 7840 17316 7868
rect 17037 7831 17095 7837
rect 11882 7800 11888 7812
rect 10974 7772 11888 7800
rect 8205 7763 8263 7769
rect 5721 7735 5779 7741
rect 5721 7701 5733 7735
rect 5767 7732 5779 7735
rect 6914 7732 6920 7744
rect 5767 7704 6920 7732
rect 5767 7701 5779 7704
rect 5721 7695 5779 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 8220 7732 8248 7763
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 14826 7760 14832 7812
rect 14884 7800 14890 7812
rect 17052 7800 17080 7831
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 20916 7868 20944 7899
rect 20990 7896 20996 7948
rect 21048 7936 21054 7948
rect 21726 7936 21732 7948
rect 21048 7908 21732 7936
rect 21048 7896 21054 7908
rect 21726 7896 21732 7908
rect 21784 7896 21790 7948
rect 21913 7939 21971 7945
rect 21913 7905 21925 7939
rect 21959 7936 21971 7939
rect 22462 7936 22468 7948
rect 21959 7908 22468 7936
rect 21959 7905 21971 7908
rect 21913 7899 21971 7905
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24118 7936 24124 7948
rect 23891 7908 24124 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24118 7896 24124 7908
rect 24176 7896 24182 7948
rect 25222 7936 25228 7948
rect 25183 7908 25228 7936
rect 25222 7896 25228 7908
rect 25280 7896 25286 7948
rect 22922 7868 22928 7880
rect 20916 7840 22928 7868
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23014 7828 23020 7880
rect 23072 7868 23078 7880
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 23072 7840 23213 7868
rect 23072 7828 23078 7840
rect 23201 7837 23213 7840
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 18049 7803 18107 7809
rect 18049 7800 18061 7803
rect 14884 7772 16896 7800
rect 17052 7772 18061 7800
rect 14884 7760 14890 7772
rect 7616 7704 8248 7732
rect 7616 7692 7622 7704
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 9950 7732 9956 7744
rect 9732 7704 9956 7732
rect 9732 7692 9738 7704
rect 9950 7692 9956 7704
rect 10008 7732 10014 7744
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 10008 7704 11253 7732
rect 10008 7692 10014 7704
rect 11241 7701 11253 7704
rect 11287 7732 11299 7735
rect 11422 7732 11428 7744
rect 11287 7704 11428 7732
rect 11287 7701 11299 7704
rect 11241 7695 11299 7701
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 14734 7732 14740 7744
rect 14507 7704 14740 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 16390 7732 16396 7744
rect 16351 7704 16396 7732
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 16868 7732 16896 7772
rect 18049 7769 18061 7772
rect 18095 7800 18107 7803
rect 20990 7800 20996 7812
rect 18095 7772 20996 7800
rect 18095 7769 18107 7772
rect 18049 7763 18107 7769
rect 20990 7760 20996 7772
rect 21048 7760 21054 7812
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 16868 7704 20637 7732
rect 20625 7701 20637 7704
rect 20671 7732 20683 7735
rect 21634 7732 21640 7744
rect 20671 7704 21640 7732
rect 20671 7701 20683 7704
rect 20625 7695 20683 7701
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 22462 7732 22468 7744
rect 22423 7704 22468 7732
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6454 7528 6460 7540
rect 5951 7500 6460 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7006 7528 7012 7540
rect 6687 7500 7012 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7650 7528 7656 7540
rect 7208 7500 7656 7528
rect 7208 7401 7236 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11020 7500 11529 7528
rect 11020 7488 11026 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11664 7500 11805 7528
rect 11664 7488 11670 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 11793 7491 11851 7497
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13630 7528 13636 7540
rect 13587 7500 13636 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 13780 7500 13829 7528
rect 13780 7488 13786 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 13817 7491 13875 7497
rect 15473 7531 15531 7537
rect 15473 7497 15485 7531
rect 15519 7528 15531 7531
rect 16022 7528 16028 7540
rect 15519 7500 16028 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 11204 7432 12848 7460
rect 11204 7420 11210 7432
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 8202 7392 8208 7404
rect 8163 7364 8208 7392
rect 7193 7355 7251 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 10778 7392 10784 7404
rect 10643 7364 10784 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 12820 7401 12848 7432
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 11848 7364 12541 7392
rect 11848 7352 11854 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 14645 7327 14703 7333
rect 5767 7296 6316 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 6288 7200 6316 7296
rect 14645 7293 14657 7327
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 8110 7256 8116 7268
rect 8023 7228 8116 7256
rect 8110 7216 8116 7228
rect 8168 7256 8174 7268
rect 8567 7259 8625 7265
rect 8567 7256 8579 7259
rect 8168 7228 8579 7256
rect 8168 7216 8174 7228
rect 8567 7225 8579 7228
rect 8613 7256 8625 7259
rect 10505 7259 10563 7265
rect 10505 7256 10517 7259
rect 8613 7228 10517 7256
rect 8613 7225 8625 7228
rect 8567 7219 8625 7225
rect 10505 7225 10517 7228
rect 10551 7256 10563 7259
rect 10959 7259 11017 7265
rect 10959 7256 10971 7259
rect 10551 7228 10971 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10959 7225 10971 7228
rect 11005 7256 11017 7259
rect 12158 7256 12164 7268
rect 11005 7228 12164 7256
rect 11005 7225 11017 7228
rect 10959 7219 11017 7225
rect 12158 7216 12164 7228
rect 12216 7216 12222 7268
rect 12621 7259 12679 7265
rect 12621 7225 12633 7259
rect 12667 7225 12679 7259
rect 12621 7219 12679 7225
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6270 7188 6276 7200
rect 6231 7160 6276 7188
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 9122 7188 9128 7200
rect 9083 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9548 7160 9689 7188
rect 9548 7148 9554 7160
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12636 7188 12664 7219
rect 14182 7216 14188 7268
rect 14240 7256 14246 7268
rect 14277 7259 14335 7265
rect 14277 7256 14289 7259
rect 14240 7228 14289 7256
rect 14240 7216 14246 7228
rect 14277 7225 14289 7228
rect 14323 7256 14335 7259
rect 14660 7256 14688 7287
rect 14734 7284 14740 7336
rect 14792 7324 14798 7336
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 14792 7296 14933 7324
rect 14792 7284 14798 7296
rect 14921 7293 14933 7296
rect 14967 7324 14979 7327
rect 15488 7324 15516 7491
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 17126 7528 17132 7540
rect 17087 7500 17132 7528
rect 17126 7488 17132 7500
rect 17184 7488 17190 7540
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 17954 7528 17960 7540
rect 17911 7500 17960 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 15746 7420 15752 7472
rect 15804 7460 15810 7472
rect 15841 7463 15899 7469
rect 15841 7460 15853 7463
rect 15804 7432 15853 7460
rect 15804 7420 15810 7432
rect 15841 7429 15853 7432
rect 15887 7460 15899 7463
rect 17880 7460 17908 7491
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 18966 7528 18972 7540
rect 18555 7500 18972 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 23290 7488 23296 7540
rect 23348 7528 23354 7540
rect 24857 7531 24915 7537
rect 24857 7528 24869 7531
rect 23348 7500 24869 7528
rect 23348 7488 23354 7500
rect 24857 7497 24869 7500
rect 24903 7497 24915 7531
rect 25222 7528 25228 7540
rect 25183 7500 25228 7528
rect 24857 7491 24915 7497
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 25866 7528 25872 7540
rect 25827 7500 25872 7528
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 19058 7460 19064 7472
rect 15887 7432 17908 7460
rect 19019 7432 19064 7460
rect 15887 7429 15899 7432
rect 15841 7423 15899 7429
rect 19058 7420 19064 7432
rect 19116 7460 19122 7472
rect 19978 7460 19984 7472
rect 19116 7432 19984 7460
rect 19116 7420 19122 7432
rect 19978 7420 19984 7432
rect 20036 7460 20042 7472
rect 20349 7463 20407 7469
rect 20349 7460 20361 7463
rect 20036 7432 20361 7460
rect 20036 7420 20042 7432
rect 20349 7429 20361 7432
rect 20395 7460 20407 7463
rect 20622 7460 20628 7472
rect 20395 7432 20628 7460
rect 20395 7429 20407 7432
rect 20349 7423 20407 7429
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 21726 7420 21732 7472
rect 21784 7460 21790 7472
rect 22281 7463 22339 7469
rect 22281 7460 22293 7463
rect 21784 7432 22293 7460
rect 21784 7420 21790 7432
rect 22281 7429 22293 7432
rect 22327 7429 22339 7463
rect 22281 7423 22339 7429
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16942 7392 16948 7404
rect 16255 7364 16948 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 18690 7352 18696 7404
rect 18748 7392 18754 7404
rect 19426 7392 19432 7404
rect 18748 7364 19288 7392
rect 19387 7364 19432 7392
rect 18748 7352 18754 7364
rect 19260 7333 19288 7364
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 21358 7392 21364 7404
rect 20364 7364 21364 7392
rect 14967 7296 15516 7324
rect 18969 7327 19027 7333
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 18969 7293 18981 7327
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 19245 7327 19303 7333
rect 19245 7293 19257 7327
rect 19291 7324 19303 7327
rect 20364 7324 20392 7364
rect 20530 7324 20536 7336
rect 19291 7296 20392 7324
rect 20491 7296 20536 7324
rect 19291 7293 19303 7296
rect 19245 7287 19303 7293
rect 16301 7259 16359 7265
rect 14323 7228 15878 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 12894 7188 12900 7200
rect 12299 7160 12900 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 15850 7188 15878 7228
rect 16301 7225 16313 7259
rect 16347 7256 16359 7259
rect 16390 7256 16396 7268
rect 16347 7228 16396 7256
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 16853 7259 16911 7265
rect 16853 7225 16865 7259
rect 16899 7256 16911 7259
rect 17402 7256 17408 7268
rect 16899 7228 17408 7256
rect 16899 7225 16911 7228
rect 16853 7219 16911 7225
rect 17402 7216 17408 7228
rect 17460 7216 17466 7268
rect 18877 7259 18935 7265
rect 18877 7225 18889 7259
rect 18923 7256 18935 7259
rect 18984 7256 19012 7287
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 20824 7333 20852 7364
rect 21358 7352 21364 7364
rect 21416 7392 21422 7404
rect 21913 7395 21971 7401
rect 21913 7392 21925 7395
rect 21416 7364 21925 7392
rect 21416 7352 21422 7364
rect 21913 7361 21925 7364
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 24210 7392 24216 7404
rect 23983 7364 24216 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7293 20867 7327
rect 20809 7287 20867 7293
rect 22097 7327 22155 7333
rect 22097 7293 22109 7327
rect 22143 7324 22155 7327
rect 25476 7327 25534 7333
rect 22143 7296 22600 7324
rect 22143 7293 22155 7296
rect 22097 7287 22155 7293
rect 20070 7256 20076 7268
rect 18923 7228 20076 7256
rect 18923 7225 18935 7228
rect 18877 7219 18935 7225
rect 20070 7216 20076 7228
rect 20128 7216 20134 7268
rect 21545 7259 21603 7265
rect 21545 7256 21557 7259
rect 20548 7228 21557 7256
rect 18230 7188 18236 7200
rect 15850 7160 18236 7188
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 20548 7188 20576 7228
rect 21545 7225 21557 7228
rect 21591 7256 21603 7259
rect 21818 7256 21824 7268
rect 21591 7228 21824 7256
rect 21591 7225 21603 7228
rect 21545 7219 21603 7225
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 22572 7200 22600 7296
rect 25476 7293 25488 7327
rect 25522 7324 25534 7327
rect 25866 7324 25872 7336
rect 25522 7296 25872 7324
rect 25522 7293 25534 7296
rect 25476 7287 25534 7293
rect 25866 7284 25872 7296
rect 25924 7284 25930 7336
rect 24026 7216 24032 7268
rect 24084 7256 24090 7268
rect 24581 7259 24639 7265
rect 24084 7228 24129 7256
rect 24084 7216 24090 7228
rect 24581 7225 24593 7259
rect 24627 7256 24639 7259
rect 24670 7256 24676 7268
rect 24627 7228 24676 7256
rect 24627 7225 24639 7228
rect 24581 7219 24639 7225
rect 24670 7216 24676 7228
rect 24728 7256 24734 7268
rect 25774 7256 25780 7268
rect 24728 7228 25780 7256
rect 24728 7216 24734 7228
rect 25774 7216 25780 7228
rect 25832 7216 25838 7268
rect 20990 7188 20996 7200
rect 19116 7160 20576 7188
rect 20951 7160 20996 7188
rect 19116 7148 19122 7160
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 22554 7188 22560 7200
rect 22515 7160 22560 7188
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 22922 7188 22928 7200
rect 22883 7160 22928 7188
rect 22922 7148 22928 7160
rect 22980 7148 22986 7200
rect 23477 7191 23535 7197
rect 23477 7157 23489 7191
rect 23523 7188 23535 7191
rect 24044 7188 24072 7216
rect 23523 7160 24072 7188
rect 23523 7157 23535 7160
rect 23477 7151 23535 7157
rect 25314 7148 25320 7200
rect 25372 7188 25378 7200
rect 25547 7191 25605 7197
rect 25547 7188 25559 7191
rect 25372 7160 25559 7188
rect 25372 7148 25378 7160
rect 25547 7157 25559 7160
rect 25593 7157 25605 7191
rect 25547 7151 25605 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 7742 6984 7748 6996
rect 7699 6956 7748 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 7742 6944 7748 6956
rect 7800 6984 7806 6996
rect 7800 6956 8064 6984
rect 7800 6944 7806 6956
rect 6457 6919 6515 6925
rect 6457 6885 6469 6919
rect 6503 6916 6515 6919
rect 6546 6916 6552 6928
rect 6503 6888 6552 6916
rect 6503 6885 6515 6888
rect 6457 6879 6515 6885
rect 6546 6876 6552 6888
rect 6604 6916 6610 6928
rect 8036 6916 8064 6956
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 8168 6956 8217 6984
rect 8168 6944 8174 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8352 6956 9045 6984
rect 8352 6944 8358 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 9033 6947 9091 6953
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12308 6956 12357 6984
rect 12308 6944 12314 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12894 6984 12900 6996
rect 12855 6956 12900 6984
rect 12345 6947 12403 6953
rect 8386 6916 8392 6928
rect 6604 6888 7742 6916
rect 8036 6888 8392 6916
rect 6604 6876 6610 6888
rect 7714 6848 7742 6888
rect 8386 6876 8392 6888
rect 8444 6916 8450 6928
rect 8849 6919 8907 6925
rect 8849 6916 8861 6919
rect 8444 6888 8861 6916
rect 8444 6876 8450 6888
rect 8849 6885 8861 6888
rect 8895 6885 8907 6919
rect 10321 6919 10379 6925
rect 10321 6916 10333 6919
rect 8849 6879 8907 6885
rect 9646 6888 10333 6916
rect 9398 6848 9404 6860
rect 7714 6820 9404 6848
rect 9398 6808 9404 6820
rect 9456 6848 9462 6860
rect 9646 6848 9674 6888
rect 10321 6885 10333 6888
rect 10367 6916 10379 6919
rect 10686 6916 10692 6928
rect 10367 6888 10692 6916
rect 10367 6885 10379 6888
rect 10321 6879 10379 6885
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 12360 6916 12388 6947
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 14645 6987 14703 6993
rect 14645 6953 14657 6987
rect 14691 6984 14703 6987
rect 15654 6984 15660 6996
rect 14691 6956 15660 6984
rect 14691 6953 14703 6956
rect 14645 6947 14703 6953
rect 14660 6916 14688 6947
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16114 6944 16120 6996
rect 16172 6984 16178 6996
rect 16485 6987 16543 6993
rect 16485 6984 16497 6987
rect 16172 6956 16497 6984
rect 16172 6944 16178 6956
rect 16485 6953 16497 6956
rect 16531 6953 16543 6987
rect 18690 6984 18696 6996
rect 16485 6947 16543 6953
rect 17052 6956 18552 6984
rect 18651 6956 18696 6984
rect 12360 6888 14688 6916
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 17052 6916 17080 6956
rect 17218 6916 17224 6928
rect 14792 6888 17080 6916
rect 17179 6888 17224 6916
rect 14792 6876 14798 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 13998 6848 14004 6860
rect 9456 6820 9674 6848
rect 13959 6820 14004 6848
rect 9456 6808 9462 6820
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 18524 6848 18552 6956
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 20530 6984 20536 6996
rect 20491 6956 20536 6984
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 23566 6984 23572 6996
rect 23527 6956 23572 6984
rect 23566 6944 23572 6956
rect 23624 6944 23630 6996
rect 18966 6876 18972 6928
rect 19024 6916 19030 6928
rect 19198 6919 19256 6925
rect 19198 6916 19210 6919
rect 19024 6888 19210 6916
rect 19024 6876 19030 6888
rect 19198 6885 19210 6888
rect 19244 6885 19256 6919
rect 19198 6879 19256 6885
rect 19794 6848 19800 6860
rect 18524 6820 19800 6848
rect 19794 6808 19800 6820
rect 19852 6848 19858 6860
rect 20073 6851 20131 6857
rect 20073 6848 20085 6851
rect 19852 6820 20085 6848
rect 19852 6808 19858 6820
rect 20073 6817 20085 6820
rect 20119 6848 20131 6851
rect 20254 6848 20260 6860
rect 20119 6820 20260 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 20254 6808 20260 6820
rect 20312 6848 20318 6860
rect 20806 6848 20812 6860
rect 20312 6820 20812 6848
rect 20312 6808 20318 6820
rect 20806 6808 20812 6820
rect 20864 6848 20870 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20864 6820 20913 6848
rect 20864 6808 20870 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 21266 6808 21272 6860
rect 21324 6848 21330 6860
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 21324 6820 21373 6848
rect 21324 6808 21330 6820
rect 21361 6817 21373 6820
rect 21407 6817 21419 6851
rect 21726 6848 21732 6860
rect 21687 6820 21732 6848
rect 21361 6811 21419 6817
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 21818 6808 21824 6860
rect 21876 6848 21882 6860
rect 22097 6851 22155 6857
rect 22097 6848 22109 6851
rect 21876 6820 22109 6848
rect 21876 6808 21882 6820
rect 22097 6817 22109 6820
rect 22143 6817 22155 6851
rect 22097 6811 22155 6817
rect 22186 6808 22192 6860
rect 22244 6848 22250 6860
rect 24949 6851 25007 6857
rect 24949 6848 24961 6851
rect 22244 6820 24961 6848
rect 22244 6808 22250 6820
rect 24949 6817 24961 6820
rect 24995 6848 25007 6851
rect 25038 6848 25044 6860
rect 24995 6820 25044 6848
rect 24995 6817 25007 6820
rect 24949 6811 25007 6817
rect 25038 6808 25044 6820
rect 25096 6808 25102 6860
rect 5166 6780 5172 6792
rect 5127 6752 5172 6780
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6454 6780 6460 6792
rect 6411 6752 6460 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7558 6780 7564 6792
rect 7055 6752 7564 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10502 6780 10508 6792
rect 10463 6752 10508 6780
rect 10229 6743 10287 6749
rect 5399 6715 5457 6721
rect 5399 6681 5411 6715
rect 5445 6712 5457 6715
rect 5445 6684 10088 6712
rect 5445 6681 5457 6684
rect 5399 6675 5457 6681
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 8846 6644 8852 6656
rect 7800 6616 8852 6644
rect 7800 6604 7806 6616
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9858 6644 9864 6656
rect 9819 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 10060 6644 10088 6684
rect 10134 6672 10140 6724
rect 10192 6712 10198 6724
rect 10244 6712 10272 6743
rect 10502 6740 10508 6752
rect 10560 6780 10566 6792
rect 11790 6780 11796 6792
rect 10560 6752 11796 6780
rect 10560 6740 10566 6752
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12526 6780 12532 6792
rect 12023 6752 12532 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6749 17187 6783
rect 17402 6780 17408 6792
rect 17363 6752 17408 6780
rect 17129 6743 17187 6749
rect 10192 6684 10272 6712
rect 14185 6715 14243 6721
rect 10192 6672 10198 6684
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 14826 6712 14832 6724
rect 14231 6684 14832 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 17144 6712 17172 6743
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 18877 6783 18935 6789
rect 17552 6752 18321 6780
rect 17552 6740 17558 6752
rect 17770 6712 17776 6724
rect 17144 6684 17776 6712
rect 17770 6672 17776 6684
rect 17828 6672 17834 6724
rect 18293 6712 18321 6752
rect 18877 6749 18889 6783
rect 18923 6780 18935 6783
rect 19426 6780 19432 6792
rect 18923 6752 19432 6780
rect 18923 6749 18935 6752
rect 18877 6743 18935 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6780 22431 6783
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 22419 6752 23213 6780
rect 22419 6749 22431 6752
rect 22373 6743 22431 6749
rect 23201 6749 23213 6752
rect 23247 6780 23259 6783
rect 23290 6780 23296 6792
rect 23247 6752 23296 6780
rect 23247 6749 23259 6752
rect 23201 6743 23259 6749
rect 23290 6740 23296 6752
rect 23348 6740 23354 6792
rect 25406 6712 25412 6724
rect 18293 6684 25412 6712
rect 25406 6672 25412 6684
rect 25464 6672 25470 6724
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10060 6616 11437 6644
rect 11425 6613 11437 6616
rect 11471 6644 11483 6647
rect 11514 6644 11520 6656
rect 11471 6616 11520 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 15930 6644 15936 6656
rect 11664 6616 15936 6644
rect 11664 6604 11670 6616
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16390 6644 16396 6656
rect 16255 6616 16396 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16390 6604 16396 6616
rect 16448 6604 16454 6656
rect 16942 6644 16948 6656
rect 16855 6616 16948 6644
rect 16942 6604 16948 6616
rect 17000 6644 17006 6656
rect 18046 6644 18052 6656
rect 17000 6616 18052 6644
rect 17000 6604 17006 6616
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 19518 6604 19524 6656
rect 19576 6644 19582 6656
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 19576 6616 19809 6644
rect 19576 6604 19582 6616
rect 19797 6613 19809 6616
rect 19843 6613 19855 6647
rect 19797 6607 19855 6613
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 22649 6647 22707 6653
rect 22649 6644 22661 6647
rect 22060 6616 22661 6644
rect 22060 6604 22066 6616
rect 22649 6613 22661 6616
rect 22695 6613 22707 6647
rect 23014 6644 23020 6656
rect 22975 6616 23020 6644
rect 22649 6607 22707 6613
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 24121 6647 24179 6653
rect 24121 6613 24133 6647
rect 24167 6644 24179 6647
rect 24210 6644 24216 6656
rect 24167 6616 24216 6644
rect 24167 6613 24179 6616
rect 24121 6607 24179 6613
rect 24210 6604 24216 6616
rect 24268 6644 24274 6656
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 24268 6616 24409 6644
rect 24268 6604 24274 6616
rect 24397 6613 24409 6616
rect 24443 6613 24455 6647
rect 24397 6607 24455 6613
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 25087 6647 25145 6653
rect 25087 6644 25099 6647
rect 24820 6616 25099 6644
rect 24820 6604 24826 6616
rect 25087 6613 25099 6616
rect 25133 6613 25145 6647
rect 25087 6607 25145 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 7098 6440 7104 6452
rect 4939 6412 7104 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7892 6412 8309 6440
rect 7892 6400 7898 6412
rect 8297 6409 8309 6412
rect 8343 6440 8355 6443
rect 9766 6440 9772 6452
rect 8343 6412 9772 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10744 6412 10885 6440
rect 10744 6400 10750 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 12250 6440 12256 6452
rect 12115 6412 12256 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 17494 6440 17500 6452
rect 14148 6412 17500 6440
rect 14148 6400 14154 6412
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18966 6440 18972 6452
rect 18927 6412 18972 6440
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 25038 6440 25044 6452
rect 24999 6412 25044 6440
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6372 4675 6375
rect 4706 6372 4712 6384
rect 4663 6344 4712 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 5859 6375 5917 6381
rect 5859 6341 5871 6375
rect 5905 6372 5917 6375
rect 9858 6372 9864 6384
rect 5905 6344 9864 6372
rect 5905 6341 5917 6344
rect 5859 6335 5917 6341
rect 9858 6332 9864 6344
rect 9916 6372 9922 6384
rect 10502 6372 10508 6384
rect 9916 6344 9996 6372
rect 10463 6344 10508 6372
rect 9916 6332 9922 6344
rect 4724 6245 4752 6332
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 5224 6276 5365 6304
rect 5224 6264 5230 6276
rect 5353 6273 5365 6276
rect 5399 6304 5411 6307
rect 5994 6304 6000 6316
rect 5399 6276 6000 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6546 6304 6552 6316
rect 6507 6276 6552 6304
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7374 6304 7380 6316
rect 6963 6276 7380 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7558 6304 7564 6316
rect 7519 6276 7564 6304
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8110 6304 8116 6316
rect 7975 6276 8116 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 9968 6313 9996 6344
rect 10502 6332 10508 6344
rect 10560 6332 10566 6384
rect 15838 6332 15844 6384
rect 15896 6372 15902 6384
rect 18187 6375 18245 6381
rect 18187 6372 18199 6375
rect 15896 6344 18199 6372
rect 15896 6332 15902 6344
rect 18187 6341 18199 6344
rect 18233 6341 18245 6375
rect 18187 6335 18245 6341
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 8444 6276 9689 6304
rect 8444 6264 8450 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 11882 6304 11888 6316
rect 11747 6276 11888 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 5788 6239 5846 6245
rect 5788 6205 5800 6239
rect 5834 6236 5846 6239
rect 8662 6236 8668 6248
rect 5834 6208 6316 6236
rect 5834 6205 5846 6208
rect 5788 6199 5846 6205
rect 6288 6112 6316 6208
rect 7576 6208 8668 6236
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 7009 6171 7067 6177
rect 7009 6168 7021 6171
rect 6972 6140 7021 6168
rect 6972 6128 6978 6140
rect 7009 6137 7021 6140
rect 7055 6168 7067 6171
rect 7576 6168 7604 6208
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 8884 6239 8942 6245
rect 8884 6205 8896 6239
rect 8930 6205 8942 6239
rect 8884 6199 8942 6205
rect 8987 6239 9045 6245
rect 8987 6205 8999 6239
rect 9033 6236 9045 6239
rect 9582 6236 9588 6248
rect 9033 6208 9588 6236
rect 9033 6205 9045 6208
rect 8987 6199 9045 6205
rect 7055 6140 7604 6168
rect 7055 6137 7067 6140
rect 7009 6131 7067 6137
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 8899 6168 8927 6199
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9692 6180 9720 6267
rect 11882 6264 11888 6276
rect 11940 6304 11946 6316
rect 13725 6307 13783 6313
rect 11940 6276 12664 6304
rect 11940 6264 11946 6276
rect 12434 6236 12440 6248
rect 12395 6208 12440 6236
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12636 6236 12664 6276
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13771 6276 14381 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14369 6273 14381 6276
rect 14415 6304 14427 6307
rect 14458 6304 14464 6316
rect 14415 6276 14464 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 18984 6304 19012 6400
rect 20898 6332 20904 6384
rect 20956 6372 20962 6384
rect 24305 6375 24363 6381
rect 20956 6344 23474 6372
rect 20956 6332 20962 6344
rect 17414 6276 19012 6304
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 12636 6208 12909 6236
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6236 15347 6239
rect 15562 6236 15568 6248
rect 15335 6208 15568 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 15562 6196 15568 6208
rect 15620 6236 15626 6248
rect 17218 6236 17224 6248
rect 15620 6208 17224 6236
rect 15620 6196 15626 6208
rect 17218 6196 17224 6208
rect 17276 6236 17282 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 17276 6208 17325 6236
rect 17276 6196 17282 6208
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 9398 6168 9404 6180
rect 7708 6140 9404 6168
rect 7708 6128 7714 6140
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 9674 6168 9680 6180
rect 9587 6140 9680 6168
rect 9674 6128 9680 6140
rect 9732 6168 9738 6180
rect 10045 6171 10103 6177
rect 10045 6168 10057 6171
rect 9732 6140 10057 6168
rect 9732 6128 9738 6140
rect 10045 6137 10057 6140
rect 10091 6137 10103 6171
rect 10045 6131 10103 6137
rect 11333 6171 11391 6177
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 14731 6171 14789 6177
rect 11379 6140 12572 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 12544 6112 12572 6140
rect 14731 6137 14743 6171
rect 14777 6168 14789 6171
rect 15654 6168 15660 6180
rect 14777 6140 15660 6168
rect 14777 6137 14789 6140
rect 14731 6131 14789 6137
rect 15654 6128 15660 6140
rect 15712 6168 15718 6180
rect 16025 6171 16083 6177
rect 16025 6168 16037 6171
rect 15712 6140 16037 6168
rect 15712 6128 15718 6140
rect 16025 6137 16037 6140
rect 16071 6168 16083 6171
rect 16479 6171 16537 6177
rect 16479 6168 16491 6171
rect 16071 6140 16491 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 16479 6137 16491 6140
rect 16525 6168 16537 6171
rect 17414 6168 17442 6276
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 21269 6307 21327 6313
rect 21269 6304 21281 6307
rect 19208 6276 21281 6304
rect 19208 6264 19214 6276
rect 18116 6239 18174 6245
rect 18116 6205 18128 6239
rect 18162 6236 18174 6239
rect 19794 6236 19800 6248
rect 18162 6208 18644 6236
rect 19755 6208 19800 6236
rect 18162 6205 18174 6208
rect 18116 6199 18174 6205
rect 16525 6140 17442 6168
rect 16525 6137 16537 6140
rect 16479 6131 16537 6137
rect 6270 6100 6276 6112
rect 6231 6072 6276 6100
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 11238 6100 11244 6112
rect 8628 6072 11244 6100
rect 8628 6060 8634 6072
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 12526 6100 12532 6112
rect 12487 6072 12532 6100
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 18616 6109 18644 6208
rect 19794 6196 19800 6208
rect 19852 6196 19858 6248
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 20364 6245 20392 6276
rect 21269 6273 21281 6276
rect 21315 6304 21327 6307
rect 21726 6304 21732 6316
rect 21315 6276 21732 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 22462 6304 22468 6316
rect 22423 6276 22468 6304
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 23446 6304 23474 6344
rect 24305 6341 24317 6375
rect 24351 6372 24363 6375
rect 24670 6372 24676 6384
rect 24351 6344 24676 6372
rect 24351 6341 24363 6344
rect 24305 6335 24363 6341
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 23446 6276 24859 6304
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6205 20407 6239
rect 20349 6199 20407 6205
rect 20717 6239 20775 6245
rect 20717 6205 20729 6239
rect 20763 6205 20775 6239
rect 22002 6236 22008 6248
rect 21963 6208 22008 6236
rect 20717 6199 20775 6205
rect 20732 6168 20760 6199
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22281 6239 22339 6245
rect 22152 6208 22197 6236
rect 22152 6196 22158 6208
rect 22281 6205 22293 6239
rect 22327 6236 22339 6239
rect 22370 6236 22376 6248
rect 22327 6208 22376 6236
rect 22327 6205 22339 6208
rect 22281 6199 22339 6205
rect 21174 6168 21180 6180
rect 19352 6140 21180 6168
rect 19352 6112 19380 6140
rect 21174 6128 21180 6140
rect 21232 6128 21238 6180
rect 21913 6171 21971 6177
rect 21913 6137 21925 6171
rect 21959 6168 21971 6171
rect 22296 6168 22324 6199
rect 22370 6196 22376 6208
rect 22428 6196 22434 6248
rect 24831 6236 24859 6276
rect 25260 6239 25318 6245
rect 25260 6236 25272 6239
rect 24831 6208 25272 6236
rect 25260 6205 25272 6208
rect 25306 6236 25318 6239
rect 25685 6239 25743 6245
rect 25685 6236 25697 6239
rect 25306 6208 25697 6236
rect 25306 6205 25318 6208
rect 25260 6199 25318 6205
rect 25685 6205 25697 6208
rect 25731 6205 25743 6239
rect 25685 6199 25743 6205
rect 23750 6168 23756 6180
rect 21959 6140 22324 6168
rect 23711 6140 23756 6168
rect 21959 6137 21971 6140
rect 21913 6131 21971 6137
rect 23750 6128 23756 6140
rect 23808 6128 23814 6180
rect 23845 6171 23903 6177
rect 23845 6137 23857 6171
rect 23891 6168 23903 6171
rect 24210 6168 24216 6180
rect 23891 6140 24216 6168
rect 23891 6137 23903 6140
rect 23845 6131 23903 6137
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 27246 6168 27252 6180
rect 24831 6140 27252 6168
rect 18601 6103 18659 6109
rect 18601 6069 18613 6103
rect 18647 6100 18659 6103
rect 18690 6100 18696 6112
rect 18647 6072 18696 6100
rect 18647 6069 18659 6072
rect 18601 6063 18659 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19334 6100 19340 6112
rect 19295 6072 19340 6100
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19426 6060 19432 6112
rect 19484 6100 19490 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19484 6072 19625 6100
rect 19484 6060 19490 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 19613 6063 19671 6069
rect 23293 6103 23351 6109
rect 23293 6069 23305 6103
rect 23339 6100 23351 6103
rect 23566 6100 23572 6112
rect 23339 6072 23572 6100
rect 23339 6069 23351 6072
rect 23293 6063 23351 6069
rect 23566 6060 23572 6072
rect 23624 6100 23630 6112
rect 24831 6100 24859 6140
rect 27246 6128 27252 6140
rect 27304 6128 27310 6180
rect 23624 6072 24859 6100
rect 23624 6060 23630 6072
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 25363 6103 25421 6109
rect 25363 6100 25375 6103
rect 25096 6072 25375 6100
rect 25096 6060 25102 6072
rect 25363 6069 25375 6072
rect 25409 6069 25421 6103
rect 25363 6063 25421 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7147 5899 7205 5905
rect 7147 5865 7159 5899
rect 7193 5896 7205 5899
rect 10134 5896 10140 5908
rect 7193 5868 10140 5896
rect 7193 5865 7205 5868
rect 7147 5859 7205 5865
rect 10134 5856 10140 5868
rect 10192 5896 10198 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10192 5868 10701 5896
rect 10192 5856 10198 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 10689 5859 10747 5865
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 12492 5868 12725 5896
rect 12492 5856 12498 5868
rect 12713 5865 12725 5868
rect 12759 5896 12771 5899
rect 13078 5896 13084 5908
rect 12759 5868 13084 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 16393 5899 16451 5905
rect 16393 5896 16405 5899
rect 16080 5868 16405 5896
rect 16080 5856 16086 5868
rect 16393 5865 16405 5868
rect 16439 5896 16451 5899
rect 16574 5896 16580 5908
rect 16439 5868 16580 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 16942 5896 16948 5908
rect 16776 5868 16948 5896
rect 5258 5828 5264 5840
rect 5067 5800 5264 5828
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 5067 5769 5095 5800
rect 5258 5788 5264 5800
rect 5316 5828 5322 5840
rect 7650 5828 7656 5840
rect 5316 5800 7656 5828
rect 5316 5788 5322 5800
rect 7650 5788 7656 5800
rect 7708 5788 7714 5840
rect 8205 5831 8263 5837
rect 8205 5797 8217 5831
rect 8251 5828 8263 5831
rect 8386 5828 8392 5840
rect 8251 5800 8392 5828
rect 8251 5797 8263 5800
rect 8205 5791 8263 5797
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 8938 5828 8944 5840
rect 8803 5800 8944 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 9180 5800 9873 5828
rect 9180 5788 9186 5800
rect 9861 5797 9873 5800
rect 9907 5828 9919 5831
rect 10042 5828 10048 5840
rect 9907 5800 10048 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 11882 5828 11888 5840
rect 11843 5800 11888 5828
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 14734 5828 14740 5840
rect 14108 5800 14740 5828
rect 5052 5763 5110 5769
rect 5052 5729 5064 5763
rect 5098 5729 5110 5763
rect 5994 5760 6000 5772
rect 5955 5732 6000 5760
rect 5052 5723 5110 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 7044 5763 7102 5769
rect 7044 5760 7056 5763
rect 6696 5732 7056 5760
rect 6696 5720 6702 5732
rect 7044 5729 7056 5732
rect 7090 5729 7102 5763
rect 7044 5723 7102 5729
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 11146 5760 11152 5772
rect 10468 5732 11152 5760
rect 10468 5720 10474 5732
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 13909 5763 13967 5769
rect 13909 5729 13921 5763
rect 13955 5760 13967 5763
rect 13998 5760 14004 5772
rect 13955 5732 14004 5760
rect 13955 5729 13967 5732
rect 13909 5723 13967 5729
rect 13998 5720 14004 5732
rect 14056 5720 14062 5772
rect 14108 5769 14136 5800
rect 14734 5788 14740 5800
rect 14792 5828 14798 5840
rect 16040 5828 16068 5856
rect 16776 5837 16804 5868
rect 16942 5856 16948 5868
rect 17000 5896 17006 5908
rect 17310 5896 17316 5908
rect 17000 5868 17316 5896
rect 17000 5856 17006 5868
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 18417 5899 18475 5905
rect 18417 5865 18429 5899
rect 18463 5896 18475 5899
rect 19426 5896 19432 5908
rect 18463 5868 19432 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 19978 5896 19984 5908
rect 19939 5868 19984 5896
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20070 5856 20076 5908
rect 20128 5896 20134 5908
rect 22649 5899 22707 5905
rect 22649 5896 22661 5899
rect 20128 5868 22661 5896
rect 20128 5856 20134 5868
rect 22649 5865 22661 5868
rect 22695 5865 22707 5899
rect 23290 5896 23296 5908
rect 23251 5868 23296 5896
rect 22649 5859 22707 5865
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 24026 5896 24032 5908
rect 23987 5868 24032 5896
rect 24026 5856 24032 5868
rect 24084 5856 24090 5908
rect 14792 5800 16068 5828
rect 16761 5831 16819 5837
rect 14792 5788 14798 5800
rect 16761 5797 16773 5831
rect 16807 5797 16819 5831
rect 16761 5791 16819 5797
rect 16853 5831 16911 5837
rect 16853 5797 16865 5831
rect 16899 5828 16911 5831
rect 17034 5828 17040 5840
rect 16899 5800 17040 5828
rect 16899 5797 16911 5800
rect 16853 5791 16911 5797
rect 17034 5788 17040 5800
rect 17092 5828 17098 5840
rect 17402 5828 17408 5840
rect 17092 5800 17408 5828
rect 17092 5788 17098 5800
rect 17402 5788 17408 5800
rect 17460 5788 17466 5840
rect 18598 5788 18604 5840
rect 18656 5828 18662 5840
rect 18693 5831 18751 5837
rect 18693 5828 18705 5831
rect 18656 5800 18705 5828
rect 18656 5788 18662 5800
rect 18693 5797 18705 5800
rect 18739 5797 18751 5831
rect 18693 5791 18751 5797
rect 19242 5788 19248 5840
rect 19300 5828 19306 5840
rect 19521 5831 19579 5837
rect 19521 5828 19533 5831
rect 19300 5800 19533 5828
rect 19300 5788 19306 5800
rect 19521 5797 19533 5800
rect 19567 5797 19579 5831
rect 19996 5828 20024 5856
rect 20625 5831 20683 5837
rect 20625 5828 20637 5831
rect 19996 5800 20637 5828
rect 19521 5791 19579 5797
rect 20625 5797 20637 5800
rect 20671 5797 20683 5831
rect 20625 5791 20683 5797
rect 21450 5788 21456 5840
rect 21508 5828 21514 5840
rect 23842 5828 23848 5840
rect 21508 5800 23848 5828
rect 21508 5788 21514 5800
rect 23842 5788 23848 5800
rect 23900 5788 23906 5840
rect 24118 5788 24124 5840
rect 24176 5828 24182 5840
rect 24176 5800 24394 5828
rect 24176 5788 24182 5800
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15378 5760 15384 5772
rect 15335 5732 15384 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 21358 5760 21364 5772
rect 21319 5732 21364 5760
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 24210 5760 24216 5772
rect 24171 5732 24216 5760
rect 24210 5720 24216 5732
rect 24268 5720 24274 5772
rect 24366 5760 24394 5800
rect 25200 5763 25258 5769
rect 25200 5760 25212 5763
rect 24366 5732 25212 5760
rect 25200 5729 25212 5732
rect 25246 5760 25258 5763
rect 25774 5760 25780 5772
rect 25246 5732 25780 5760
rect 25246 5729 25258 5732
rect 25200 5723 25258 5729
rect 25774 5720 25780 5732
rect 25832 5720 25838 5772
rect 1535 5695 1593 5701
rect 1535 5661 1547 5695
rect 1581 5692 1593 5695
rect 7834 5692 7840 5704
rect 1581 5664 7840 5692
rect 1581 5661 1593 5664
rect 1535 5655 1593 5661
rect 7834 5652 7840 5664
rect 7892 5692 7898 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7892 5664 8125 5692
rect 7892 5652 7898 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 8113 5655 8171 5661
rect 8541 5664 9413 5692
rect 6135 5627 6193 5633
rect 6135 5593 6147 5627
rect 6181 5624 6193 5627
rect 6730 5624 6736 5636
rect 6181 5596 6736 5624
rect 6181 5593 6193 5596
rect 6135 5587 6193 5593
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 8541 5624 8569 5664
rect 9401 5661 9413 5664
rect 9447 5692 9459 5695
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9447 5664 9781 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 10870 5692 10876 5704
rect 10192 5664 10876 5692
rect 10192 5652 10198 5664
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11790 5692 11796 5704
rect 11751 5664 11796 5692
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5692 12495 5695
rect 13538 5692 13544 5704
rect 12483 5664 13544 5692
rect 12483 5661 12495 5664
rect 12437 5655 12495 5661
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 14182 5692 14188 5704
rect 14143 5664 14188 5692
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19610 5692 19616 5704
rect 19291 5664 19616 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 7616 5596 8569 5624
rect 8817 5596 9254 5624
rect 7616 5584 7622 5596
rect 5123 5559 5181 5565
rect 5123 5525 5135 5559
rect 5169 5556 5181 5559
rect 6270 5556 6276 5568
rect 5169 5528 6276 5556
rect 5169 5525 5181 5528
rect 5123 5519 5181 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6454 5556 6460 5568
rect 6415 5528 6460 5556
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 7469 5559 7527 5565
rect 7469 5556 7481 5559
rect 7432 5528 7481 5556
rect 7432 5516 7438 5528
rect 7469 5525 7481 5528
rect 7515 5525 7527 5559
rect 7469 5519 7527 5525
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 8817 5556 8845 5596
rect 9122 5556 9128 5568
rect 7708 5528 8845 5556
rect 9083 5528 9128 5556
rect 7708 5516 7714 5528
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9226 5556 9254 5596
rect 12526 5584 12532 5636
rect 12584 5624 12590 5636
rect 15286 5624 15292 5636
rect 12584 5596 15292 5624
rect 12584 5584 12590 5596
rect 15286 5584 15292 5596
rect 15344 5624 15350 5636
rect 15841 5627 15899 5633
rect 15841 5624 15853 5627
rect 15344 5596 15853 5624
rect 15344 5584 15350 5596
rect 15841 5593 15853 5596
rect 15887 5593 15899 5627
rect 15841 5587 15899 5593
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 17052 5624 17080 5655
rect 16724 5596 17080 5624
rect 16724 5584 16730 5596
rect 11422 5556 11428 5568
rect 9226 5528 11428 5556
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 15654 5556 15660 5568
rect 15519 5528 15660 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 17954 5556 17960 5568
rect 17915 5528 17960 5556
rect 17954 5516 17960 5528
rect 18012 5556 18018 5568
rect 18616 5556 18644 5655
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 23017 5695 23075 5701
rect 23017 5661 23029 5695
rect 23063 5692 23075 5695
rect 23658 5692 23664 5704
rect 23063 5664 23664 5692
rect 23063 5661 23075 5664
rect 23017 5655 23075 5661
rect 23658 5652 23664 5664
rect 23716 5652 23722 5704
rect 23750 5652 23756 5704
rect 23808 5692 23814 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23808 5664 24593 5692
rect 23808 5652 23814 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 25271 5627 25329 5633
rect 25271 5624 25283 5627
rect 23446 5596 25283 5624
rect 18012 5528 18644 5556
rect 21361 5559 21419 5565
rect 18012 5516 18018 5528
rect 21361 5525 21373 5559
rect 21407 5556 21419 5559
rect 21450 5556 21456 5568
rect 21407 5528 21456 5556
rect 21407 5525 21419 5528
rect 21361 5519 21419 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 22094 5556 22100 5568
rect 22055 5528 22100 5556
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 23446 5556 23474 5596
rect 25271 5593 25283 5596
rect 25317 5593 25329 5627
rect 25271 5587 25329 5593
rect 22796 5528 23474 5556
rect 22796 5516 22802 5528
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 3283 5355 3341 5361
rect 3283 5321 3295 5355
rect 3329 5352 3341 5355
rect 6454 5352 6460 5364
rect 3329 5324 6460 5352
rect 3329 5321 3341 5324
rect 3283 5315 3341 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7190 5352 7196 5364
rect 6604 5324 7196 5352
rect 6604 5312 6610 5324
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 8168 5324 8309 5352
rect 8168 5312 8174 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 9674 5352 9680 5364
rect 9635 5324 9680 5352
rect 8297 5315 8355 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10042 5352 10048 5364
rect 10003 5324 10048 5352
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15436 5324 15577 5352
rect 15436 5312 15442 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 15565 5315 15623 5321
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5352 17926 5364
rect 17920 5324 18920 5352
rect 17920 5312 17926 5324
rect 5258 5284 5264 5296
rect 5219 5256 5264 5284
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 6273 5287 6331 5293
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 6362 5284 6368 5296
rect 6319 5256 6368 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 6288 5216 6316 5247
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 9950 5284 9956 5296
rect 7524 5256 9956 5284
rect 7524 5244 7530 5256
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 13633 5287 13691 5293
rect 13633 5284 13645 5287
rect 11256 5256 13645 5284
rect 5787 5188 6316 5216
rect 5787 5157 5815 5188
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 9490 5216 9496 5228
rect 6512 5188 9496 5216
rect 6512 5176 6518 5188
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 11256 5160 11284 5256
rect 13633 5253 13645 5256
rect 13679 5284 13691 5287
rect 14734 5284 14740 5296
rect 13679 5256 14740 5284
rect 13679 5253 13691 5256
rect 13633 5247 13691 5253
rect 14734 5244 14740 5256
rect 14792 5244 14798 5296
rect 15930 5244 15936 5296
rect 15988 5284 15994 5296
rect 18782 5284 18788 5296
rect 15988 5256 18788 5284
rect 15988 5244 15994 5256
rect 18782 5244 18788 5256
rect 18840 5244 18846 5296
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 12526 5216 12532 5228
rect 11563 5188 12532 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 18892 5225 18920 5324
rect 19058 5312 19064 5364
rect 19116 5352 19122 5364
rect 19797 5355 19855 5361
rect 19797 5352 19809 5355
rect 19116 5324 19809 5352
rect 19116 5312 19122 5324
rect 19797 5321 19809 5324
rect 19843 5352 19855 5355
rect 19978 5352 19984 5364
rect 19843 5324 19984 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 21358 5352 21364 5364
rect 20456 5324 21364 5352
rect 20456 5296 20484 5324
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22520 5324 23029 5352
rect 22520 5312 22526 5324
rect 23017 5321 23029 5324
rect 23063 5352 23075 5355
rect 23063 5324 23474 5352
rect 23063 5321 23075 5324
rect 23017 5315 23075 5321
rect 20438 5284 20444 5296
rect 20351 5256 20444 5284
rect 20438 5244 20444 5256
rect 20496 5244 20502 5296
rect 18877 5219 18935 5225
rect 18877 5185 18889 5219
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 21913 5219 21971 5225
rect 21913 5185 21925 5219
rect 21959 5216 21971 5219
rect 22554 5216 22560 5228
rect 21959 5188 22140 5216
rect 22515 5188 22560 5216
rect 21959 5185 21971 5188
rect 21913 5179 21971 5185
rect 22112 5160 22140 5188
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 23446 5216 23474 5324
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 25041 5355 25099 5361
rect 25041 5352 25053 5355
rect 24268 5324 25053 5352
rect 24268 5312 24274 5324
rect 25041 5321 25053 5324
rect 25087 5321 25099 5355
rect 25041 5315 25099 5321
rect 23842 5244 23848 5296
rect 23900 5284 23906 5296
rect 26510 5284 26516 5296
rect 23900 5256 26516 5284
rect 23900 5244 23906 5256
rect 26510 5244 26516 5256
rect 26568 5244 26574 5296
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 23446 5188 24133 5216
rect 24121 5185 24133 5188
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 3212 5151 3270 5157
rect 3212 5117 3224 5151
rect 3258 5148 3270 5151
rect 4776 5151 4834 5157
rect 3258 5120 3740 5148
rect 3258 5117 3270 5120
rect 3212 5111 3270 5117
rect 3712 5024 3740 5120
rect 4776 5117 4788 5151
rect 4822 5148 4834 5151
rect 5772 5151 5830 5157
rect 4822 5120 5488 5148
rect 4822 5117 4834 5120
rect 4776 5111 4834 5117
rect 5460 5024 5488 5120
rect 5772 5117 5784 5151
rect 5818 5117 5830 5151
rect 5772 5111 5830 5117
rect 5859 5151 5917 5157
rect 5859 5117 5871 5151
rect 5905 5148 5917 5151
rect 6178 5148 6184 5160
rect 5905 5120 6184 5148
rect 5905 5117 5917 5120
rect 5859 5111 5917 5117
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 7024 5080 7052 5111
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 7156 5120 7389 5148
rect 7156 5108 7162 5120
rect 7377 5117 7389 5120
rect 7423 5148 7435 5151
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7423 5120 7941 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7929 5117 7941 5120
rect 7975 5148 7987 5151
rect 8294 5148 8300 5160
rect 7975 5120 8300 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 8478 5148 8484 5160
rect 8439 5120 8484 5148
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 10962 5148 10968 5160
rect 10735 5120 10968 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11238 5148 11244 5160
rect 11199 5120 11244 5148
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 13786 5120 14473 5148
rect 7466 5080 7472 5092
rect 7024 5052 7472 5080
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 7650 5080 7656 5092
rect 7611 5052 7656 5080
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 8662 5080 8668 5092
rect 8168 5052 8668 5080
rect 8168 5040 8174 5052
rect 8662 5040 8668 5052
rect 8720 5080 8726 5092
rect 8802 5083 8860 5089
rect 8802 5080 8814 5083
rect 8720 5052 8814 5080
rect 8720 5040 8726 5052
rect 8802 5049 8814 5052
rect 8848 5049 8860 5083
rect 12161 5083 12219 5089
rect 12161 5080 12173 5083
rect 8802 5043 8860 5049
rect 9416 5052 12173 5080
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 1452 4984 1593 5012
rect 1452 4972 1458 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 3694 5012 3700 5024
rect 3655 4984 3700 5012
rect 1581 4975 1639 4981
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4847 5015 4905 5021
rect 4847 4981 4859 5015
rect 4893 5012 4905 5015
rect 5074 5012 5080 5024
rect 4893 4984 5080 5012
rect 4893 4981 4905 4984
rect 4847 4975 4905 4981
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5500 4984 5549 5012
rect 5500 4972 5506 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 6638 5012 6644 5024
rect 6599 4984 6644 5012
rect 5537 4975 5595 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 9416 5021 9444 5052
rect 12161 5049 12173 5052
rect 12207 5080 12219 5083
rect 12342 5080 12348 5092
rect 12207 5052 12348 5080
rect 12207 5049 12219 5052
rect 12161 5043 12219 5049
rect 12342 5040 12348 5052
rect 12400 5040 12406 5092
rect 12526 5080 12532 5092
rect 12487 5052 12532 5080
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 12621 5083 12679 5089
rect 12621 5049 12633 5083
rect 12667 5049 12679 5083
rect 13170 5080 13176 5092
rect 13131 5052 13176 5080
rect 12621 5043 12679 5049
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 9272 4984 9413 5012
rect 9272 4972 9278 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 11882 5012 11888 5024
rect 11843 4984 11888 5012
rect 9401 4975 9459 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12360 5012 12388 5040
rect 12636 5012 12664 5043
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 12360 4984 12664 5012
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 13078 5012 13084 5024
rect 12768 4984 13084 5012
rect 12768 4972 12774 4984
rect 13078 4972 13084 4984
rect 13136 5012 13142 5024
rect 13786 5012 13814 5120
rect 14461 5117 14473 5120
rect 14507 5148 14519 5151
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14507 5120 14565 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 14734 5108 14740 5160
rect 14792 5148 14798 5160
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14792 5120 15025 5148
rect 14792 5108 14798 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 16301 5151 16359 5157
rect 16301 5117 16313 5151
rect 16347 5148 16359 5151
rect 16482 5148 16488 5160
rect 16347 5120 16488 5148
rect 16347 5117 16359 5120
rect 16301 5111 16359 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16853 5151 16911 5157
rect 16853 5148 16865 5151
rect 16632 5120 16865 5148
rect 16632 5108 16638 5120
rect 16853 5117 16865 5120
rect 16899 5117 16911 5151
rect 16853 5111 16911 5117
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 19610 5148 19616 5160
rect 19567 5120 19616 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 19610 5108 19616 5120
rect 19668 5108 19674 5160
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 20036 5120 20361 5148
rect 20036 5108 20042 5120
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20349 5111 20407 5117
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5148 20683 5151
rect 21542 5148 21548 5160
rect 20671 5120 21548 5148
rect 20671 5117 20683 5120
rect 20625 5111 20683 5117
rect 15289 5083 15347 5089
rect 15289 5049 15301 5083
rect 15335 5080 15347 5083
rect 15470 5080 15476 5092
rect 15335 5052 15476 5080
rect 15335 5049 15347 5052
rect 15289 5043 15347 5049
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 17126 5080 17132 5092
rect 17087 5052 17132 5080
rect 17126 5040 17132 5052
rect 17184 5040 17190 5092
rect 18969 5083 19027 5089
rect 18969 5049 18981 5083
rect 19015 5080 19027 5083
rect 19334 5080 19340 5092
rect 19015 5052 19340 5080
rect 19015 5049 19027 5052
rect 18969 5043 19027 5049
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 20257 5083 20315 5089
rect 20257 5049 20269 5083
rect 20303 5080 20315 5083
rect 20640 5080 20668 5111
rect 21542 5108 21548 5120
rect 21600 5108 21606 5160
rect 22002 5148 22008 5160
rect 21915 5120 22008 5148
rect 22002 5108 22008 5120
rect 22060 5108 22066 5160
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22278 5148 22284 5160
rect 22152 5120 22197 5148
rect 22239 5120 22284 5148
rect 22152 5108 22158 5120
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 23658 5148 23664 5160
rect 23619 5120 23664 5148
rect 23658 5108 23664 5120
rect 23716 5108 23722 5160
rect 23750 5108 23756 5160
rect 23808 5148 23814 5160
rect 23937 5151 23995 5157
rect 23808 5120 23853 5148
rect 23808 5108 23814 5120
rect 23937 5117 23949 5151
rect 23983 5148 23995 5151
rect 24026 5148 24032 5160
rect 23983 5120 24032 5148
rect 23983 5117 23995 5120
rect 23937 5111 23995 5117
rect 20303 5052 20668 5080
rect 22020 5080 22048 5108
rect 23474 5080 23480 5092
rect 22020 5052 22140 5080
rect 23387 5052 23480 5080
rect 20303 5049 20315 5052
rect 20257 5043 20315 5049
rect 13998 5012 14004 5024
rect 13136 4984 13814 5012
rect 13959 4984 14004 5012
rect 13136 4972 13142 4984
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 18506 5012 18512 5024
rect 18467 4984 18512 5012
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 20806 5012 20812 5024
rect 20767 4984 20812 5012
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 22112 5012 22140 5052
rect 23474 5040 23480 5052
rect 23532 5080 23538 5092
rect 23952 5080 23980 5111
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 23532 5052 23980 5080
rect 23532 5040 23538 5052
rect 24854 5040 24860 5092
rect 24912 5080 24918 5092
rect 25225 5083 25283 5089
rect 25225 5080 25237 5083
rect 24912 5052 25237 5080
rect 24912 5040 24918 5052
rect 25225 5049 25237 5052
rect 25271 5049 25283 5083
rect 25774 5080 25780 5092
rect 25735 5052 25780 5080
rect 25225 5043 25283 5049
rect 25774 5040 25780 5052
rect 25832 5040 25838 5092
rect 23658 5012 23664 5024
rect 22112 4984 23664 5012
rect 23658 4972 23664 4984
rect 23716 5012 23722 5024
rect 24670 5012 24676 5024
rect 23716 4984 24676 5012
rect 23716 4972 23722 4984
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 4571 4811 4629 4817
rect 4571 4777 4583 4811
rect 4617 4808 4629 4811
rect 7558 4808 7564 4820
rect 4617 4780 7564 4808
rect 4617 4777 4629 4780
rect 4571 4771 4629 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 7834 4808 7840 4820
rect 7795 4780 7840 4808
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8478 4808 8484 4820
rect 8343 4780 8484 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8478 4768 8484 4780
rect 8536 4808 8542 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8536 4780 9045 4808
rect 8536 4768 8542 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 9766 4768 9772 4820
rect 9824 4768 9830 4820
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 11238 4808 11244 4820
rect 10919 4780 11244 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 12526 4768 12532 4820
rect 12584 4808 12590 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12584 4780 12909 4808
rect 12584 4768 12590 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 12897 4771 12955 4777
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 14734 4808 14740 4820
rect 14691 4780 14740 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4808 15715 4811
rect 15746 4808 15752 4820
rect 15703 4780 15752 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16942 4808 16948 4820
rect 16903 4780 16948 4808
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 19518 4808 19524 4820
rect 19479 4780 19524 4808
rect 19518 4768 19524 4780
rect 19576 4768 19582 4820
rect 19978 4808 19984 4820
rect 19939 4780 19984 4808
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 20438 4808 20444 4820
rect 20399 4780 20444 4808
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22152 4780 24624 4808
rect 22152 4768 22158 4780
rect 9493 4743 9551 4749
rect 5368 4712 8616 4740
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 4500 4675 4558 4681
rect 4500 4672 4512 4675
rect 3660 4644 4512 4672
rect 3660 4632 3666 4644
rect 4500 4641 4512 4644
rect 4546 4672 4558 4675
rect 5368 4672 5396 4712
rect 4546 4644 5396 4672
rect 5445 4675 5503 4681
rect 4546 4641 4558 4644
rect 4500 4635 4558 4641
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 5534 4672 5540 4684
rect 5491 4644 5540 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6733 4675 6791 4681
rect 6733 4641 6745 4675
rect 6779 4672 6791 4675
rect 6822 4672 6828 4684
rect 6779 4644 6828 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6972 4644 7021 4672
rect 6972 4632 6978 4644
rect 7009 4641 7021 4644
rect 7055 4672 7067 4675
rect 7098 4672 7104 4684
rect 7055 4644 7104 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7466 4672 7472 4684
rect 7427 4644 7472 4672
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 8202 4672 8208 4684
rect 8163 4644 8208 4672
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8481 4675 8539 4681
rect 8481 4672 8493 4675
rect 8352 4644 8493 4672
rect 8352 4632 8358 4644
rect 8481 4641 8493 4644
rect 8527 4641 8539 4675
rect 8481 4635 8539 4641
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4604 7251 4607
rect 8386 4604 8392 4616
rect 7239 4576 8392 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 5583 4539 5641 4545
rect 5583 4505 5595 4539
rect 5629 4536 5641 4539
rect 7558 4536 7564 4548
rect 5629 4508 7564 4536
rect 5629 4505 5641 4508
rect 5583 4499 5641 4505
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 8588 4536 8616 4712
rect 9493 4709 9505 4743
rect 9539 4740 9551 4743
rect 9784 4740 9812 4768
rect 9953 4743 10011 4749
rect 9953 4740 9965 4743
rect 9539 4712 9965 4740
rect 9539 4709 9551 4712
rect 9493 4703 9551 4709
rect 9953 4709 9965 4712
rect 9999 4709 10011 4743
rect 9953 4703 10011 4709
rect 11695 4743 11753 4749
rect 11695 4709 11707 4743
rect 11741 4740 11753 4743
rect 12250 4740 12256 4752
rect 11741 4712 12256 4740
rect 11741 4709 11753 4712
rect 11695 4703 11753 4709
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 13262 4740 13268 4752
rect 13223 4712 13268 4740
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 18506 4740 18512 4752
rect 18467 4712 18512 4740
rect 18506 4700 18512 4712
rect 18564 4700 18570 4752
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 11514 4672 11520 4684
rect 10551 4644 11520 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9306 4604 9312 4616
rect 9180 4576 9312 4604
rect 9180 4564 9186 4576
rect 9306 4564 9312 4576
rect 9364 4604 9370 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9364 4576 9873 4604
rect 9364 4564 9370 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10520 4536 10548 4635
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 16758 4632 16764 4684
rect 16816 4672 16822 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16816 4644 17049 4672
rect 16816 4632 16822 4644
rect 17037 4641 17049 4644
rect 17083 4641 17095 4675
rect 19150 4672 19156 4684
rect 19063 4644 19156 4672
rect 17037 4635 17095 4641
rect 19150 4632 19156 4644
rect 19208 4672 19214 4684
rect 19536 4672 19564 4768
rect 24118 4740 24124 4752
rect 23952 4712 24124 4740
rect 19208 4644 19564 4672
rect 19208 4632 19214 4644
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20864 4644 20913 4672
rect 20864 4632 20870 4644
rect 20901 4641 20913 4644
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 22554 4632 22560 4684
rect 22612 4672 22618 4684
rect 23017 4675 23075 4681
rect 23017 4672 23029 4675
rect 22612 4644 23029 4672
rect 22612 4632 22618 4644
rect 23017 4641 23029 4644
rect 23063 4672 23075 4675
rect 23474 4672 23480 4684
rect 23063 4644 23480 4672
rect 23063 4641 23075 4644
rect 23017 4635 23075 4641
rect 23474 4632 23480 4644
rect 23532 4632 23538 4684
rect 23750 4672 23756 4684
rect 23663 4644 23756 4672
rect 23750 4632 23756 4644
rect 23808 4672 23814 4684
rect 23952 4681 23980 4712
rect 24118 4700 24124 4712
rect 24176 4700 24182 4752
rect 24596 4681 24624 4780
rect 23937 4675 23995 4681
rect 23937 4672 23949 4675
rect 23808 4644 23949 4672
rect 23808 4632 23814 4644
rect 23937 4641 23949 4644
rect 23983 4641 23995 4675
rect 23937 4635 23995 4641
rect 24581 4675 24639 4681
rect 24581 4641 24593 4675
rect 24627 4672 24639 4675
rect 24946 4672 24952 4684
rect 24627 4644 24952 4672
rect 24627 4641 24639 4644
rect 24581 4635 24639 4641
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11296 4576 11345 4604
rect 11296 4564 11302 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 11333 4567 11391 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13173 4567 13231 4573
rect 8588 4508 10548 4536
rect 10870 4496 10876 4548
rect 10928 4536 10934 4548
rect 11149 4539 11207 4545
rect 11149 4536 11161 4539
rect 10928 4508 11161 4536
rect 10928 4496 10934 4508
rect 11149 4505 11161 4508
rect 11195 4536 11207 4539
rect 13078 4536 13084 4548
rect 11195 4508 13084 4536
rect 11195 4505 11207 4508
rect 11149 4499 11207 4505
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 13188 4536 13216 4567
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 15470 4604 15476 4616
rect 15335 4576 15476 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4604 22155 4607
rect 22278 4604 22284 4616
rect 22143 4576 22284 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 22278 4564 22284 4576
rect 22336 4604 22342 4616
rect 23109 4607 23167 4613
rect 23109 4604 23121 4607
rect 22336 4576 23121 4604
rect 22336 4564 22342 4576
rect 23109 4573 23121 4576
rect 23155 4604 23167 4607
rect 24210 4604 24216 4616
rect 23155 4576 24216 4604
rect 23155 4573 23167 4576
rect 23109 4567 23167 4573
rect 24210 4564 24216 4576
rect 24268 4564 24274 4616
rect 13446 4536 13452 4548
rect 13188 4508 13452 4536
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 18138 4536 18144 4548
rect 18051 4508 18144 4536
rect 18138 4496 18144 4508
rect 18196 4536 18202 4548
rect 22738 4536 22744 4548
rect 18196 4508 22744 4536
rect 18196 4496 18202 4508
rect 22738 4496 22744 4508
rect 22796 4496 22802 4548
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9122 4468 9128 4480
rect 8260 4440 9128 4468
rect 8260 4428 8266 4440
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 11388 4440 12265 4468
rect 11388 4428 11394 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 16206 4468 16212 4480
rect 16167 4440 16212 4468
rect 12253 4431 12311 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16574 4468 16580 4480
rect 16535 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 17221 4471 17279 4477
rect 17221 4437 17233 4471
rect 17267 4468 17279 4471
rect 17954 4468 17960 4480
rect 17267 4440 17960 4468
rect 17267 4437 17279 4440
rect 17221 4431 17279 4437
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 18230 4428 18236 4480
rect 18288 4468 18294 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 18288 4440 21097 4468
rect 18288 4428 18294 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21542 4468 21548 4480
rect 21503 4440 21548 4468
rect 21085 4431 21143 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 3602 4264 3608 4276
rect 3563 4236 3608 4264
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 3970 4264 3976 4276
rect 3931 4236 3976 4264
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 5534 4264 5540 4276
rect 5447 4236 5540 4264
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 8938 4264 8944 4276
rect 5592 4236 8944 4264
rect 5592 4224 5598 4236
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9180 4236 9781 4264
rect 9180 4224 9186 4236
rect 9769 4233 9781 4236
rect 9815 4264 9827 4267
rect 10962 4264 10968 4276
rect 9815 4236 10968 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 11756 4236 11897 4264
rect 11756 4224 11762 4236
rect 11885 4233 11897 4236
rect 11931 4264 11943 4267
rect 12250 4264 12256 4276
rect 11931 4236 12256 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12250 4224 12256 4236
rect 12308 4264 12314 4276
rect 16206 4264 16212 4276
rect 12308 4236 14412 4264
rect 16167 4236 16212 4264
rect 12308 4224 12314 4236
rect 4617 4199 4675 4205
rect 4617 4165 4629 4199
rect 4663 4196 4675 4199
rect 5350 4196 5356 4208
rect 4663 4168 5356 4196
rect 4663 4165 4675 4168
rect 4617 4159 4675 4165
rect 4759 4069 4787 4168
rect 5350 4156 5356 4168
rect 5408 4156 5414 4208
rect 5859 4199 5917 4205
rect 5859 4165 5871 4199
rect 5905 4196 5917 4199
rect 5994 4196 6000 4208
rect 5905 4168 6000 4196
rect 5905 4165 5917 4168
rect 5859 4159 5917 4165
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 8389 4199 8447 4205
rect 6880 4168 7512 4196
rect 6880 4156 6886 4168
rect 3764 4063 3822 4069
rect 3764 4029 3776 4063
rect 3810 4060 3822 4063
rect 4744 4063 4802 4069
rect 3810 4032 4154 4060
rect 3810 4029 3822 4032
rect 3764 4023 3822 4029
rect 4126 3924 4154 4032
rect 4744 4029 4756 4063
rect 4790 4029 4802 4063
rect 4744 4023 4802 4029
rect 5788 4063 5846 4069
rect 5788 4029 5800 4063
rect 5834 4060 5846 4063
rect 6917 4063 6975 4069
rect 5834 4032 6316 4060
rect 5834 4029 5846 4032
rect 5788 4023 5846 4029
rect 4246 3924 4252 3936
rect 4126 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4847 3927 4905 3933
rect 4847 3893 4859 3927
rect 4893 3924 4905 3927
rect 5166 3924 5172 3936
rect 4893 3896 5172 3924
rect 4893 3893 4905 3896
rect 4847 3887 4905 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6288 3933 6316 4032
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 6932 3992 6960 4023
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7064 4032 7389 4060
rect 7064 4020 7070 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7484 4060 7512 4168
rect 8389 4165 8401 4199
rect 8435 4196 8447 4199
rect 8662 4196 8668 4208
rect 8435 4168 8668 4196
rect 8435 4165 8447 4168
rect 8389 4159 8447 4165
rect 8662 4156 8668 4168
rect 8720 4196 8726 4208
rect 10042 4196 10048 4208
rect 8720 4168 10048 4196
rect 8720 4156 8726 4168
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 14093 4199 14151 4205
rect 14093 4165 14105 4199
rect 14139 4196 14151 4199
rect 14182 4196 14188 4208
rect 14139 4168 14188 4196
rect 14139 4165 14151 4168
rect 14093 4159 14151 4165
rect 14182 4156 14188 4168
rect 14240 4156 14246 4208
rect 14384 4205 14412 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 19150 4264 19156 4276
rect 19111 4236 19156 4264
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 21174 4224 21180 4276
rect 21232 4264 21238 4276
rect 21269 4267 21327 4273
rect 21269 4264 21281 4267
rect 21232 4236 21281 4264
rect 21232 4224 21238 4236
rect 21269 4233 21281 4236
rect 21315 4233 21327 4267
rect 22833 4267 22891 4273
rect 22833 4264 22845 4267
rect 21269 4227 21327 4233
rect 21560 4236 22845 4264
rect 14369 4199 14427 4205
rect 14369 4196 14381 4199
rect 14279 4168 14381 4196
rect 14369 4165 14381 4168
rect 14415 4165 14427 4199
rect 14369 4159 14427 4165
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 9122 4128 9128 4140
rect 7699 4100 9128 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 11238 4128 11244 4140
rect 10704 4100 11244 4128
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7484 4032 7941 4060
rect 7377 4023 7435 4029
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8444 4032 8493 4060
rect 8444 4020 8450 4032
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 8527 4032 10057 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 7098 3992 7104 4004
rect 6687 3964 7104 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 8662 3992 8668 4004
rect 8575 3964 8668 3992
rect 8662 3952 8668 3964
rect 8720 3992 8726 4004
rect 8802 3995 8860 4001
rect 8802 3992 8814 3995
rect 8720 3964 8814 3992
rect 8720 3952 8726 3964
rect 8802 3961 8814 3964
rect 8848 3961 8860 3995
rect 10704 3992 10732 4100
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 10870 3992 10876 4004
rect 8802 3955 8860 3961
rect 9226 3964 10732 3992
rect 10831 3964 10876 3992
rect 6273 3927 6331 3933
rect 6273 3893 6285 3927
rect 6319 3924 6331 3927
rect 6822 3924 6828 3936
rect 6319 3896 6828 3924
rect 6319 3893 6331 3896
rect 6273 3887 6331 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 9226 3924 9254 3964
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3992 11023 3995
rect 11330 3992 11336 4004
rect 11011 3964 11336 3992
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 9398 3924 9404 3936
rect 7708 3896 9254 3924
rect 9359 3896 9404 3924
rect 7708 3884 7714 3896
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 10689 3927 10747 3933
rect 10689 3893 10701 3927
rect 10735 3924 10747 3927
rect 10980 3924 11008 3955
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 11514 3992 11520 4004
rect 11475 3964 11520 3992
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 12526 3992 12532 4004
rect 12487 3964 12532 3992
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3992 12679 3995
rect 13262 3992 13268 4004
rect 12667 3964 13268 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 12158 3924 12164 3936
rect 10735 3896 11008 3924
rect 12119 3896 12164 3924
rect 10735 3893 10747 3896
rect 10689 3887 10747 3893
rect 12158 3884 12164 3896
rect 12216 3924 12222 3936
rect 12636 3924 12664 3955
rect 13262 3952 13268 3964
rect 13320 3992 13326 4004
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 13320 3964 13461 3992
rect 13320 3952 13326 3964
rect 13449 3961 13461 3964
rect 13495 3961 13507 3995
rect 14384 3992 14412 4159
rect 14458 4156 14464 4208
rect 14516 4196 14522 4208
rect 16574 4196 16580 4208
rect 14516 4168 14596 4196
rect 14516 4156 14522 4168
rect 14568 4137 14596 4168
rect 16408 4168 16580 4196
rect 16408 4137 16436 4168
rect 16574 4156 16580 4168
rect 16632 4196 16638 4208
rect 19797 4199 19855 4205
rect 16632 4168 18276 4196
rect 16632 4156 16638 4168
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4097 14611 4131
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 16371 4100 16405 4128
rect 14553 4091 14611 4097
rect 16393 4097 16405 4100
rect 16439 4097 16451 4131
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 16393 4091 16451 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 16816 4100 17325 4128
rect 16816 4088 16822 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 18138 4128 18144 4140
rect 18099 4100 18144 4128
rect 17313 4091 17371 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18248 4128 18276 4168
rect 19797 4165 19809 4199
rect 19843 4196 19855 4199
rect 19981 4199 20039 4205
rect 19981 4196 19993 4199
rect 19843 4168 19993 4196
rect 19843 4165 19855 4168
rect 19797 4159 19855 4165
rect 19981 4165 19993 4168
rect 20027 4196 20039 4199
rect 20438 4196 20444 4208
rect 20027 4168 20444 4196
rect 20027 4165 20039 4168
rect 19981 4159 20039 4165
rect 20438 4156 20444 4168
rect 20496 4156 20502 4208
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 18248 4100 18429 4128
rect 18417 4097 18429 4100
rect 18463 4097 18475 4131
rect 18417 4091 18475 4097
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4060 19947 4063
rect 20070 4060 20076 4072
rect 19935 4032 20076 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20254 4060 20260 4072
rect 20211 4032 20260 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 21284 4060 21312 4227
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 21560 4205 21588 4236
rect 22833 4233 22845 4236
rect 22879 4264 22891 4267
rect 25406 4264 25412 4276
rect 22879 4236 23474 4264
rect 25367 4236 25412 4264
rect 22879 4233 22891 4236
rect 22833 4227 22891 4233
rect 21545 4199 21603 4205
rect 21545 4196 21557 4199
rect 21508 4168 21557 4196
rect 21508 4156 21514 4168
rect 21545 4165 21557 4168
rect 21591 4165 21603 4199
rect 22554 4196 22560 4208
rect 22515 4168 22560 4196
rect 21545 4159 21603 4165
rect 22554 4156 22560 4168
rect 22612 4156 22618 4208
rect 23446 4196 23474 4236
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 23658 4196 23664 4208
rect 23446 4168 23664 4196
rect 23658 4156 23664 4168
rect 23716 4196 23722 4208
rect 23753 4199 23811 4205
rect 23753 4196 23765 4199
rect 23716 4168 23765 4196
rect 23716 4156 23722 4168
rect 23753 4165 23765 4168
rect 23799 4165 23811 4199
rect 23753 4159 23811 4165
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4128 22247 4131
rect 22922 4128 22928 4140
rect 22235 4100 22928 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22922 4088 22928 4100
rect 22980 4088 22986 4140
rect 25041 4131 25099 4137
rect 25041 4128 25053 4131
rect 23676 4100 25053 4128
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 21284 4032 21465 4060
rect 21453 4029 21465 4032
rect 21499 4029 21511 4063
rect 21726 4060 21732 4072
rect 21687 4032 21732 4060
rect 21453 4023 21511 4029
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 21818 4020 21824 4072
rect 21876 4060 21882 4072
rect 23676 4069 23704 4100
rect 25041 4097 25053 4100
rect 25087 4097 25099 4131
rect 25041 4091 25099 4097
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 21876 4032 23673 4060
rect 21876 4020 21882 4032
rect 23661 4029 23673 4032
rect 23707 4029 23719 4063
rect 23661 4023 23719 4029
rect 23937 4063 23995 4069
rect 23937 4029 23949 4063
rect 23983 4029 23995 4063
rect 23937 4023 23995 4029
rect 24397 4063 24455 4069
rect 24397 4029 24409 4063
rect 24443 4060 24455 4063
rect 25225 4063 25283 4069
rect 25225 4060 25237 4063
rect 24443 4032 25237 4060
rect 24443 4029 24455 4032
rect 24397 4023 24455 4029
rect 25225 4029 25237 4032
rect 25271 4060 25283 4063
rect 25685 4063 25743 4069
rect 25685 4060 25697 4063
rect 25271 4032 25697 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25685 4029 25697 4032
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 14915 3995 14973 4001
rect 14915 3992 14927 3995
rect 14384 3964 14927 3992
rect 13449 3955 13507 3961
rect 14915 3961 14927 3964
rect 14961 3992 14973 3995
rect 14961 3964 15792 3992
rect 14961 3961 14973 3964
rect 14915 3955 14973 3961
rect 15764 3936 15792 3964
rect 16206 3952 16212 4004
rect 16264 3992 16270 4004
rect 16485 3995 16543 4001
rect 16485 3992 16497 3995
rect 16264 3964 16497 3992
rect 16264 3952 16270 3964
rect 16485 3961 16497 3964
rect 16531 3961 16543 3995
rect 17678 3992 17684 4004
rect 16485 3955 16543 3961
rect 17144 3964 17684 3992
rect 12216 3896 12664 3924
rect 12216 3884 12222 3896
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 15473 3927 15531 3933
rect 15473 3924 15485 3927
rect 13872 3896 15485 3924
rect 13872 3884 13878 3896
rect 15473 3893 15485 3896
rect 15519 3893 15531 3927
rect 15473 3887 15531 3893
rect 15746 3884 15752 3936
rect 15804 3924 15810 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15804 3896 15853 3924
rect 15804 3884 15810 3896
rect 15841 3893 15853 3896
rect 15887 3924 15899 3927
rect 17144 3924 17172 3964
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 17865 3995 17923 4001
rect 17865 3961 17877 3995
rect 17911 3992 17923 3995
rect 18233 3995 18291 4001
rect 18233 3992 18245 3995
rect 17911 3964 18245 3992
rect 17911 3961 17923 3964
rect 17865 3955 17923 3961
rect 18233 3961 18245 3964
rect 18279 3992 18291 3995
rect 18506 3992 18512 4004
rect 18279 3964 18512 3992
rect 18279 3961 18291 3964
rect 18233 3955 18291 3961
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 20625 3995 20683 4001
rect 20625 3961 20637 3995
rect 20671 3992 20683 3995
rect 22738 3992 22744 4004
rect 20671 3964 22744 3992
rect 20671 3961 20683 3964
rect 20625 3955 20683 3961
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 15887 3896 17172 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 20070 3884 20076 3936
rect 20128 3924 20134 3936
rect 21818 3924 21824 3936
rect 20128 3896 21824 3924
rect 20128 3884 20134 3896
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 23014 3884 23020 3936
rect 23072 3924 23078 3936
rect 23385 3927 23443 3933
rect 23385 3924 23397 3927
rect 23072 3896 23397 3924
rect 23072 3884 23078 3896
rect 23385 3893 23397 3896
rect 23431 3924 23443 3927
rect 23952 3924 23980 4023
rect 23431 3896 23980 3924
rect 24765 3927 24823 3933
rect 23431 3893 23443 3896
rect 23385 3887 23443 3893
rect 24765 3893 24777 3927
rect 24811 3924 24823 3927
rect 24946 3924 24952 3936
rect 24811 3896 24952 3924
rect 24811 3893 24823 3896
rect 24765 3887 24823 3893
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 7064 3692 7481 3720
rect 7064 3680 7070 3692
rect 7469 3689 7481 3692
rect 7515 3720 7527 3723
rect 7834 3720 7840 3732
rect 7515 3692 7840 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 9824 3692 10609 3720
rect 9824 3680 9830 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 10597 3683 10655 3689
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 11296 3692 11345 3720
rect 11296 3680 11302 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 13596 3692 15025 3720
rect 13596 3680 13602 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15470 3720 15476 3732
rect 15431 3692 15476 3720
rect 15013 3683 15071 3689
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 16666 3720 16672 3732
rect 15764 3692 16672 3720
rect 6365 3655 6423 3661
rect 6365 3621 6377 3655
rect 6411 3652 6423 3655
rect 7024 3652 7052 3680
rect 6411 3624 7052 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 2866 3584 2872 3596
rect 2827 3556 2872 3584
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 4500 3587 4558 3593
rect 4500 3553 4512 3587
rect 4546 3584 4558 3587
rect 4614 3584 4620 3596
rect 4546 3556 4620 3584
rect 4546 3553 4558 3556
rect 4500 3547 4558 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5480 3587 5538 3593
rect 5480 3584 5492 3587
rect 5408 3556 5492 3584
rect 5408 3544 5414 3556
rect 5480 3553 5492 3556
rect 5526 3553 5538 3587
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 5480 3547 5538 3553
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 7024 3593 7052 3624
rect 8205 3655 8263 3661
rect 8205 3621 8217 3655
rect 8251 3652 8263 3655
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8251 3624 9045 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 9033 3621 9045 3624
rect 9079 3652 9091 3655
rect 9398 3652 9404 3664
rect 9079 3624 9404 3652
rect 9079 3621 9091 3624
rect 9033 3615 9091 3621
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 9930 3655 9988 3661
rect 9930 3621 9942 3655
rect 9976 3652 9988 3655
rect 10042 3652 10048 3664
rect 9976 3624 10048 3652
rect 9976 3621 9988 3624
rect 9930 3615 9988 3621
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 12206 3655 12264 3661
rect 12206 3652 12218 3655
rect 11756 3624 12218 3652
rect 11756 3612 11762 3624
rect 12206 3621 12218 3624
rect 12252 3621 12264 3655
rect 12206 3615 12264 3621
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 13814 3652 13820 3664
rect 13780 3624 13820 3652
rect 13780 3612 13786 3624
rect 13814 3612 13820 3624
rect 13872 3652 13878 3664
rect 13872 3624 13917 3652
rect 13872 3612 13878 3624
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 9180 3556 11897 3584
rect 9180 3544 9186 3556
rect 11885 3553 11897 3556
rect 11931 3584 11943 3587
rect 11974 3584 11980 3596
rect 11931 3556 11980 3584
rect 11931 3553 11943 3556
rect 11885 3547 11943 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 5583 3519 5641 3525
rect 5583 3485 5595 3519
rect 5629 3516 5641 3519
rect 6914 3516 6920 3528
rect 5629 3488 6920 3516
rect 5629 3485 5641 3488
rect 5583 3479 5641 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7190 3516 7196 3528
rect 7151 3488 7196 3516
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 8754 3516 8760 3528
rect 8715 3488 8760 3516
rect 8113 3479 8171 3485
rect 5994 3448 6000 3460
rect 4126 3420 6000 3448
rect 3099 3383 3157 3389
rect 3099 3349 3111 3383
rect 3145 3380 3157 3383
rect 4126 3380 4154 3420
rect 5994 3408 6000 3420
rect 6052 3448 6058 3460
rect 8128 3448 8156 3479
rect 8754 3476 8760 3488
rect 8812 3516 8818 3528
rect 9306 3516 9312 3528
rect 8812 3488 9312 3516
rect 8812 3476 8818 3488
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9674 3516 9680 3528
rect 9635 3488 9680 3516
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 13906 3516 13912 3528
rect 13771 3488 13912 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 14090 3476 14096 3488
rect 14148 3516 14154 3528
rect 15764 3516 15792 3692
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 17126 3680 17132 3732
rect 17184 3720 17190 3732
rect 17405 3723 17463 3729
rect 17405 3720 17417 3723
rect 17184 3692 17417 3720
rect 17184 3680 17190 3692
rect 17405 3689 17417 3692
rect 17451 3720 17463 3723
rect 18506 3720 18512 3732
rect 17451 3692 17632 3720
rect 18467 3692 18512 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15988 3624 16037 3652
rect 15988 3612 15994 3624
rect 16025 3621 16037 3624
rect 16071 3652 16083 3655
rect 16390 3652 16396 3664
rect 16071 3624 16396 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 16574 3652 16580 3664
rect 16535 3624 16580 3652
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 17604 3593 17632 3692
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 23658 3720 23664 3732
rect 23619 3692 23664 3720
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 24670 3720 24676 3732
rect 24044 3692 24676 3720
rect 17678 3612 17684 3664
rect 17736 3652 17742 3664
rect 17910 3655 17968 3661
rect 17910 3652 17922 3655
rect 17736 3624 17922 3652
rect 17736 3612 17742 3624
rect 17910 3621 17922 3624
rect 17956 3621 17968 3655
rect 17910 3615 17968 3621
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3553 17647 3587
rect 17589 3547 17647 3553
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19334 3584 19340 3596
rect 18380 3556 19340 3584
rect 18380 3544 18386 3556
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 21545 3587 21603 3593
rect 21545 3553 21557 3587
rect 21591 3584 21603 3587
rect 21726 3584 21732 3596
rect 21591 3556 21732 3584
rect 21591 3553 21603 3556
rect 21545 3547 21603 3553
rect 21726 3544 21732 3556
rect 21784 3544 21790 3596
rect 22278 3544 22284 3596
rect 22336 3584 22342 3596
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22336 3556 22477 3584
rect 22336 3544 22342 3556
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 23014 3584 23020 3596
rect 22787 3556 23020 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 23014 3544 23020 3556
rect 23072 3544 23078 3596
rect 24044 3593 24072 3692
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 24268 3624 24348 3652
rect 24268 3612 24274 3624
rect 24029 3587 24087 3593
rect 24029 3553 24041 3587
rect 24075 3553 24087 3587
rect 24029 3547 24087 3553
rect 24118 3544 24124 3596
rect 24176 3584 24182 3596
rect 24320 3593 24348 3624
rect 24305 3587 24363 3593
rect 24176 3556 24221 3584
rect 24176 3544 24182 3556
rect 24305 3553 24317 3587
rect 24351 3553 24363 3587
rect 24305 3547 24363 3553
rect 14148 3488 15792 3516
rect 15933 3519 15991 3525
rect 14148 3476 14154 3488
rect 15933 3485 15945 3519
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 11701 3451 11759 3457
rect 11701 3448 11713 3451
rect 6052 3420 8156 3448
rect 8817 3420 11713 3448
rect 6052 3408 6058 3420
rect 3145 3352 4154 3380
rect 4571 3383 4629 3389
rect 3145 3349 3157 3352
rect 3099 3343 3157 3349
rect 4571 3349 4583 3383
rect 4617 3380 4629 3383
rect 5442 3380 5448 3392
rect 4617 3352 5448 3380
rect 4617 3349 4629 3352
rect 4571 3343 4629 3349
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 6086 3380 6092 3392
rect 5951 3352 6092 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 8817 3380 8845 3420
rect 11701 3417 11713 3420
rect 11747 3448 11759 3451
rect 12526 3448 12532 3460
rect 11747 3420 12532 3448
rect 11747 3417 11759 3420
rect 11701 3411 11759 3417
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 13446 3448 13452 3460
rect 13407 3420 13452 3448
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 15948 3448 15976 3479
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 22925 3519 22983 3525
rect 22925 3516 22937 3519
rect 20220 3488 22937 3516
rect 20220 3476 20226 3488
rect 22925 3485 22937 3488
rect 22971 3485 22983 3519
rect 22925 3479 22983 3485
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 24489 3519 24547 3525
rect 24489 3516 24501 3519
rect 23164 3488 24501 3516
rect 23164 3476 23170 3488
rect 24489 3485 24501 3488
rect 24535 3485 24547 3519
rect 24489 3479 24547 3485
rect 16482 3448 16488 3460
rect 15948 3420 16488 3448
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17310 3408 17316 3460
rect 17368 3448 17374 3460
rect 19521 3451 19579 3457
rect 19521 3448 19533 3451
rect 17368 3420 19533 3448
rect 17368 3408 17374 3420
rect 19521 3417 19533 3420
rect 19567 3417 19579 3451
rect 22554 3448 22560 3460
rect 22515 3420 22560 3448
rect 19521 3411 19579 3417
rect 22554 3408 22560 3420
rect 22612 3408 22618 3460
rect 9398 3380 9404 3392
rect 6236 3352 8845 3380
rect 9359 3352 9404 3380
rect 6236 3340 6242 3352
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 10686 3340 10692 3392
rect 10744 3380 10750 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10744 3352 10885 3380
rect 10744 3340 10750 3352
rect 10873 3349 10885 3352
rect 10919 3349 10931 3383
rect 10873 3343 10931 3349
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 12805 3383 12863 3389
rect 12805 3380 12817 3383
rect 12676 3352 12817 3380
rect 12676 3340 12682 3352
rect 12805 3349 12817 3352
rect 12851 3380 12863 3383
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 12851 3352 13093 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 13081 3349 13093 3352
rect 13127 3349 13139 3383
rect 13081 3343 13139 3349
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 14608 3352 14657 3380
rect 14608 3340 14614 3352
rect 14645 3349 14657 3352
rect 14691 3349 14703 3383
rect 18874 3380 18880 3392
rect 18835 3352 18880 3380
rect 14645 3343 14703 3349
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3380 20039 3383
rect 20254 3380 20260 3392
rect 20027 3352 20260 3380
rect 20027 3349 20039 3352
rect 19981 3343 20039 3349
rect 20254 3340 20260 3352
rect 20312 3380 20318 3392
rect 21358 3380 21364 3392
rect 20312 3352 21364 3380
rect 20312 3340 20318 3352
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 22186 3380 22192 3392
rect 22147 3352 22192 3380
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 4614 3176 4620 3188
rect 3292 3148 4154 3176
rect 4575 3148 4620 3176
rect 3292 3136 3298 3148
rect 4126 3108 4154 3148
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6454 3176 6460 3188
rect 6415 3148 6460 3176
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8662 3176 8668 3188
rect 8623 3148 8668 3176
rect 8662 3136 8668 3148
rect 8720 3176 8726 3188
rect 10042 3176 10048 3188
rect 8720 3148 10048 3176
rect 8720 3136 8726 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11756 3148 11897 3176
rect 11756 3136 11762 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 13722 3176 13728 3188
rect 13683 3148 13728 3176
rect 11885 3139 11943 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 15562 3176 15568 3188
rect 15523 3148 15568 3176
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 15930 3176 15936 3188
rect 15891 3148 15936 3176
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 17678 3176 17684 3188
rect 17639 3148 17684 3176
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 19334 3176 19340 3188
rect 19295 3148 19340 3176
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 20162 3176 20168 3188
rect 20123 3148 20168 3176
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 21726 3176 21732 3188
rect 21639 3148 21732 3176
rect 21726 3136 21732 3148
rect 21784 3176 21790 3188
rect 23014 3176 23020 3188
rect 21784 3148 23020 3176
rect 21784 3136 21790 3148
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 24118 3136 24124 3188
rect 24176 3176 24182 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 24176 3148 24409 3176
rect 24176 3136 24182 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24397 3139 24455 3145
rect 4126 3080 9536 3108
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2924 3012 3065 3040
rect 2924 3000 2930 3012
rect 3053 3009 3065 3012
rect 3099 3040 3111 3043
rect 4890 3040 4896 3052
rect 3099 3012 4896 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5408 3012 5641 3040
rect 5408 3000 5414 3012
rect 5629 3009 5641 3012
rect 5675 3040 5687 3043
rect 6270 3040 6276 3052
rect 5675 3012 6276 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 7248 3012 8861 3040
rect 7248 3000 7254 3012
rect 8849 3009 8861 3012
rect 8895 3040 8907 3043
rect 9398 3040 9404 3052
rect 8895 3012 9404 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2972 2375 2975
rect 2406 2972 2412 2984
rect 2464 2981 2470 2984
rect 2464 2975 2502 2981
rect 2363 2944 2412 2972
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 2406 2932 2412 2944
rect 2490 2941 2502 2975
rect 2464 2935 2502 2941
rect 3764 2975 3822 2981
rect 3764 2941 3776 2975
rect 3810 2972 3822 2975
rect 4776 2975 4834 2981
rect 3810 2944 4154 2972
rect 3810 2941 3822 2944
rect 3764 2935 3822 2941
rect 2464 2932 2470 2935
rect 4126 2848 4154 2944
rect 4776 2941 4788 2975
rect 4822 2972 4834 2975
rect 5258 2972 5264 2984
rect 4822 2944 5264 2972
rect 4822 2941 4834 2944
rect 4776 2935 4834 2941
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 5788 2975 5846 2981
rect 5788 2941 5800 2975
rect 5834 2972 5846 2975
rect 6086 2972 6092 2984
rect 5834 2944 6092 2972
rect 5834 2941 5846 2944
rect 5788 2935 5846 2941
rect 6086 2932 6092 2944
rect 6144 2972 6150 2984
rect 6362 2972 6368 2984
rect 6144 2944 6368 2972
rect 6144 2932 6150 2944
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 7282 2932 7288 2984
rect 7340 2972 7346 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7340 2944 7573 2972
rect 7340 2932 7346 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7834 2972 7840 2984
rect 7795 2944 7840 2972
rect 7561 2935 7619 2941
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 7374 2904 7380 2916
rect 5132 2876 7380 2904
rect 5132 2864 5138 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7576 2904 7604 2935
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8067 2944 9352 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 7576 2876 8432 2904
rect 8404 2848 8432 2876
rect 8662 2864 8668 2916
rect 8720 2904 8726 2916
rect 9170 2907 9228 2913
rect 9170 2904 9182 2907
rect 8720 2876 9182 2904
rect 8720 2864 8726 2876
rect 9170 2873 9182 2876
rect 9216 2873 9228 2907
rect 9170 2867 9228 2873
rect 2547 2839 2605 2845
rect 2547 2805 2559 2839
rect 2593 2836 2605 2839
rect 3694 2836 3700 2848
rect 2593 2808 3700 2836
rect 2593 2805 2605 2808
rect 2547 2799 2605 2805
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 3835 2839 3893 2845
rect 3835 2805 3847 2839
rect 3881 2836 3893 2839
rect 3970 2836 3976 2848
rect 3881 2808 3976 2836
rect 3881 2805 3893 2808
rect 3835 2799 3893 2805
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 4126 2808 4160 2848
rect 4154 2796 4160 2808
rect 4212 2836 4218 2848
rect 4847 2839 4905 2845
rect 4212 2808 4257 2836
rect 4212 2796 4218 2808
rect 4847 2805 4859 2839
rect 4893 2836 4905 2839
rect 4982 2836 4988 2848
rect 4893 2808 4988 2836
rect 4893 2805 4905 2808
rect 4847 2799 4905 2805
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5859 2839 5917 2845
rect 5859 2805 5871 2839
rect 5905 2836 5917 2839
rect 6638 2836 6644 2848
rect 5905 2808 6644 2836
rect 5905 2805 5917 2808
rect 5859 2799 5917 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 8386 2836 8392 2848
rect 8347 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 9324 2836 9352 2944
rect 9508 2904 9536 3080
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 19797 3111 19855 3117
rect 19797 3108 19809 3111
rect 18656 3080 19809 3108
rect 18656 3068 18662 3080
rect 19797 3077 19809 3080
rect 19843 3077 19855 3111
rect 22370 3108 22376 3120
rect 22331 3080 22376 3108
rect 19797 3071 19855 3077
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 23842 3068 23848 3120
rect 23900 3108 23906 3120
rect 24765 3111 24823 3117
rect 24765 3108 24777 3111
rect 23900 3080 24777 3108
rect 23900 3068 23906 3080
rect 24765 3077 24777 3080
rect 24811 3077 24823 3111
rect 24765 3071 24823 3077
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 10928 3012 11161 3040
rect 10928 3000 10934 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11514 3000 11520 3052
rect 11572 3040 11578 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 11572 3012 12817 3040
rect 11572 3000 11578 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 16574 3040 16580 3052
rect 16535 3012 16580 3040
rect 12805 3003 12863 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18874 3040 18880 3052
rect 18187 3012 18880 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3040 21419 3043
rect 21818 3040 21824 3052
rect 21407 3012 21824 3040
rect 21407 3009 21419 3012
rect 21361 3003 21419 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22094 3040 22100 3052
rect 22007 3012 22100 3040
rect 22094 3000 22100 3012
rect 22152 3040 22158 3052
rect 22554 3040 22560 3052
rect 22152 3012 22560 3040
rect 22152 3000 22158 3012
rect 22554 3000 22560 3012
rect 22612 3040 22618 3052
rect 23382 3040 23388 3052
rect 22612 3012 23388 3040
rect 22612 3000 22618 3012
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 24121 3043 24179 3049
rect 24121 3009 24133 3043
rect 24167 3040 24179 3043
rect 24210 3040 24216 3052
rect 24167 3012 24216 3040
rect 24167 3009 24179 3012
rect 24121 3003 24179 3009
rect 24210 3000 24216 3012
rect 24268 3000 24274 3052
rect 16942 2932 16948 2984
rect 17000 2972 17006 2984
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 17000 2944 17877 2972
rect 17000 2932 17006 2944
rect 17865 2941 17877 2944
rect 17911 2941 17923 2975
rect 17865 2935 17923 2941
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 20162 2972 20168 2984
rect 19659 2944 20168 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2941 21327 2975
rect 22186 2972 22192 2984
rect 22147 2944 22192 2972
rect 21269 2935 21327 2941
rect 10686 2904 10692 2916
rect 9508 2876 10692 2904
rect 10686 2864 10692 2876
rect 10744 2904 10750 2916
rect 10873 2907 10931 2913
rect 10873 2904 10885 2907
rect 10744 2876 10885 2904
rect 10744 2864 10750 2876
rect 10873 2873 10885 2876
rect 10919 2873 10931 2907
rect 10873 2867 10931 2873
rect 10965 2907 11023 2913
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 11882 2904 11888 2916
rect 11011 2876 11888 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 9674 2836 9680 2848
rect 9324 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 9950 2836 9956 2848
rect 9815 2808 9956 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 9950 2796 9956 2808
rect 10008 2836 10014 2848
rect 10597 2839 10655 2845
rect 10597 2836 10609 2839
rect 10008 2808 10609 2836
rect 10008 2796 10014 2808
rect 10597 2805 10609 2808
rect 10643 2836 10655 2839
rect 10980 2836 11008 2867
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 12529 2907 12587 2913
rect 12529 2873 12541 2907
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 10643 2808 11008 2836
rect 12544 2836 12572 2867
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 14550 2904 14556 2916
rect 12676 2876 12721 2904
rect 14511 2876 14556 2904
rect 12676 2864 12682 2876
rect 14550 2864 14556 2876
rect 14608 2864 14614 2916
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2873 14703 2907
rect 14645 2867 14703 2873
rect 15197 2907 15255 2913
rect 15197 2873 15209 2907
rect 15243 2904 15255 2907
rect 15746 2904 15752 2916
rect 15243 2876 15752 2904
rect 15243 2873 15255 2876
rect 15197 2867 15255 2873
rect 13538 2836 13544 2848
rect 12544 2808 13544 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 14660 2836 14688 2867
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16114 2904 16120 2916
rect 16075 2876 16120 2904
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 16209 2907 16267 2913
rect 16209 2873 16221 2907
rect 16255 2873 16267 2907
rect 16209 2867 16267 2873
rect 17313 2907 17371 2913
rect 17313 2873 17325 2907
rect 17359 2904 17371 2907
rect 18233 2907 18291 2913
rect 18233 2904 18245 2907
rect 17359 2876 18245 2904
rect 17359 2873 17371 2876
rect 17313 2867 17371 2873
rect 18233 2873 18245 2876
rect 18279 2904 18291 2907
rect 18506 2904 18512 2916
rect 18279 2876 18512 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 15562 2836 15568 2848
rect 14415 2808 15568 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 15562 2796 15568 2808
rect 15620 2836 15626 2848
rect 16224 2836 16252 2867
rect 18506 2864 18512 2876
rect 18564 2864 18570 2916
rect 18785 2907 18843 2913
rect 18785 2873 18797 2907
rect 18831 2873 18843 2907
rect 18785 2867 18843 2873
rect 20533 2907 20591 2913
rect 20533 2873 20545 2907
rect 20579 2904 20591 2907
rect 21174 2904 21180 2916
rect 20579 2876 21180 2904
rect 20579 2873 20591 2876
rect 20533 2867 20591 2873
rect 15620 2808 16252 2836
rect 17865 2839 17923 2845
rect 15620 2796 15626 2808
rect 17865 2805 17877 2839
rect 17911 2836 17923 2839
rect 18800 2836 18828 2867
rect 21174 2864 21180 2876
rect 21232 2904 21238 2916
rect 21284 2904 21312 2935
rect 22186 2932 22192 2944
rect 22244 2932 22250 2984
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2972 24639 2975
rect 24627 2944 25268 2972
rect 24627 2941 24639 2944
rect 24581 2935 24639 2941
rect 22278 2904 22284 2916
rect 21232 2876 22284 2904
rect 21232 2864 21238 2876
rect 22278 2864 22284 2876
rect 22336 2904 22342 2916
rect 22649 2907 22707 2913
rect 22649 2904 22661 2907
rect 22336 2876 22661 2904
rect 22336 2864 22342 2876
rect 22649 2873 22661 2876
rect 22695 2873 22707 2907
rect 22649 2867 22707 2873
rect 23477 2907 23535 2913
rect 23477 2873 23489 2907
rect 23523 2904 23535 2907
rect 24670 2904 24676 2916
rect 23523 2876 24676 2904
rect 23523 2873 23535 2876
rect 23477 2867 23535 2873
rect 24670 2864 24676 2876
rect 24728 2864 24734 2916
rect 25240 2848 25268 2944
rect 23014 2836 23020 2848
rect 17911 2808 18828 2836
rect 22975 2808 23020 2836
rect 17911 2805 17923 2808
rect 17865 2799 17923 2805
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 25222 2836 25228 2848
rect 25183 2808 25228 2836
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 3694 2592 3700 2644
rect 3752 2632 3758 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 3752 2604 6285 2632
rect 3752 2592 3758 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 6638 2632 6644 2644
rect 6599 2604 6644 2632
rect 6273 2595 6331 2601
rect 3234 2564 3240 2576
rect 3195 2536 3240 2564
rect 3234 2524 3240 2536
rect 3292 2524 3298 2576
rect 5074 2564 5080 2576
rect 5035 2536 5080 2564
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5721 2567 5779 2573
rect 5721 2533 5733 2567
rect 5767 2564 5779 2567
rect 5994 2564 6000 2576
rect 5767 2536 6000 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 1648 2499 1706 2505
rect 1648 2465 1660 2499
rect 1694 2496 1706 2499
rect 2038 2496 2044 2508
rect 1694 2468 2044 2496
rect 1694 2465 1706 2468
rect 1648 2459 1706 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2465 3086 2499
rect 3028 2459 3086 2465
rect 4868 2499 4926 2505
rect 4868 2465 4880 2499
rect 4914 2496 4926 2499
rect 6288 2496 6316 2595
rect 6638 2592 6644 2604
rect 6696 2632 6702 2644
rect 7653 2635 7711 2641
rect 6696 2604 7052 2632
rect 6696 2592 6702 2604
rect 6914 2496 6920 2508
rect 4914 2468 5396 2496
rect 6288 2468 6920 2496
rect 4914 2465 4926 2468
rect 4868 2459 4926 2465
rect 658 2388 664 2440
rect 716 2428 722 2440
rect 3043 2428 3071 2459
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 716 2400 3433 2428
rect 716 2388 722 2400
rect 3421 2397 3433 2400
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 1719 2363 1777 2369
rect 1719 2329 1731 2363
rect 1765 2360 1777 2363
rect 2958 2360 2964 2372
rect 1765 2332 2964 2360
rect 1765 2329 1777 2332
rect 1719 2323 1777 2329
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 2038 2292 2044 2304
rect 1999 2264 2044 2292
rect 2038 2252 2044 2264
rect 2096 2252 2102 2304
rect 5368 2301 5396 2468
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7024 2505 7052 2604
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 7834 2632 7840 2644
rect 7699 2604 7840 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 9125 2635 9183 2641
rect 8067 2604 8340 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8312 2573 8340 2604
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9171 2604 9628 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 8297 2567 8355 2573
rect 8297 2533 8309 2567
rect 8343 2564 8355 2567
rect 9214 2564 9220 2576
rect 8343 2536 9220 2564
rect 8343 2533 8355 2536
rect 8297 2527 8355 2533
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 9600 2564 9628 2604
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 9732 2604 10793 2632
rect 9732 2592 9738 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 10781 2595 10839 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 12342 2592 12348 2604
rect 12400 2632 12406 2644
rect 16390 2632 16396 2644
rect 12400 2604 12848 2632
rect 12400 2592 12406 2604
rect 9950 2564 9956 2576
rect 9600 2536 9956 2564
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 12820 2573 12848 2604
rect 13786 2604 16396 2632
rect 11241 2567 11299 2573
rect 11241 2564 11253 2567
rect 10100 2536 11253 2564
rect 10100 2524 10106 2536
rect 11241 2533 11253 2536
rect 11287 2564 11299 2567
rect 12713 2567 12771 2573
rect 12713 2564 12725 2567
rect 11287 2536 12725 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 12713 2533 12725 2536
rect 12759 2533 12771 2567
rect 12713 2527 12771 2533
rect 12805 2567 12863 2573
rect 12805 2533 12817 2567
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 13538 2564 13544 2576
rect 13403 2536 13544 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 13538 2524 13544 2536
rect 13596 2524 13602 2576
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 7009 2459 7067 2465
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 5859 2400 7052 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 7024 2360 7052 2400
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7156 2400 8217 2428
rect 7156 2388 7162 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 8205 2391 8263 2397
rect 8404 2400 9505 2428
rect 8404 2360 8432 2400
rect 9493 2397 9505 2400
rect 9539 2428 9551 2431
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9539 2400 9873 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9861 2391 9919 2397
rect 10060 2400 10149 2428
rect 8754 2360 8760 2372
rect 7024 2332 8432 2360
rect 8667 2332 8760 2360
rect 8754 2320 8760 2332
rect 8812 2360 8818 2372
rect 10060 2360 10088 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 13786 2428 13814 2604
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 17313 2635 17371 2641
rect 17313 2601 17325 2635
rect 17359 2632 17371 2635
rect 19518 2632 19524 2644
rect 17359 2604 19524 2632
rect 17359 2601 17371 2604
rect 17313 2595 17371 2601
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 20990 2592 20996 2644
rect 21048 2632 21054 2644
rect 23017 2635 23075 2641
rect 23017 2632 23029 2635
rect 21048 2604 23029 2632
rect 21048 2592 21054 2604
rect 23017 2601 23029 2604
rect 23063 2601 23075 2635
rect 23017 2595 23075 2601
rect 15289 2567 15347 2573
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15335 2536 15669 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15657 2533 15669 2536
rect 15703 2564 15715 2567
rect 15930 2564 15936 2576
rect 15703 2536 15936 2564
rect 15703 2533 15715 2536
rect 15657 2527 15715 2533
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2564 17831 2567
rect 18506 2564 18512 2576
rect 17819 2536 18512 2564
rect 17819 2533 17831 2536
rect 17773 2527 17831 2533
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 18782 2524 18788 2576
rect 18840 2564 18846 2576
rect 19705 2567 19763 2573
rect 19705 2564 19717 2567
rect 18840 2536 19717 2564
rect 18840 2524 18846 2536
rect 19705 2533 19717 2536
rect 19751 2533 19763 2567
rect 19705 2527 19763 2533
rect 21913 2567 21971 2573
rect 21913 2533 21925 2567
rect 21959 2564 21971 2567
rect 22186 2564 22192 2576
rect 21959 2536 22192 2564
rect 21959 2533 21971 2536
rect 21913 2527 21971 2533
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 14182 2456 14188 2468
rect 14240 2496 14246 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14240 2468 14749 2496
rect 14240 2456 14246 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 14737 2459 14795 2465
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 19720 2496 19748 2527
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 24670 2524 24676 2576
rect 24728 2564 24734 2576
rect 24765 2567 24823 2573
rect 24765 2564 24777 2567
rect 24728 2536 24777 2564
rect 24728 2524 24734 2536
rect 24765 2533 24777 2536
rect 24811 2533 24823 2567
rect 24765 2527 24823 2533
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19720 2468 19901 2496
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 21174 2496 21180 2508
rect 21039 2468 21180 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 21358 2456 21364 2508
rect 21416 2496 21422 2508
rect 21453 2499 21511 2505
rect 21453 2496 21465 2499
rect 21416 2468 21465 2496
rect 21416 2456 21422 2468
rect 21453 2465 21465 2468
rect 21499 2496 21511 2499
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 21499 2468 22293 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22738 2496 22744 2508
rect 22699 2468 22744 2496
rect 22281 2459 22339 2465
rect 22738 2456 22744 2468
rect 22796 2496 22802 2508
rect 23201 2499 23259 2505
rect 23201 2496 23213 2499
rect 22796 2468 23213 2496
rect 22796 2456 22802 2468
rect 23201 2465 23213 2468
rect 23247 2465 23259 2499
rect 23845 2499 23903 2505
rect 23845 2496 23857 2499
rect 23201 2459 23259 2465
rect 23446 2468 23857 2496
rect 10137 2391 10195 2397
rect 12820 2400 13814 2428
rect 8812 2332 10088 2360
rect 11609 2363 11667 2369
rect 8812 2320 8818 2332
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 12820 2360 12848 2400
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13964 2400 14105 2428
rect 13964 2388 13970 2400
rect 14093 2397 14105 2400
rect 14139 2428 14151 2431
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 14139 2400 15577 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 15746 2388 15752 2440
rect 15804 2428 15810 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15804 2400 16037 2428
rect 15804 2388 15810 2400
rect 16025 2397 16037 2400
rect 16071 2428 16083 2431
rect 18141 2431 18199 2437
rect 16071 2400 16988 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 11655 2332 12848 2360
rect 13725 2363 13783 2369
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 13725 2329 13737 2363
rect 13771 2360 13783 2363
rect 13998 2360 14004 2372
rect 13771 2332 14004 2360
rect 13771 2329 13783 2332
rect 13725 2323 13783 2329
rect 13998 2320 14004 2332
rect 14056 2360 14062 2372
rect 15764 2360 15792 2388
rect 14056 2332 15792 2360
rect 14056 2320 14062 2332
rect 16206 2320 16212 2372
rect 16264 2360 16270 2372
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 16264 2332 16865 2360
rect 16264 2320 16270 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 16960 2360 16988 2400
rect 18141 2397 18153 2431
rect 18187 2428 18199 2431
rect 18414 2428 18420 2440
rect 18187 2400 18420 2428
rect 18187 2397 18199 2400
rect 18141 2391 18199 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18524 2400 18705 2428
rect 18524 2360 18552 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 21266 2428 21272 2440
rect 20671 2400 21272 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 21266 2388 21272 2400
rect 21324 2428 21330 2440
rect 22094 2428 22100 2440
rect 21324 2400 22100 2428
rect 21324 2388 21330 2400
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 16960 2332 18552 2360
rect 16853 2323 16911 2329
rect 19242 2320 19248 2372
rect 19300 2360 19306 2372
rect 20073 2363 20131 2369
rect 20073 2360 20085 2363
rect 19300 2332 20085 2360
rect 19300 2320 19306 2332
rect 20073 2329 20085 2332
rect 20119 2329 20131 2363
rect 20073 2323 20131 2329
rect 21634 2320 21640 2372
rect 21692 2360 21698 2372
rect 23446 2360 23474 2468
rect 23845 2465 23857 2468
rect 23891 2496 23903 2499
rect 24121 2499 24179 2505
rect 24121 2496 24133 2499
rect 23891 2468 24133 2496
rect 23891 2465 23903 2468
rect 23845 2459 23903 2465
rect 24121 2465 24133 2468
rect 24167 2465 24179 2499
rect 24121 2459 24179 2465
rect 25660 2499 25718 2505
rect 25660 2465 25672 2499
rect 25706 2496 25718 2499
rect 26142 2496 26148 2508
rect 25706 2468 26148 2496
rect 25706 2465 25718 2468
rect 25660 2459 25718 2465
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 25731 2363 25789 2369
rect 25731 2360 25743 2363
rect 21692 2332 23474 2360
rect 23676 2332 25743 2360
rect 21692 2320 21698 2332
rect 5353 2295 5411 2301
rect 5353 2261 5365 2295
rect 5399 2292 5411 2295
rect 5534 2292 5540 2304
rect 5399 2264 5540 2292
rect 5399 2261 5411 2264
rect 5353 2255 5411 2261
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 7190 2292 7196 2304
rect 7151 2264 7196 2292
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 14369 2295 14427 2301
rect 14369 2261 14381 2295
rect 14415 2292 14427 2295
rect 14458 2292 14464 2304
rect 14415 2264 14464 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 16482 2292 16488 2304
rect 16443 2264 16488 2292
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 17184 2264 19349 2292
rect 17184 2252 17190 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 22922 2292 22928 2304
rect 22883 2264 22928 2292
rect 19337 2255 19395 2261
rect 22922 2252 22928 2264
rect 22980 2252 22986 2304
rect 23017 2295 23075 2301
rect 23017 2261 23029 2295
rect 23063 2292 23075 2295
rect 23676 2292 23704 2332
rect 25731 2329 25743 2332
rect 25777 2329 25789 2363
rect 25731 2323 25789 2329
rect 26142 2292 26148 2304
rect 23063 2264 23704 2292
rect 26103 2264 26148 2292
rect 23063 2261 23075 2264
rect 23017 2255 23075 2261
rect 26142 2252 26148 2264
rect 26200 2252 26206 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 4246 2048 4252 2100
rect 4304 2088 4310 2100
rect 12526 2088 12532 2100
rect 4304 2060 12532 2088
rect 4304 2048 4310 2060
rect 12526 2048 12532 2060
rect 12584 2048 12590 2100
rect 7190 76 7196 128
rect 7248 116 7254 128
rect 13538 116 13544 128
rect 7248 88 13544 116
rect 7248 76 7254 88
rect 13538 76 13544 88
rect 13596 76 13602 128
rect 9674 8 9680 60
rect 9732 48 9738 60
rect 10778 48 10784 60
rect 9732 20 10784 48
rect 9732 8 9738 20
rect 10778 8 10784 20
rect 10836 8 10842 60
<< via1 >>
rect 8300 27480 8352 27532
rect 9036 27480 9088 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 26240 24896 26292 24948
rect 6920 24760 6972 24812
rect 12348 24760 12400 24812
rect 23480 24692 23532 24744
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 20904 24352 20956 24404
rect 27344 24352 27396 24404
rect 4712 24216 4764 24268
rect 8116 24216 8168 24268
rect 17684 24216 17736 24268
rect 19156 24216 19208 24268
rect 19984 24216 20036 24268
rect 23112 24259 23164 24268
rect 23112 24225 23121 24259
rect 23121 24225 23155 24259
rect 23155 24225 23164 24259
rect 23112 24216 23164 24225
rect 25136 24216 25188 24268
rect 24860 24080 24912 24132
rect 8024 24012 8076 24064
rect 18880 24012 18932 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2872 23851 2924 23860
rect 2872 23817 2881 23851
rect 2881 23817 2915 23851
rect 2915 23817 2924 23851
rect 2872 23808 2924 23817
rect 3884 23851 3936 23860
rect 3884 23817 3893 23851
rect 3893 23817 3927 23851
rect 3927 23817 3936 23851
rect 3884 23808 3936 23817
rect 8116 23851 8168 23860
rect 8116 23817 8125 23851
rect 8125 23817 8159 23851
rect 8159 23817 8168 23851
rect 8116 23808 8168 23817
rect 19524 23808 19576 23860
rect 21916 23808 21968 23860
rect 24124 23808 24176 23860
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 1492 23740 1544 23792
rect 480 23604 532 23656
rect 2872 23604 2924 23656
rect 3884 23604 3936 23656
rect 6184 23740 6236 23792
rect 7932 23604 7984 23656
rect 18512 23740 18564 23792
rect 19156 23783 19208 23792
rect 19156 23749 19165 23783
rect 19165 23749 19199 23783
rect 19199 23749 19208 23783
rect 19156 23740 19208 23749
rect 22744 23740 22796 23792
rect 12348 23604 12400 23656
rect 15568 23604 15620 23656
rect 6736 23536 6788 23588
rect 7840 23536 7892 23588
rect 12072 23536 12124 23588
rect 17316 23604 17368 23656
rect 17500 23536 17552 23588
rect 20904 23604 20956 23656
rect 20812 23536 20864 23588
rect 2412 23468 2464 23520
rect 2688 23468 2740 23520
rect 6828 23468 6880 23520
rect 12164 23468 12216 23520
rect 19984 23468 20036 23520
rect 20720 23468 20772 23520
rect 23112 23468 23164 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 25596 23128 25648 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 25228 22720 25280 22772
rect 24124 22380 24176 22432
rect 25596 22380 25648 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 25504 21292 25556 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 20812 21088 20864 21140
rect 22008 21088 22060 21140
rect 11152 21020 11204 21072
rect 14832 21020 14884 21072
rect 20812 20952 20864 21004
rect 20168 20748 20220 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 24768 20587 24820 20596
rect 24768 20553 24777 20587
rect 24777 20553 24811 20587
rect 24811 20553 24820 20587
rect 24768 20544 24820 20553
rect 19340 20340 19392 20392
rect 24584 20383 24636 20392
rect 24584 20349 24593 20383
rect 24593 20349 24627 20383
rect 24627 20349 24636 20383
rect 24584 20340 24636 20349
rect 19524 20204 19576 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 20812 20204 20864 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 12532 20000 12584 20052
rect 13360 20000 13412 20052
rect 18880 20000 18932 20052
rect 20076 20000 20128 20052
rect 24584 20000 24636 20052
rect 15936 19864 15988 19916
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 19064 19796 19116 19848
rect 19984 19796 20036 19848
rect 22560 19864 22612 19916
rect 23848 19864 23900 19916
rect 16304 19660 16356 19712
rect 19248 19660 19300 19712
rect 21180 19703 21232 19712
rect 21180 19669 21189 19703
rect 21189 19669 21223 19703
rect 21223 19669 21232 19703
rect 21180 19660 21232 19669
rect 22468 19660 22520 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 16948 19499 17000 19508
rect 16948 19465 16957 19499
rect 16957 19465 16991 19499
rect 16991 19465 17000 19499
rect 16948 19456 17000 19465
rect 19064 19456 19116 19508
rect 22560 19499 22612 19508
rect 22560 19465 22569 19499
rect 22569 19465 22603 19499
rect 22603 19465 22612 19499
rect 22560 19456 22612 19465
rect 24768 19499 24820 19508
rect 24768 19465 24777 19499
rect 24777 19465 24811 19499
rect 24811 19465 24820 19499
rect 24768 19456 24820 19465
rect 16028 19388 16080 19440
rect 17500 19388 17552 19440
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 20260 19320 20312 19372
rect 20996 19363 21048 19372
rect 20996 19329 21005 19363
rect 21005 19329 21039 19363
rect 21039 19329 21048 19363
rect 20996 19320 21048 19329
rect 16948 19252 17000 19304
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 21640 19295 21692 19304
rect 21640 19261 21649 19295
rect 21649 19261 21683 19295
rect 21683 19261 21692 19295
rect 21640 19252 21692 19261
rect 24860 19252 24912 19304
rect 20720 19227 20772 19236
rect 16488 19116 16540 19168
rect 18604 19159 18656 19168
rect 18604 19125 18613 19159
rect 18613 19125 18647 19159
rect 18647 19125 18656 19159
rect 18604 19116 18656 19125
rect 20720 19193 20729 19227
rect 20729 19193 20763 19227
rect 20763 19193 20772 19227
rect 20720 19184 20772 19193
rect 21180 19184 21232 19236
rect 21548 19227 21600 19236
rect 21548 19193 21557 19227
rect 21557 19193 21591 19227
rect 21591 19193 21600 19227
rect 21548 19184 21600 19193
rect 23848 19159 23900 19168
rect 23848 19125 23857 19159
rect 23857 19125 23891 19159
rect 23891 19125 23900 19159
rect 23848 19116 23900 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 19248 18912 19300 18964
rect 16488 18844 16540 18896
rect 17132 18887 17184 18896
rect 17132 18853 17141 18887
rect 17141 18853 17175 18887
rect 17175 18853 17184 18887
rect 17132 18844 17184 18853
rect 17408 18844 17460 18896
rect 19432 18887 19484 18896
rect 19432 18853 19441 18887
rect 19441 18853 19475 18887
rect 19475 18853 19484 18887
rect 19432 18844 19484 18853
rect 20444 18844 20496 18896
rect 20996 18887 21048 18896
rect 20996 18853 21005 18887
rect 21005 18853 21039 18887
rect 21039 18853 21048 18887
rect 20996 18844 21048 18853
rect 21180 18844 21232 18896
rect 16120 18776 16172 18828
rect 23020 18776 23072 18828
rect 24768 18776 24820 18828
rect 17224 18708 17276 18760
rect 20720 18708 20772 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 18144 18572 18196 18624
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 24216 18572 24268 18624
rect 24676 18572 24728 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 21548 18411 21600 18420
rect 21548 18377 21557 18411
rect 21557 18377 21591 18411
rect 21591 18377 21600 18411
rect 21548 18368 21600 18377
rect 25412 18411 25464 18420
rect 25412 18377 25421 18411
rect 25421 18377 25455 18411
rect 25455 18377 25464 18411
rect 25412 18368 25464 18377
rect 9680 18300 9732 18352
rect 13544 18300 13596 18352
rect 12808 18232 12860 18284
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 18512 18275 18564 18284
rect 18512 18241 18521 18275
rect 18521 18241 18555 18275
rect 18555 18241 18564 18275
rect 18512 18232 18564 18241
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 21456 18232 21508 18284
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 23020 18275 23072 18284
rect 22192 18232 22244 18241
rect 23020 18241 23029 18275
rect 23029 18241 23063 18275
rect 23063 18241 23072 18275
rect 23020 18232 23072 18241
rect 12256 18164 12308 18216
rect 14464 18207 14516 18216
rect 14464 18173 14482 18207
rect 14482 18173 14516 18207
rect 14464 18164 14516 18173
rect 13544 18096 13596 18148
rect 14372 18028 14424 18080
rect 15384 18028 15436 18080
rect 15844 18028 15896 18080
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 17960 18028 18012 18080
rect 19432 18096 19484 18148
rect 20260 18139 20312 18148
rect 20260 18105 20269 18139
rect 20269 18105 20303 18139
rect 20303 18105 20312 18139
rect 20260 18096 20312 18105
rect 21548 18028 21600 18080
rect 23112 18096 23164 18148
rect 24216 18164 24268 18216
rect 25136 18096 25188 18148
rect 24032 18028 24084 18080
rect 24584 18028 24636 18080
rect 24768 18028 24820 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 17132 17824 17184 17876
rect 18144 17824 18196 17876
rect 20168 17867 20220 17876
rect 20168 17833 20177 17867
rect 20177 17833 20211 17867
rect 20211 17833 20220 17867
rect 20168 17824 20220 17833
rect 20996 17824 21048 17876
rect 24124 17867 24176 17876
rect 24124 17833 24133 17867
rect 24133 17833 24167 17867
rect 24167 17833 24176 17867
rect 24124 17824 24176 17833
rect 27528 17824 27580 17876
rect 13084 17799 13136 17808
rect 13084 17765 13093 17799
rect 13093 17765 13127 17799
rect 13127 17765 13136 17799
rect 13084 17756 13136 17765
rect 13176 17799 13228 17808
rect 13176 17765 13185 17799
rect 13185 17765 13219 17799
rect 13219 17765 13228 17799
rect 13176 17756 13228 17765
rect 17408 17756 17460 17808
rect 18604 17799 18656 17808
rect 18604 17765 18613 17799
rect 18613 17765 18647 17799
rect 18647 17765 18656 17799
rect 18604 17756 18656 17765
rect 21640 17799 21692 17808
rect 21640 17765 21649 17799
rect 21649 17765 21683 17799
rect 21683 17765 21692 17799
rect 21640 17756 21692 17765
rect 22192 17799 22244 17808
rect 22192 17765 22201 17799
rect 22201 17765 22235 17799
rect 22235 17765 22244 17799
rect 22192 17756 22244 17765
rect 23112 17756 23164 17808
rect 8300 17688 8352 17740
rect 9128 17688 9180 17740
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 24676 17688 24728 17740
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 20720 17620 20772 17672
rect 22192 17620 22244 17672
rect 23572 17663 23624 17672
rect 13636 17595 13688 17604
rect 13636 17561 13645 17595
rect 13645 17561 13679 17595
rect 13679 17561 13688 17595
rect 13636 17552 13688 17561
rect 14372 17552 14424 17604
rect 23572 17629 23581 17663
rect 23581 17629 23615 17663
rect 23615 17629 23624 17663
rect 23572 17620 23624 17629
rect 23388 17552 23440 17604
rect 16488 17527 16540 17536
rect 16488 17493 16497 17527
rect 16497 17493 16531 17527
rect 16531 17493 16540 17527
rect 16488 17484 16540 17493
rect 18512 17484 18564 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 13084 17280 13136 17332
rect 15568 17280 15620 17332
rect 15844 17323 15896 17332
rect 15844 17289 15853 17323
rect 15853 17289 15887 17323
rect 15887 17289 15896 17323
rect 17408 17323 17460 17332
rect 15844 17280 15896 17289
rect 13176 17212 13228 17264
rect 13636 17255 13688 17264
rect 13636 17221 13645 17255
rect 13645 17221 13679 17255
rect 13679 17221 13688 17255
rect 13636 17212 13688 17221
rect 12164 17144 12216 17196
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 18604 17280 18656 17332
rect 21640 17280 21692 17332
rect 22192 17280 22244 17332
rect 23112 17323 23164 17332
rect 23112 17289 23121 17323
rect 23121 17289 23155 17323
rect 23155 17289 23164 17323
rect 23112 17280 23164 17289
rect 23388 17323 23440 17332
rect 23388 17289 23397 17323
rect 23397 17289 23431 17323
rect 23431 17289 23440 17323
rect 23388 17280 23440 17289
rect 24676 17280 24728 17332
rect 17224 17144 17276 17196
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 19156 17187 19208 17196
rect 19156 17153 19165 17187
rect 19165 17153 19199 17187
rect 19199 17153 19208 17187
rect 19156 17144 19208 17153
rect 19248 17144 19300 17196
rect 15936 17076 15988 17128
rect 20996 17076 21048 17128
rect 24124 17144 24176 17196
rect 16488 17008 16540 17060
rect 17960 17008 18012 17060
rect 18604 17051 18656 17060
rect 18604 17017 18613 17051
rect 18613 17017 18647 17051
rect 18647 17017 18656 17051
rect 18604 17008 18656 17017
rect 20536 17008 20588 17060
rect 21272 17051 21324 17060
rect 21272 17017 21275 17051
rect 21275 17017 21309 17051
rect 21309 17017 21324 17051
rect 21272 17008 21324 17017
rect 23020 17008 23072 17060
rect 24032 17008 24084 17060
rect 24768 17008 24820 17060
rect 14740 16940 14792 16992
rect 18420 16940 18472 16992
rect 20168 16940 20220 16992
rect 24492 16940 24544 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 11152 16779 11204 16788
rect 11152 16745 11161 16779
rect 11161 16745 11195 16779
rect 11195 16745 11204 16779
rect 11152 16736 11204 16745
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 17960 16779 18012 16788
rect 17960 16745 17969 16779
rect 17969 16745 18003 16779
rect 18003 16745 18012 16779
rect 17960 16736 18012 16745
rect 18604 16736 18656 16788
rect 20260 16736 20312 16788
rect 22100 16736 22152 16788
rect 24032 16779 24084 16788
rect 6828 16668 6880 16720
rect 8116 16711 8168 16720
rect 8116 16677 8125 16711
rect 8125 16677 8159 16711
rect 8159 16677 8168 16711
rect 8116 16668 8168 16677
rect 8208 16711 8260 16720
rect 8208 16677 8217 16711
rect 8217 16677 8251 16711
rect 8251 16677 8260 16711
rect 13176 16711 13228 16720
rect 8208 16668 8260 16677
rect 13176 16677 13185 16711
rect 13185 16677 13219 16711
rect 13219 16677 13228 16711
rect 13176 16668 13228 16677
rect 17776 16668 17828 16720
rect 19156 16668 19208 16720
rect 19524 16668 19576 16720
rect 19984 16711 20036 16720
rect 19984 16677 19993 16711
rect 19993 16677 20027 16711
rect 20027 16677 20036 16711
rect 19984 16668 20036 16677
rect 21272 16668 21324 16720
rect 23020 16711 23072 16720
rect 23020 16677 23029 16711
rect 23029 16677 23063 16711
rect 23063 16677 23072 16711
rect 23020 16668 23072 16677
rect 24032 16745 24041 16779
rect 24041 16745 24075 16779
rect 24075 16745 24084 16779
rect 24032 16736 24084 16745
rect 23572 16711 23624 16720
rect 23572 16677 23581 16711
rect 23581 16677 23615 16711
rect 23615 16677 23624 16711
rect 23572 16668 23624 16677
rect 24492 16711 24544 16720
rect 24492 16677 24501 16711
rect 24501 16677 24535 16711
rect 24535 16677 24544 16711
rect 24492 16668 24544 16677
rect 25136 16668 25188 16720
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 11796 16600 11848 16652
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 16212 16575 16264 16584
rect 6736 16464 6788 16516
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 17500 16532 17552 16584
rect 18604 16532 18656 16584
rect 13452 16464 13504 16516
rect 13636 16507 13688 16516
rect 13636 16473 13645 16507
rect 13645 16473 13679 16507
rect 13679 16473 13688 16507
rect 13636 16464 13688 16473
rect 15568 16464 15620 16516
rect 22192 16532 22244 16584
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 9772 16396 9824 16448
rect 14004 16439 14056 16448
rect 14004 16405 14013 16439
rect 14013 16405 14047 16439
rect 14047 16405 14056 16439
rect 14004 16396 14056 16405
rect 18144 16396 18196 16448
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 20720 16439 20772 16448
rect 20720 16405 20729 16439
rect 20729 16405 20763 16439
rect 20763 16405 20772 16439
rect 20720 16396 20772 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 8116 16192 8168 16244
rect 13268 16192 13320 16244
rect 14096 16192 14148 16244
rect 22192 16192 22244 16244
rect 23020 16235 23072 16244
rect 23020 16201 23029 16235
rect 23029 16201 23063 16235
rect 23063 16201 23072 16235
rect 23020 16192 23072 16201
rect 25136 16235 25188 16244
rect 25136 16201 25145 16235
rect 25145 16201 25179 16235
rect 25179 16201 25188 16235
rect 25136 16192 25188 16201
rect 7472 16124 7524 16176
rect 8208 16124 8260 16176
rect 10140 16167 10192 16176
rect 10140 16133 10149 16167
rect 10149 16133 10183 16167
rect 10183 16133 10192 16167
rect 10140 16124 10192 16133
rect 13360 16124 13412 16176
rect 13452 16167 13504 16176
rect 13452 16133 13461 16167
rect 13461 16133 13495 16167
rect 13495 16133 13504 16167
rect 19156 16167 19208 16176
rect 13452 16124 13504 16133
rect 19156 16133 19165 16167
rect 19165 16133 19199 16167
rect 19199 16133 19208 16167
rect 19156 16124 19208 16133
rect 21916 16124 21968 16176
rect 8024 16099 8076 16108
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 8024 16056 8076 16065
rect 9772 16056 9824 16108
rect 11336 16056 11388 16108
rect 12256 16056 12308 16108
rect 14004 16099 14056 16108
rect 14004 16065 14013 16099
rect 14013 16065 14047 16099
rect 14047 16065 14056 16099
rect 14004 16056 14056 16065
rect 15292 16056 15344 16108
rect 15568 16099 15620 16108
rect 15568 16065 15577 16099
rect 15577 16065 15611 16099
rect 15611 16065 15620 16099
rect 15568 16056 15620 16065
rect 18604 16056 18656 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 22100 16099 22152 16108
rect 22100 16065 22109 16099
rect 22109 16065 22143 16099
rect 22143 16065 22152 16099
rect 22100 16056 22152 16065
rect 24768 16124 24820 16176
rect 24308 16056 24360 16108
rect 8760 15920 8812 15972
rect 10048 15920 10100 15972
rect 11244 15920 11296 15972
rect 19984 16031 20036 16040
rect 13176 15920 13228 15972
rect 13820 15920 13872 15972
rect 14096 15963 14148 15972
rect 14096 15929 14105 15963
rect 14105 15929 14139 15963
rect 14139 15929 14148 15963
rect 14648 15963 14700 15972
rect 14096 15920 14148 15929
rect 14648 15929 14657 15963
rect 14657 15929 14691 15963
rect 14691 15929 14700 15963
rect 14648 15920 14700 15929
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 14832 15852 14884 15904
rect 15936 15920 15988 15972
rect 17500 15963 17552 15972
rect 17500 15929 17509 15963
rect 17509 15929 17543 15963
rect 17543 15929 17552 15963
rect 17500 15920 17552 15929
rect 16120 15852 16172 15904
rect 16672 15852 16724 15904
rect 17776 15852 17828 15904
rect 19524 15920 19576 15972
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20168 16031 20220 16040
rect 20168 15997 20177 16031
rect 20177 15997 20211 16031
rect 20211 15997 20220 16031
rect 20168 15988 20220 15997
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 22192 15963 22244 15972
rect 22192 15929 22201 15963
rect 22201 15929 22235 15963
rect 22235 15929 22244 15963
rect 22192 15920 22244 15929
rect 24216 15920 24268 15972
rect 20812 15852 20864 15904
rect 24124 15852 24176 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 7840 15691 7892 15700
rect 7840 15657 7849 15691
rect 7849 15657 7883 15691
rect 7883 15657 7892 15691
rect 7840 15648 7892 15657
rect 9772 15648 9824 15700
rect 10140 15648 10192 15700
rect 13360 15648 13412 15700
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 8208 15623 8260 15632
rect 8208 15589 8217 15623
rect 8217 15589 8251 15623
rect 8251 15589 8260 15623
rect 11060 15623 11112 15632
rect 8208 15580 8260 15589
rect 11060 15589 11069 15623
rect 11069 15589 11103 15623
rect 11103 15589 11112 15623
rect 11060 15580 11112 15589
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 13820 15580 13872 15589
rect 14004 15580 14056 15632
rect 14648 15580 14700 15632
rect 14740 15580 14792 15632
rect 17500 15580 17552 15632
rect 18696 15580 18748 15632
rect 19524 15648 19576 15700
rect 20536 15648 20588 15700
rect 20996 15691 21048 15700
rect 20996 15657 21005 15691
rect 21005 15657 21039 15691
rect 21039 15657 21048 15691
rect 20996 15648 21048 15657
rect 24032 15648 24084 15700
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 25136 15691 25188 15700
rect 25136 15657 25145 15691
rect 25145 15657 25179 15691
rect 25179 15657 25188 15691
rect 25136 15648 25188 15657
rect 9588 15555 9640 15564
rect 9588 15521 9597 15555
rect 9597 15521 9631 15555
rect 9631 15521 9640 15555
rect 9588 15512 9640 15521
rect 12716 15512 12768 15564
rect 8760 15487 8812 15496
rect 8760 15453 8769 15487
rect 8769 15453 8803 15487
rect 8803 15453 8812 15487
rect 10968 15487 11020 15496
rect 8760 15444 8812 15453
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 15384 15512 15436 15564
rect 19432 15512 19484 15564
rect 20168 15580 20220 15632
rect 20444 15580 20496 15632
rect 23388 15580 23440 15632
rect 24676 15580 24728 15632
rect 15660 15444 15712 15496
rect 17132 15444 17184 15496
rect 18880 15444 18932 15496
rect 20812 15512 20864 15564
rect 21732 15555 21784 15564
rect 20352 15444 20404 15496
rect 21732 15521 21741 15555
rect 21741 15521 21775 15555
rect 21775 15521 21784 15555
rect 21732 15512 21784 15521
rect 21824 15512 21876 15564
rect 24952 15555 25004 15564
rect 24952 15521 24961 15555
rect 24961 15521 24995 15555
rect 24995 15521 25004 15555
rect 24952 15512 25004 15521
rect 20168 15376 20220 15428
rect 21088 15376 21140 15428
rect 22928 15444 22980 15496
rect 13084 15351 13136 15360
rect 13084 15317 13093 15351
rect 13093 15317 13127 15351
rect 13127 15317 13136 15351
rect 13084 15308 13136 15317
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 20812 15308 20864 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 9588 15104 9640 15156
rect 10876 15104 10928 15156
rect 11060 15104 11112 15156
rect 11980 15104 12032 15156
rect 12440 15104 12492 15156
rect 12716 15147 12768 15156
rect 12716 15113 12725 15147
rect 12725 15113 12759 15147
rect 12759 15113 12768 15147
rect 12716 15104 12768 15113
rect 13912 15104 13964 15156
rect 15384 15104 15436 15156
rect 19432 15104 19484 15156
rect 20168 15104 20220 15156
rect 22192 15104 22244 15156
rect 23940 15104 23992 15156
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 14832 15036 14884 15088
rect 15660 15036 15712 15088
rect 17684 15036 17736 15088
rect 20720 15036 20772 15088
rect 21916 15036 21968 15088
rect 23388 15079 23440 15088
rect 23388 15045 23397 15079
rect 23397 15045 23431 15079
rect 23431 15045 23440 15079
rect 23388 15036 23440 15045
rect 10140 14968 10192 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 14648 14968 14700 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 18420 14968 18472 15020
rect 18880 14968 18932 15020
rect 11336 14900 11388 14952
rect 7380 14875 7432 14884
rect 7380 14841 7389 14875
rect 7389 14841 7423 14875
rect 7423 14841 7432 14875
rect 7380 14832 7432 14841
rect 7472 14875 7524 14884
rect 7472 14841 7481 14875
rect 7481 14841 7515 14875
rect 7515 14841 7524 14875
rect 7472 14832 7524 14841
rect 8944 14875 8996 14884
rect 8944 14841 8953 14875
rect 8953 14841 8987 14875
rect 8987 14841 8996 14875
rect 8944 14832 8996 14841
rect 9036 14875 9088 14884
rect 9036 14841 9045 14875
rect 9045 14841 9079 14875
rect 9079 14841 9088 14875
rect 9036 14832 9088 14841
rect 8208 14764 8260 14816
rect 11244 14832 11296 14884
rect 13636 14832 13688 14884
rect 14004 14900 14056 14952
rect 20812 14968 20864 15020
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 14924 14875 14976 14884
rect 14924 14841 14933 14875
rect 14933 14841 14967 14875
rect 14967 14841 14976 14875
rect 14924 14832 14976 14841
rect 16488 14875 16540 14884
rect 10692 14764 10744 14816
rect 12716 14764 12768 14816
rect 13912 14764 13964 14816
rect 14740 14764 14792 14816
rect 16488 14841 16497 14875
rect 16497 14841 16531 14875
rect 16531 14841 16540 14875
rect 16488 14832 16540 14841
rect 16672 14832 16724 14884
rect 17500 14875 17552 14884
rect 17500 14841 17509 14875
rect 17509 14841 17543 14875
rect 17543 14841 17552 14875
rect 17500 14832 17552 14841
rect 17960 14832 18012 14884
rect 18144 14875 18196 14884
rect 18144 14841 18153 14875
rect 18153 14841 18187 14875
rect 18187 14841 18196 14875
rect 18144 14832 18196 14841
rect 17868 14764 17920 14816
rect 19064 14832 19116 14884
rect 20628 14900 20680 14952
rect 20996 14900 21048 14952
rect 23664 14943 23716 14952
rect 21732 14832 21784 14884
rect 23664 14909 23673 14943
rect 23673 14909 23707 14943
rect 23707 14909 23716 14943
rect 23664 14900 23716 14909
rect 23112 14832 23164 14884
rect 18880 14764 18932 14816
rect 20352 14764 20404 14816
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 22192 14807 22244 14816
rect 22192 14773 22201 14807
rect 22201 14773 22235 14807
rect 22235 14773 22244 14807
rect 22192 14764 22244 14773
rect 24216 14900 24268 14952
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 8944 14560 8996 14612
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 11428 14603 11480 14612
rect 11428 14569 11437 14603
rect 11437 14569 11471 14603
rect 11471 14569 11480 14603
rect 11428 14560 11480 14569
rect 11980 14603 12032 14612
rect 11980 14569 11989 14603
rect 11989 14569 12023 14603
rect 12023 14569 12032 14603
rect 11980 14560 12032 14569
rect 12716 14560 12768 14612
rect 14924 14603 14976 14612
rect 14924 14569 14933 14603
rect 14933 14569 14967 14603
rect 14967 14569 14976 14603
rect 14924 14560 14976 14569
rect 15292 14560 15344 14612
rect 9036 14492 9088 14544
rect 13636 14492 13688 14544
rect 8852 14424 8904 14476
rect 11152 14424 11204 14476
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 15384 14467 15436 14476
rect 15384 14433 15402 14467
rect 15402 14433 15436 14467
rect 17316 14560 17368 14612
rect 17868 14560 17920 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 23664 14603 23716 14612
rect 16672 14535 16724 14544
rect 16672 14501 16681 14535
rect 16681 14501 16715 14535
rect 16715 14501 16724 14535
rect 16672 14492 16724 14501
rect 17224 14535 17276 14544
rect 17224 14501 17233 14535
rect 17233 14501 17267 14535
rect 17267 14501 17276 14535
rect 17224 14492 17276 14501
rect 18144 14492 18196 14544
rect 18236 14535 18288 14544
rect 18236 14501 18245 14535
rect 18245 14501 18279 14535
rect 18279 14501 18288 14535
rect 18236 14492 18288 14501
rect 21824 14492 21876 14544
rect 15384 14424 15436 14433
rect 19432 14424 19484 14476
rect 21732 14467 21784 14476
rect 21732 14433 21741 14467
rect 21741 14433 21775 14467
rect 21775 14433 21784 14467
rect 21732 14424 21784 14433
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 15476 14356 15528 14408
rect 17408 14356 17460 14408
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 18420 14356 18472 14365
rect 21088 14356 21140 14408
rect 22192 14424 22244 14476
rect 22376 14467 22428 14476
rect 22376 14433 22385 14467
rect 22385 14433 22419 14467
rect 22419 14433 22428 14467
rect 22376 14424 22428 14433
rect 23664 14569 23673 14603
rect 23673 14569 23707 14603
rect 23707 14569 23716 14603
rect 23664 14560 23716 14569
rect 24124 14603 24176 14612
rect 24124 14569 24133 14603
rect 24133 14569 24167 14603
rect 24167 14569 24176 14603
rect 24124 14560 24176 14569
rect 22836 14424 22888 14476
rect 23940 14467 23992 14476
rect 23940 14433 23949 14467
rect 23949 14433 23983 14467
rect 23983 14433 23992 14467
rect 23940 14424 23992 14433
rect 25412 14467 25464 14476
rect 25412 14433 25421 14467
rect 25421 14433 25455 14467
rect 25455 14433 25464 14467
rect 25412 14424 25464 14433
rect 18972 14288 19024 14340
rect 20076 14288 20128 14340
rect 20812 14288 20864 14340
rect 7932 14263 7984 14272
rect 7932 14229 7941 14263
rect 7941 14229 7975 14263
rect 7975 14229 7984 14263
rect 7932 14220 7984 14229
rect 9496 14220 9548 14272
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 18144 14220 18196 14272
rect 22928 14220 22980 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 10692 14016 10744 14068
rect 11152 14016 11204 14068
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 15476 14016 15528 14068
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 16396 14016 16448 14068
rect 18236 14016 18288 14068
rect 19340 14016 19392 14068
rect 19524 14016 19576 14068
rect 21088 14016 21140 14068
rect 22836 14016 22888 14068
rect 23940 14059 23992 14068
rect 23940 14025 23949 14059
rect 23949 14025 23983 14059
rect 23983 14025 23992 14059
rect 23940 14016 23992 14025
rect 24860 14016 24912 14068
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 6736 13812 6788 13864
rect 7932 13855 7984 13864
rect 7932 13821 7941 13855
rect 7941 13821 7975 13855
rect 7975 13821 7984 13855
rect 7932 13812 7984 13821
rect 11796 13948 11848 14000
rect 13084 13948 13136 14000
rect 14372 13948 14424 14000
rect 18972 13948 19024 14000
rect 20444 13948 20496 14000
rect 20904 13948 20956 14000
rect 25412 13948 25464 14000
rect 14648 13880 14700 13932
rect 16304 13880 16356 13932
rect 17224 13880 17276 13932
rect 19156 13880 19208 13932
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 8484 13676 8536 13728
rect 8852 13676 8904 13728
rect 10140 13744 10192 13796
rect 11428 13744 11480 13796
rect 11888 13787 11940 13796
rect 11888 13753 11897 13787
rect 11897 13753 11931 13787
rect 11931 13753 11940 13787
rect 11888 13744 11940 13753
rect 12256 13787 12308 13796
rect 12256 13753 12265 13787
rect 12265 13753 12299 13787
rect 12299 13753 12308 13787
rect 13084 13812 13136 13864
rect 17316 13812 17368 13864
rect 20812 13880 20864 13932
rect 19616 13812 19668 13864
rect 20076 13855 20128 13864
rect 20076 13821 20085 13855
rect 20085 13821 20119 13855
rect 20119 13821 20128 13855
rect 20076 13812 20128 13821
rect 13636 13787 13688 13796
rect 12256 13744 12308 13753
rect 13636 13753 13645 13787
rect 13645 13753 13679 13787
rect 13679 13753 13688 13787
rect 13636 13744 13688 13753
rect 14280 13744 14332 13796
rect 15936 13744 15988 13796
rect 16304 13744 16356 13796
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 17960 13676 18012 13728
rect 19340 13719 19392 13728
rect 19340 13685 19349 13719
rect 19349 13685 19383 13719
rect 19383 13685 19392 13719
rect 19340 13676 19392 13685
rect 20352 13812 20404 13864
rect 22008 13812 22060 13864
rect 24952 13812 25004 13864
rect 25504 13812 25556 13864
rect 21548 13719 21600 13728
rect 21548 13685 21557 13719
rect 21557 13685 21591 13719
rect 21591 13685 21600 13719
rect 21548 13676 21600 13685
rect 21732 13676 21784 13728
rect 22100 13676 22152 13728
rect 24216 13676 24268 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 8116 13472 8168 13524
rect 12808 13472 12860 13524
rect 13360 13472 13412 13524
rect 14372 13472 14424 13524
rect 16212 13472 16264 13524
rect 19524 13472 19576 13524
rect 21088 13472 21140 13524
rect 9036 13404 9088 13456
rect 15752 13447 15804 13456
rect 15752 13413 15761 13447
rect 15761 13413 15795 13447
rect 15795 13413 15804 13447
rect 15752 13404 15804 13413
rect 18788 13404 18840 13456
rect 25596 13472 25648 13524
rect 22928 13447 22980 13456
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 11980 13336 12032 13388
rect 12808 13336 12860 13388
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 17500 13336 17552 13388
rect 19340 13336 19392 13388
rect 21732 13379 21784 13388
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 9956 13268 10008 13320
rect 13176 13311 13228 13320
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 15476 13268 15528 13320
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16028 13268 16080 13320
rect 18144 13268 18196 13320
rect 18972 13268 19024 13320
rect 21732 13345 21741 13379
rect 21741 13345 21775 13379
rect 21775 13345 21784 13379
rect 21732 13336 21784 13345
rect 22928 13413 22937 13447
rect 22937 13413 22971 13447
rect 22971 13413 22980 13447
rect 22928 13404 22980 13413
rect 21548 13268 21600 13320
rect 22376 13336 22428 13388
rect 9680 13200 9732 13252
rect 11796 13200 11848 13252
rect 16120 13200 16172 13252
rect 24124 13379 24176 13388
rect 24124 13345 24133 13379
rect 24133 13345 24167 13379
rect 24167 13345 24176 13379
rect 24124 13336 24176 13345
rect 25780 13336 25832 13388
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 13820 13132 13872 13184
rect 14556 13132 14608 13184
rect 16672 13175 16724 13184
rect 16672 13141 16681 13175
rect 16681 13141 16715 13175
rect 16715 13141 16724 13175
rect 16672 13132 16724 13141
rect 18144 13132 18196 13184
rect 18880 13175 18932 13184
rect 18880 13141 18889 13175
rect 18889 13141 18923 13175
rect 18923 13141 18932 13175
rect 18880 13132 18932 13141
rect 20260 13175 20312 13184
rect 20260 13141 20269 13175
rect 20269 13141 20303 13175
rect 20303 13141 20312 13175
rect 20260 13132 20312 13141
rect 20352 13132 20404 13184
rect 20996 13132 21048 13184
rect 21732 13132 21784 13184
rect 22468 13132 22520 13184
rect 24032 13175 24084 13184
rect 24032 13141 24041 13175
rect 24041 13141 24075 13175
rect 24075 13141 24084 13175
rect 24032 13132 24084 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 9036 12928 9088 12980
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 14096 12928 14148 12980
rect 15752 12928 15804 12980
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 7840 12860 7892 12912
rect 12992 12860 13044 12912
rect 13268 12860 13320 12912
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 11244 12835 11296 12844
rect 8300 12792 8352 12801
rect 8392 12767 8444 12776
rect 6920 12656 6972 12708
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 13176 12792 13228 12844
rect 8484 12656 8536 12708
rect 10876 12699 10928 12708
rect 10876 12665 10885 12699
rect 10885 12665 10919 12699
rect 10919 12665 10928 12699
rect 10876 12656 10928 12665
rect 12808 12699 12860 12708
rect 7840 12588 7892 12640
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 12808 12665 12817 12699
rect 12817 12665 12851 12699
rect 12851 12665 12860 12699
rect 12808 12656 12860 12665
rect 13636 12656 13688 12708
rect 11428 12588 11480 12640
rect 11980 12588 12032 12640
rect 12900 12588 12952 12640
rect 15200 12792 15252 12844
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 17408 12792 17460 12844
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 20628 12792 20680 12844
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 18972 12724 19024 12776
rect 19156 12724 19208 12776
rect 19524 12724 19576 12776
rect 18880 12588 18932 12640
rect 19340 12631 19392 12640
rect 19340 12597 19349 12631
rect 19349 12597 19383 12631
rect 19383 12597 19392 12631
rect 19340 12588 19392 12597
rect 20352 12724 20404 12776
rect 22100 12699 22152 12708
rect 22100 12665 22109 12699
rect 22109 12665 22143 12699
rect 22143 12665 22152 12699
rect 22100 12656 22152 12665
rect 20536 12588 20588 12640
rect 21548 12588 21600 12640
rect 22284 12656 22336 12708
rect 22744 12699 22796 12708
rect 22744 12665 22753 12699
rect 22753 12665 22787 12699
rect 22787 12665 22796 12699
rect 22744 12656 22796 12665
rect 22468 12588 22520 12640
rect 24032 12656 24084 12708
rect 25780 12631 25832 12640
rect 25780 12597 25789 12631
rect 25789 12597 25823 12631
rect 25823 12597 25832 12631
rect 25780 12588 25832 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 8392 12384 8444 12436
rect 9956 12427 10008 12436
rect 9956 12393 9965 12427
rect 9965 12393 9999 12427
rect 9999 12393 10008 12427
rect 9956 12384 10008 12393
rect 10140 12384 10192 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 13912 12427 13964 12436
rect 13912 12393 13921 12427
rect 13921 12393 13955 12427
rect 13955 12393 13964 12427
rect 13912 12384 13964 12393
rect 15200 12384 15252 12436
rect 15752 12384 15804 12436
rect 16672 12384 16724 12436
rect 19156 12384 19208 12436
rect 22100 12384 22152 12436
rect 24124 12384 24176 12436
rect 13636 12316 13688 12368
rect 15936 12316 15988 12368
rect 17316 12359 17368 12368
rect 17316 12325 17325 12359
rect 17325 12325 17359 12359
rect 17359 12325 17368 12359
rect 17316 12316 17368 12325
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 8760 12248 8812 12300
rect 10692 12248 10744 12300
rect 11888 12248 11940 12300
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 14464 12180 14516 12232
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 19064 12248 19116 12300
rect 20628 12316 20680 12368
rect 21916 12316 21968 12368
rect 23020 12316 23072 12368
rect 20168 12248 20220 12300
rect 22652 12248 22704 12300
rect 24768 12316 24820 12368
rect 15200 12112 15252 12164
rect 15844 12112 15896 12164
rect 19524 12112 19576 12164
rect 21180 12180 21232 12232
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 23020 12180 23072 12232
rect 24676 12180 24728 12232
rect 20260 12112 20312 12164
rect 22008 12112 22060 12164
rect 23756 12112 23808 12164
rect 12900 12044 12952 12096
rect 18696 12044 18748 12096
rect 20352 12044 20404 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 8484 11840 8536 11892
rect 10140 11883 10192 11892
rect 8300 11815 8352 11824
rect 8300 11781 8309 11815
rect 8309 11781 8343 11815
rect 8343 11781 8352 11815
rect 8300 11772 8352 11781
rect 8576 11704 8628 11756
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 12808 11883 12860 11892
rect 12808 11849 12817 11883
rect 12817 11849 12851 11883
rect 12851 11849 12860 11883
rect 12808 11840 12860 11849
rect 14096 11840 14148 11892
rect 14556 11840 14608 11892
rect 10048 11772 10100 11824
rect 7472 11568 7524 11620
rect 8024 11543 8076 11552
rect 8024 11509 8033 11543
rect 8033 11509 8067 11543
rect 8067 11509 8076 11543
rect 8024 11500 8076 11509
rect 9220 11500 9272 11552
rect 9588 11500 9640 11552
rect 13728 11636 13780 11688
rect 10140 11568 10192 11620
rect 12808 11568 12860 11620
rect 17040 11840 17092 11892
rect 19340 11840 19392 11892
rect 15476 11772 15528 11824
rect 15936 11772 15988 11824
rect 17316 11772 17368 11824
rect 20628 11815 20680 11824
rect 20628 11781 20637 11815
rect 20637 11781 20671 11815
rect 20671 11781 20680 11815
rect 20628 11772 20680 11781
rect 24768 11840 24820 11892
rect 24676 11772 24728 11824
rect 18052 11747 18104 11756
rect 18052 11713 18061 11747
rect 18061 11713 18095 11747
rect 18095 11713 18104 11747
rect 18052 11704 18104 11713
rect 19524 11704 19576 11756
rect 22744 11704 22796 11756
rect 23756 11747 23808 11756
rect 23756 11713 23765 11747
rect 23765 11713 23799 11747
rect 23799 11713 23808 11747
rect 23756 11704 23808 11713
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 18144 11679 18196 11688
rect 18144 11645 18153 11679
rect 18153 11645 18187 11679
rect 18187 11645 18196 11679
rect 18144 11636 18196 11645
rect 18604 11636 18656 11688
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 22008 11679 22060 11688
rect 18788 11568 18840 11620
rect 22008 11645 22017 11679
rect 22017 11645 22051 11679
rect 22051 11645 22060 11679
rect 22008 11636 22060 11645
rect 23020 11568 23072 11620
rect 24124 11568 24176 11620
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 21732 11500 21784 11552
rect 22928 11500 22980 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 8576 11296 8628 11348
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 12348 11296 12400 11348
rect 12808 11296 12860 11348
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 13912 11296 13964 11348
rect 9588 11228 9640 11280
rect 10048 11228 10100 11280
rect 10784 11228 10836 11280
rect 12256 11271 12308 11280
rect 12256 11237 12265 11271
rect 12265 11237 12299 11271
rect 12299 11237 12308 11271
rect 18144 11296 18196 11348
rect 19064 11339 19116 11348
rect 19064 11305 19073 11339
rect 19073 11305 19107 11339
rect 19107 11305 19116 11339
rect 19064 11296 19116 11305
rect 21364 11296 21416 11348
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 23020 11339 23072 11348
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 24124 11296 24176 11348
rect 25044 11296 25096 11348
rect 12256 11228 12308 11237
rect 15752 11228 15804 11280
rect 17868 11271 17920 11280
rect 17868 11237 17877 11271
rect 17877 11237 17911 11271
rect 17911 11237 17920 11271
rect 17868 11228 17920 11237
rect 20352 11228 20404 11280
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 7932 11160 7984 11212
rect 8484 11160 8536 11212
rect 9404 11160 9456 11212
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 13912 11160 13964 11212
rect 19340 11160 19392 11212
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 21180 11160 21232 11212
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 23204 11160 23256 11212
rect 25136 11160 25188 11212
rect 8576 10956 8628 11008
rect 9312 10956 9364 11008
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10876 11092 10928 11144
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 11428 11024 11480 11076
rect 12992 11024 13044 11076
rect 14648 10956 14700 11008
rect 15476 11092 15528 11144
rect 17316 11092 17368 11144
rect 15568 11024 15620 11076
rect 24216 11092 24268 11144
rect 18328 11067 18380 11076
rect 18328 11033 18337 11067
rect 18337 11033 18371 11067
rect 18371 11033 18380 11067
rect 18328 11024 18380 11033
rect 16212 10956 16264 11008
rect 17316 10956 17368 11008
rect 17500 10956 17552 11008
rect 17684 10956 17736 11008
rect 24676 10999 24728 11008
rect 24676 10965 24685 10999
rect 24685 10965 24719 10999
rect 24719 10965 24728 10999
rect 24676 10956 24728 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 7012 10752 7064 10804
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 10048 10752 10100 10804
rect 10784 10752 10836 10804
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 13636 10752 13688 10804
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 18880 10752 18932 10804
rect 21180 10752 21232 10804
rect 22284 10795 22336 10804
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 6552 10616 6604 10668
rect 7932 10616 7984 10668
rect 9956 10684 10008 10736
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 10232 10684 10284 10693
rect 10692 10684 10744 10736
rect 12440 10684 12492 10736
rect 13268 10684 13320 10736
rect 17868 10684 17920 10736
rect 19524 10684 19576 10736
rect 20904 10684 20956 10736
rect 11520 10616 11572 10668
rect 12072 10616 12124 10668
rect 12532 10659 12584 10668
rect 12532 10625 12541 10659
rect 12541 10625 12575 10659
rect 12575 10625 12584 10659
rect 12532 10616 12584 10625
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 13360 10616 13412 10668
rect 13912 10616 13964 10668
rect 14556 10616 14608 10668
rect 23480 10616 23532 10668
rect 24676 10616 24728 10668
rect 24952 10659 25004 10668
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 8576 10591 8628 10600
rect 8576 10557 8585 10591
rect 8585 10557 8619 10591
rect 8619 10557 8628 10591
rect 8576 10548 8628 10557
rect 11244 10548 11296 10600
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 9496 10480 9548 10532
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 9220 10412 9272 10464
rect 12348 10480 12400 10532
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 12624 10480 12676 10489
rect 12900 10480 12952 10532
rect 13728 10480 13780 10532
rect 14832 10548 14884 10600
rect 16396 10548 16448 10600
rect 17776 10548 17828 10600
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 16488 10480 16540 10532
rect 18788 10480 18840 10532
rect 20168 10548 20220 10600
rect 22652 10591 22704 10600
rect 22652 10557 22661 10591
rect 22661 10557 22695 10591
rect 22695 10557 22704 10591
rect 22652 10548 22704 10557
rect 9864 10412 9916 10464
rect 13360 10412 13412 10464
rect 14464 10412 14516 10464
rect 16304 10412 16356 10464
rect 17776 10412 17828 10464
rect 19248 10455 19300 10464
rect 19248 10421 19257 10455
rect 19257 10421 19291 10455
rect 19291 10421 19300 10455
rect 19248 10412 19300 10421
rect 19524 10412 19576 10464
rect 20076 10412 20128 10464
rect 21732 10412 21784 10464
rect 23204 10455 23256 10464
rect 23204 10421 23213 10455
rect 23213 10421 23247 10455
rect 23247 10421 23256 10455
rect 23204 10412 23256 10421
rect 24860 10412 24912 10464
rect 25136 10412 25188 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 9312 10208 9364 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 11520 10251 11572 10260
rect 11520 10217 11529 10251
rect 11529 10217 11563 10251
rect 11563 10217 11572 10251
rect 11520 10208 11572 10217
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 17224 10208 17276 10260
rect 9956 10140 10008 10192
rect 6644 10072 6696 10124
rect 7104 10072 7156 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 9864 10072 9916 10124
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 11428 10140 11480 10192
rect 11152 10072 11204 10124
rect 12256 10140 12308 10192
rect 12348 10140 12400 10192
rect 13544 10183 13596 10192
rect 13544 10149 13553 10183
rect 13553 10149 13587 10183
rect 13587 10149 13596 10183
rect 13544 10140 13596 10149
rect 13636 10183 13688 10192
rect 13636 10149 13645 10183
rect 13645 10149 13679 10183
rect 13679 10149 13688 10183
rect 13636 10140 13688 10149
rect 15936 10140 15988 10192
rect 12532 10072 12584 10124
rect 15568 10072 15620 10124
rect 12440 10004 12492 10056
rect 12808 10004 12860 10056
rect 17316 10140 17368 10192
rect 18052 10208 18104 10260
rect 18972 10208 19024 10260
rect 23204 10140 23256 10192
rect 23480 10183 23532 10192
rect 23480 10149 23489 10183
rect 23489 10149 23523 10183
rect 23523 10149 23532 10183
rect 23480 10140 23532 10149
rect 24216 10140 24268 10192
rect 19064 10115 19116 10124
rect 19064 10081 19073 10115
rect 19073 10081 19107 10115
rect 19107 10081 19116 10115
rect 19064 10072 19116 10081
rect 19248 10115 19300 10124
rect 19248 10081 19257 10115
rect 19257 10081 19291 10115
rect 19291 10081 19300 10115
rect 19248 10072 19300 10081
rect 20444 10072 20496 10124
rect 10416 9936 10468 9988
rect 14096 9979 14148 9988
rect 14096 9945 14105 9979
rect 14105 9945 14139 9979
rect 14139 9945 14148 9979
rect 14096 9936 14148 9945
rect 10140 9868 10192 9920
rect 12900 9868 12952 9920
rect 14280 9868 14332 9920
rect 14832 9868 14884 9920
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 18328 10004 18380 10056
rect 18788 10004 18840 10056
rect 21364 10072 21416 10124
rect 22836 10047 22888 10056
rect 22836 10013 22845 10047
rect 22845 10013 22879 10047
rect 22879 10013 22888 10047
rect 22836 10004 22888 10013
rect 18696 9936 18748 9988
rect 20628 9979 20680 9988
rect 20628 9945 20637 9979
rect 20637 9945 20671 9979
rect 20671 9945 20680 9979
rect 20628 9936 20680 9945
rect 20996 9979 21048 9988
rect 20996 9945 21005 9979
rect 21005 9945 21039 9979
rect 21039 9945 21048 9979
rect 20996 9936 21048 9945
rect 24768 10004 24820 10056
rect 25228 10004 25280 10056
rect 23572 9936 23624 9988
rect 24124 9936 24176 9988
rect 17040 9868 17092 9877
rect 20076 9868 20128 9920
rect 20168 9868 20220 9920
rect 21364 9868 21416 9920
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 23296 9868 23348 9920
rect 24216 9868 24268 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 7104 9707 7156 9716
rect 7104 9673 7113 9707
rect 7113 9673 7147 9707
rect 7147 9673 7156 9707
rect 7104 9664 7156 9673
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 9220 9664 9272 9716
rect 9864 9707 9916 9716
rect 9864 9673 9873 9707
rect 9873 9673 9907 9707
rect 9907 9673 9916 9707
rect 9864 9664 9916 9673
rect 9956 9664 10008 9716
rect 10232 9664 10284 9716
rect 12256 9707 12308 9716
rect 12256 9673 12265 9707
rect 12265 9673 12299 9707
rect 12299 9673 12308 9707
rect 12256 9664 12308 9673
rect 13636 9707 13688 9716
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 14648 9664 14700 9716
rect 15660 9664 15712 9716
rect 15936 9664 15988 9716
rect 17224 9707 17276 9716
rect 17224 9673 17233 9707
rect 17233 9673 17267 9707
rect 17267 9673 17276 9707
rect 17224 9664 17276 9673
rect 19064 9707 19116 9716
rect 19064 9673 19073 9707
rect 19073 9673 19107 9707
rect 19107 9673 19116 9707
rect 19064 9664 19116 9673
rect 23572 9664 23624 9716
rect 24216 9707 24268 9716
rect 24216 9673 24225 9707
rect 24225 9673 24259 9707
rect 24259 9673 24268 9707
rect 24216 9664 24268 9673
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 11980 9596 12032 9648
rect 13544 9596 13596 9648
rect 22192 9596 22244 9648
rect 9312 9528 9364 9580
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 11060 9528 11112 9580
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 14096 9528 14148 9580
rect 17040 9528 17092 9580
rect 18236 9528 18288 9580
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 19524 9528 19576 9580
rect 22284 9528 22336 9580
rect 24124 9528 24176 9580
rect 24952 9571 25004 9580
rect 24952 9537 24961 9571
rect 24961 9537 24995 9571
rect 24995 9537 25004 9571
rect 24952 9528 25004 9537
rect 8116 9460 8168 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 8760 9392 8812 9444
rect 9220 9460 9272 9512
rect 10232 9460 10284 9512
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 6092 9324 6144 9376
rect 8024 9324 8076 9376
rect 8668 9324 8720 9376
rect 10784 9392 10836 9444
rect 12256 9392 12308 9444
rect 14188 9392 14240 9444
rect 11612 9324 11664 9376
rect 15660 9324 15712 9376
rect 16212 9392 16264 9444
rect 17960 9324 18012 9376
rect 19524 9392 19576 9444
rect 20996 9435 21048 9444
rect 20996 9401 21005 9435
rect 21005 9401 21039 9435
rect 21039 9401 21048 9435
rect 20996 9392 21048 9401
rect 21456 9392 21508 9444
rect 22928 9392 22980 9444
rect 23572 9392 23624 9444
rect 21364 9367 21416 9376
rect 21364 9333 21373 9367
rect 21373 9333 21407 9367
rect 21407 9333 21416 9367
rect 21364 9324 21416 9333
rect 23204 9324 23256 9376
rect 24676 9392 24728 9444
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 6092 9120 6144 9172
rect 10140 9120 10192 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 15476 9120 15528 9172
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 16396 9120 16448 9172
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 8576 9052 8628 9104
rect 9772 9095 9824 9104
rect 9772 9061 9781 9095
rect 9781 9061 9815 9095
rect 9815 9061 9824 9095
rect 9772 9052 9824 9061
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 12624 9052 12676 9104
rect 14096 9095 14148 9104
rect 14096 9061 14105 9095
rect 14105 9061 14139 9095
rect 14139 9061 14148 9095
rect 14096 9052 14148 9061
rect 17224 9052 17276 9104
rect 17776 9052 17828 9104
rect 18972 9052 19024 9104
rect 5448 9027 5500 9036
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 7380 8984 7432 9036
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 11888 8984 11940 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 16304 8984 16356 9036
rect 19984 9052 20036 9104
rect 20444 9120 20496 9172
rect 20628 9163 20680 9172
rect 20628 9129 20637 9163
rect 20637 9129 20671 9163
rect 20671 9129 20680 9163
rect 20628 9120 20680 9129
rect 24768 9120 24820 9172
rect 23572 9052 23624 9104
rect 19708 8984 19760 9036
rect 20812 8984 20864 9036
rect 21272 8984 21324 9036
rect 21916 9027 21968 9036
rect 21916 8993 21925 9027
rect 21925 8993 21959 9027
rect 21959 8993 21968 9027
rect 21916 8984 21968 8993
rect 6736 8916 6788 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 8760 8916 8812 8968
rect 13176 8916 13228 8968
rect 17684 8916 17736 8968
rect 17776 8916 17828 8968
rect 21640 8916 21692 8968
rect 22008 8916 22060 8968
rect 24032 8916 24084 8968
rect 24216 8916 24268 8968
rect 8944 8848 8996 8900
rect 10324 8891 10376 8900
rect 10324 8857 10333 8891
rect 10333 8857 10367 8891
rect 10367 8857 10376 8891
rect 10324 8848 10376 8857
rect 10784 8848 10836 8900
rect 11152 8848 11204 8900
rect 14188 8848 14240 8900
rect 19524 8848 19576 8900
rect 8116 8780 8168 8832
rect 11060 8780 11112 8832
rect 16580 8780 16632 8832
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 24860 8780 24912 8832
rect 25228 8780 25280 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 9772 8576 9824 8628
rect 12624 8576 12676 8628
rect 13544 8576 13596 8628
rect 15292 8576 15344 8628
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 20904 8576 20956 8628
rect 23296 8576 23348 8628
rect 23848 8576 23900 8628
rect 24032 8576 24084 8628
rect 9588 8508 9640 8560
rect 13728 8508 13780 8560
rect 21364 8508 21416 8560
rect 8576 8440 8628 8492
rect 10324 8440 10376 8492
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 16580 8440 16632 8492
rect 20628 8440 20680 8492
rect 22284 8483 22336 8492
rect 6000 8372 6052 8424
rect 6736 8372 6788 8424
rect 7288 8372 7340 8424
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 15016 8372 15068 8424
rect 15660 8372 15712 8424
rect 5448 8304 5500 8356
rect 6092 8304 6144 8356
rect 8208 8304 8260 8356
rect 9220 8304 9272 8356
rect 10968 8347 11020 8356
rect 10968 8313 10977 8347
rect 10977 8313 11011 8347
rect 11011 8313 11020 8347
rect 10968 8304 11020 8313
rect 11152 8304 11204 8356
rect 13544 8347 13596 8356
rect 13544 8313 13553 8347
rect 13553 8313 13587 8347
rect 13587 8313 13596 8347
rect 14096 8347 14148 8356
rect 13544 8304 13596 8313
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 16396 8347 16448 8356
rect 14096 8304 14148 8313
rect 6368 8236 6420 8288
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 6828 8236 6880 8288
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 9864 8236 9916 8288
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 13452 8236 13504 8288
rect 15016 8236 15068 8288
rect 16120 8236 16172 8288
rect 16396 8313 16405 8347
rect 16405 8313 16439 8347
rect 16439 8313 16448 8347
rect 16396 8304 16448 8313
rect 18236 8304 18288 8356
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 21272 8415 21324 8424
rect 21272 8381 21281 8415
rect 21281 8381 21315 8415
rect 21315 8381 21324 8415
rect 21272 8372 21324 8381
rect 19984 8304 20036 8356
rect 21916 8372 21968 8424
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 23388 8440 23440 8492
rect 22560 8372 22612 8424
rect 25044 8372 25096 8424
rect 23756 8347 23808 8356
rect 23756 8313 23765 8347
rect 23765 8313 23799 8347
rect 23799 8313 23808 8347
rect 23756 8304 23808 8313
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 17684 8279 17736 8288
rect 17684 8245 17693 8279
rect 17693 8245 17727 8279
rect 17727 8245 17736 8279
rect 17684 8236 17736 8245
rect 18420 8236 18472 8288
rect 20628 8279 20680 8288
rect 20628 8245 20637 8279
rect 20637 8245 20671 8279
rect 20671 8245 20680 8279
rect 20628 8236 20680 8245
rect 21732 8236 21784 8288
rect 22468 8236 22520 8288
rect 23572 8236 23624 8288
rect 25688 8279 25740 8288
rect 25688 8245 25697 8279
rect 25697 8245 25731 8279
rect 25731 8245 25740 8279
rect 25688 8236 25740 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8576 8032 8628 8084
rect 9772 8075 9824 8084
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 11336 8032 11388 8084
rect 11428 8032 11480 8084
rect 13176 8075 13228 8084
rect 7748 8007 7800 8016
rect 7748 7973 7757 8007
rect 7757 7973 7791 8007
rect 7791 7973 7800 8007
rect 7748 7964 7800 7973
rect 7840 7964 7892 8016
rect 5540 7939 5592 7948
rect 5540 7905 5549 7939
rect 5549 7905 5583 7939
rect 5583 7905 5592 7939
rect 5540 7896 5592 7905
rect 8484 7964 8536 8016
rect 11612 8007 11664 8016
rect 11612 7973 11621 8007
rect 11621 7973 11655 8007
rect 11655 7973 11664 8007
rect 11612 7964 11664 7973
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 14280 8032 14332 8084
rect 13636 7964 13688 8016
rect 14096 8007 14148 8016
rect 14096 7973 14105 8007
rect 14105 7973 14139 8007
rect 14139 7973 14148 8007
rect 14096 7964 14148 7973
rect 9496 7896 9548 7948
rect 10140 7896 10192 7948
rect 16396 8032 16448 8084
rect 17684 8032 17736 8084
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 17132 8007 17184 8016
rect 17132 7973 17141 8007
rect 17141 7973 17175 8007
rect 17175 7973 17184 8007
rect 17132 7964 17184 7973
rect 21916 8032 21968 8084
rect 23756 8032 23808 8084
rect 7012 7828 7064 7880
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 8116 7760 8168 7812
rect 15752 7896 15804 7948
rect 16028 7896 16080 7948
rect 17960 7896 18012 7948
rect 20628 7964 20680 8016
rect 21272 7964 21324 8016
rect 23296 8007 23348 8016
rect 23296 7973 23305 8007
rect 23305 7973 23339 8007
rect 23339 7973 23348 8007
rect 23296 7964 23348 7973
rect 24216 8007 24268 8016
rect 24216 7973 24225 8007
rect 24225 7973 24259 8007
rect 24259 7973 24268 8007
rect 24216 7964 24268 7973
rect 24676 8007 24728 8016
rect 24676 7973 24685 8007
rect 24685 7973 24719 8007
rect 24719 7973 24728 8007
rect 24676 7964 24728 7973
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 13728 7828 13780 7880
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 17316 7871 17368 7880
rect 6920 7692 6972 7744
rect 7564 7692 7616 7744
rect 11888 7760 11940 7812
rect 14832 7760 14884 7812
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 20996 7896 21048 7948
rect 21732 7939 21784 7948
rect 21732 7905 21741 7939
rect 21741 7905 21775 7939
rect 21775 7905 21784 7939
rect 21732 7896 21784 7905
rect 22468 7896 22520 7948
rect 24124 7896 24176 7948
rect 25228 7939 25280 7948
rect 25228 7905 25237 7939
rect 25237 7905 25271 7939
rect 25271 7905 25280 7939
rect 25228 7896 25280 7905
rect 22928 7828 22980 7880
rect 23020 7828 23072 7880
rect 9680 7692 9732 7744
rect 9956 7692 10008 7744
rect 11428 7692 11480 7744
rect 14740 7692 14792 7744
rect 16396 7735 16448 7744
rect 16396 7701 16405 7735
rect 16405 7701 16439 7735
rect 16439 7701 16448 7735
rect 16396 7692 16448 7701
rect 20996 7760 21048 7812
rect 21640 7692 21692 7744
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 6460 7488 6512 7540
rect 7012 7488 7064 7540
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 10968 7488 11020 7540
rect 11612 7488 11664 7540
rect 13636 7488 13688 7540
rect 13728 7488 13780 7540
rect 11152 7420 11204 7472
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 10784 7352 10836 7404
rect 11796 7352 11848 7404
rect 8116 7259 8168 7268
rect 8116 7225 8125 7259
rect 8125 7225 8159 7259
rect 8159 7225 8168 7259
rect 8116 7216 8168 7225
rect 12164 7216 12216 7268
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 9496 7148 9548 7200
rect 14188 7216 14240 7268
rect 14740 7284 14792 7336
rect 16028 7488 16080 7540
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 15752 7420 15804 7472
rect 17960 7488 18012 7540
rect 18972 7488 19024 7540
rect 23296 7488 23348 7540
rect 25228 7531 25280 7540
rect 25228 7497 25237 7531
rect 25237 7497 25271 7531
rect 25271 7497 25280 7531
rect 25228 7488 25280 7497
rect 25872 7531 25924 7540
rect 25872 7497 25881 7531
rect 25881 7497 25915 7531
rect 25915 7497 25924 7531
rect 25872 7488 25924 7497
rect 19064 7463 19116 7472
rect 19064 7429 19073 7463
rect 19073 7429 19107 7463
rect 19107 7429 19116 7463
rect 19984 7463 20036 7472
rect 19064 7420 19116 7429
rect 19984 7429 19993 7463
rect 19993 7429 20027 7463
rect 20027 7429 20036 7463
rect 19984 7420 20036 7429
rect 20628 7463 20680 7472
rect 20628 7429 20637 7463
rect 20637 7429 20671 7463
rect 20671 7429 20680 7463
rect 20628 7420 20680 7429
rect 21732 7420 21784 7472
rect 16948 7352 17000 7404
rect 18696 7352 18748 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 20536 7327 20588 7336
rect 12900 7148 12952 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 16396 7216 16448 7268
rect 17408 7216 17460 7268
rect 20536 7293 20545 7327
rect 20545 7293 20579 7327
rect 20579 7293 20588 7327
rect 20536 7284 20588 7293
rect 21364 7352 21416 7404
rect 24216 7352 24268 7404
rect 20076 7216 20128 7268
rect 18236 7148 18288 7200
rect 19064 7148 19116 7200
rect 21824 7216 21876 7268
rect 25872 7284 25924 7336
rect 24032 7259 24084 7268
rect 24032 7225 24041 7259
rect 24041 7225 24075 7259
rect 24075 7225 24084 7259
rect 24032 7216 24084 7225
rect 24676 7216 24728 7268
rect 25780 7216 25832 7268
rect 20996 7191 21048 7200
rect 20996 7157 21005 7191
rect 21005 7157 21039 7191
rect 21039 7157 21048 7191
rect 20996 7148 21048 7157
rect 22560 7191 22612 7200
rect 22560 7157 22569 7191
rect 22569 7157 22603 7191
rect 22603 7157 22612 7191
rect 22560 7148 22612 7157
rect 22928 7191 22980 7200
rect 22928 7157 22937 7191
rect 22937 7157 22971 7191
rect 22971 7157 22980 7191
rect 22928 7148 22980 7157
rect 25320 7148 25372 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 7748 6944 7800 6996
rect 6552 6876 6604 6928
rect 8116 6944 8168 6996
rect 8300 6944 8352 6996
rect 12256 6944 12308 6996
rect 12900 6987 12952 6996
rect 8392 6876 8444 6928
rect 9404 6808 9456 6860
rect 10692 6876 10744 6928
rect 12900 6953 12909 6987
rect 12909 6953 12943 6987
rect 12943 6953 12952 6987
rect 12900 6944 12952 6953
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 16120 6944 16172 6996
rect 18696 6987 18748 6996
rect 14740 6876 14792 6928
rect 17224 6919 17276 6928
rect 17224 6885 17233 6919
rect 17233 6885 17267 6919
rect 17267 6885 17276 6919
rect 17224 6876 17276 6885
rect 14004 6851 14056 6860
rect 14004 6817 14013 6851
rect 14013 6817 14047 6851
rect 14047 6817 14056 6851
rect 14004 6808 14056 6817
rect 18696 6953 18705 6987
rect 18705 6953 18739 6987
rect 18739 6953 18748 6987
rect 18696 6944 18748 6953
rect 20536 6987 20588 6996
rect 20536 6953 20545 6987
rect 20545 6953 20579 6987
rect 20579 6953 20588 6987
rect 20536 6944 20588 6953
rect 23572 6987 23624 6996
rect 23572 6953 23581 6987
rect 23581 6953 23615 6987
rect 23615 6953 23624 6987
rect 23572 6944 23624 6953
rect 18972 6876 19024 6928
rect 19800 6808 19852 6860
rect 20260 6808 20312 6860
rect 20812 6808 20864 6860
rect 21272 6808 21324 6860
rect 21732 6851 21784 6860
rect 21732 6817 21741 6851
rect 21741 6817 21775 6851
rect 21775 6817 21784 6851
rect 21732 6808 21784 6817
rect 21824 6808 21876 6860
rect 22192 6808 22244 6860
rect 25044 6808 25096 6860
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 6460 6740 6512 6792
rect 7564 6740 7616 6792
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 10508 6783 10560 6792
rect 7748 6604 7800 6656
rect 8852 6604 8904 6656
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 10140 6672 10192 6724
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11796 6740 11848 6792
rect 12532 6740 12584 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 17408 6783 17460 6792
rect 14832 6672 14884 6724
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 17500 6740 17552 6792
rect 17776 6672 17828 6724
rect 19432 6740 19484 6792
rect 23296 6740 23348 6792
rect 25412 6672 25464 6724
rect 11520 6604 11572 6656
rect 11612 6604 11664 6656
rect 15936 6604 15988 6656
rect 16396 6604 16448 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 18052 6604 18104 6656
rect 19524 6604 19576 6656
rect 22008 6604 22060 6656
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 24216 6604 24268 6656
rect 24768 6604 24820 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 7104 6400 7156 6452
rect 7840 6400 7892 6452
rect 9772 6400 9824 6452
rect 10692 6400 10744 6452
rect 12256 6400 12308 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14096 6400 14148 6452
rect 17500 6400 17552 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18972 6443 19024 6452
rect 18972 6409 18981 6443
rect 18981 6409 19015 6443
rect 19015 6409 19024 6443
rect 18972 6400 19024 6409
rect 25044 6443 25096 6452
rect 25044 6409 25053 6443
rect 25053 6409 25087 6443
rect 25087 6409 25096 6443
rect 25044 6400 25096 6409
rect 4712 6332 4764 6384
rect 9864 6332 9916 6384
rect 10508 6375 10560 6384
rect 5172 6264 5224 6316
rect 6000 6264 6052 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7380 6264 7432 6316
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 8116 6264 8168 6316
rect 8392 6264 8444 6316
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 15844 6332 15896 6384
rect 6920 6128 6972 6180
rect 8668 6196 8720 6248
rect 7656 6128 7708 6180
rect 9588 6196 9640 6248
rect 11888 6264 11940 6316
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 14464 6264 14516 6316
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 20904 6332 20956 6384
rect 15568 6196 15620 6248
rect 17224 6196 17276 6248
rect 9404 6171 9456 6180
rect 9404 6137 9413 6171
rect 9413 6137 9447 6171
rect 9447 6137 9456 6171
rect 9404 6128 9456 6137
rect 9680 6128 9732 6180
rect 15660 6171 15712 6180
rect 15660 6137 15669 6171
rect 15669 6137 15703 6171
rect 15703 6137 15712 6171
rect 15660 6128 15712 6137
rect 19156 6264 19208 6316
rect 19800 6239 19852 6248
rect 6276 6103 6328 6112
rect 6276 6069 6285 6103
rect 6285 6069 6319 6103
rect 6319 6069 6328 6103
rect 6276 6060 6328 6069
rect 8576 6060 8628 6112
rect 11244 6060 11296 6112
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 19800 6205 19809 6239
rect 19809 6205 19843 6239
rect 19843 6205 19852 6239
rect 19800 6196 19852 6205
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 21732 6264 21784 6316
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 24676 6332 24728 6384
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22100 6196 22152 6205
rect 21180 6128 21232 6180
rect 22376 6196 22428 6248
rect 23756 6171 23808 6180
rect 23756 6137 23765 6171
rect 23765 6137 23799 6171
rect 23799 6137 23808 6171
rect 23756 6128 23808 6137
rect 24216 6128 24268 6180
rect 18696 6060 18748 6112
rect 19340 6103 19392 6112
rect 19340 6069 19349 6103
rect 19349 6069 19383 6103
rect 19383 6069 19392 6103
rect 19340 6060 19392 6069
rect 19432 6060 19484 6112
rect 23572 6060 23624 6112
rect 27252 6128 27304 6180
rect 25044 6060 25096 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 10140 5856 10192 5908
rect 12440 5856 12492 5908
rect 13084 5856 13136 5908
rect 16028 5856 16080 5908
rect 16580 5856 16632 5908
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 5264 5788 5316 5840
rect 7656 5788 7708 5840
rect 8392 5788 8444 5840
rect 8944 5788 8996 5840
rect 9128 5788 9180 5840
rect 10048 5788 10100 5840
rect 11888 5831 11940 5840
rect 11888 5797 11897 5831
rect 11897 5797 11931 5831
rect 11931 5797 11940 5831
rect 11888 5788 11940 5797
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 6644 5720 6696 5772
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 11152 5720 11204 5772
rect 14004 5720 14056 5772
rect 14740 5788 14792 5840
rect 16948 5856 17000 5908
rect 17316 5856 17368 5908
rect 19432 5856 19484 5908
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 20076 5856 20128 5908
rect 23296 5899 23348 5908
rect 23296 5865 23305 5899
rect 23305 5865 23339 5899
rect 23339 5865 23348 5899
rect 23296 5856 23348 5865
rect 24032 5899 24084 5908
rect 24032 5865 24041 5899
rect 24041 5865 24075 5899
rect 24075 5865 24084 5899
rect 24032 5856 24084 5865
rect 17040 5788 17092 5840
rect 17408 5788 17460 5840
rect 18604 5788 18656 5840
rect 19248 5788 19300 5840
rect 21456 5788 21508 5840
rect 23848 5788 23900 5840
rect 24124 5788 24176 5840
rect 15384 5720 15436 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 21364 5763 21416 5772
rect 21364 5729 21373 5763
rect 21373 5729 21407 5763
rect 21407 5729 21416 5763
rect 21364 5720 21416 5729
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 24216 5763 24268 5772
rect 24216 5729 24225 5763
rect 24225 5729 24259 5763
rect 24259 5729 24268 5763
rect 24216 5720 24268 5729
rect 25780 5720 25832 5772
rect 7840 5652 7892 5704
rect 6736 5584 6788 5636
rect 7564 5584 7616 5636
rect 10140 5652 10192 5704
rect 10876 5652 10928 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 13544 5652 13596 5704
rect 14188 5695 14240 5704
rect 14188 5661 14197 5695
rect 14197 5661 14231 5695
rect 14231 5661 14240 5695
rect 14188 5652 14240 5661
rect 6276 5516 6328 5568
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 7380 5516 7432 5568
rect 7656 5516 7708 5568
rect 9128 5559 9180 5568
rect 9128 5525 9137 5559
rect 9137 5525 9171 5559
rect 9171 5525 9180 5559
rect 9128 5516 9180 5525
rect 12532 5584 12584 5636
rect 15292 5584 15344 5636
rect 16672 5584 16724 5636
rect 11428 5559 11480 5568
rect 11428 5525 11437 5559
rect 11437 5525 11471 5559
rect 11471 5525 11480 5559
rect 11428 5516 11480 5525
rect 15660 5516 15712 5568
rect 17960 5559 18012 5568
rect 17960 5525 17969 5559
rect 17969 5525 18003 5559
rect 18003 5525 18012 5559
rect 19616 5652 19668 5704
rect 23664 5652 23716 5704
rect 23756 5652 23808 5704
rect 17960 5516 18012 5525
rect 21456 5516 21508 5568
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 22744 5516 22796 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 6460 5312 6512 5364
rect 6552 5312 6604 5364
rect 7196 5312 7248 5364
rect 8116 5312 8168 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 10048 5355 10100 5364
rect 10048 5321 10057 5355
rect 10057 5321 10091 5355
rect 10091 5321 10100 5355
rect 10048 5312 10100 5321
rect 15384 5312 15436 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 5264 5287 5316 5296
rect 5264 5253 5273 5287
rect 5273 5253 5307 5287
rect 5307 5253 5316 5287
rect 5264 5244 5316 5253
rect 6368 5244 6420 5296
rect 7472 5244 7524 5296
rect 9956 5244 10008 5296
rect 6460 5176 6512 5228
rect 9496 5176 9548 5228
rect 14740 5244 14792 5296
rect 15936 5244 15988 5296
rect 18788 5244 18840 5296
rect 12532 5176 12584 5228
rect 19064 5312 19116 5364
rect 19984 5312 20036 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 22468 5312 22520 5364
rect 20444 5287 20496 5296
rect 20444 5253 20453 5287
rect 20453 5253 20487 5287
rect 20487 5253 20496 5287
rect 20444 5244 20496 5253
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 24216 5312 24268 5364
rect 23848 5244 23900 5296
rect 26516 5244 26568 5296
rect 6184 5108 6236 5160
rect 7104 5108 7156 5160
rect 8300 5108 8352 5160
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 7472 5040 7524 5092
rect 7656 5083 7708 5092
rect 7656 5049 7665 5083
rect 7665 5049 7699 5083
rect 7699 5049 7708 5083
rect 7656 5040 7708 5049
rect 8116 5040 8168 5092
rect 8668 5040 8720 5092
rect 1400 4972 1452 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 5080 4972 5132 5024
rect 5448 4972 5500 5024
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 9220 4972 9272 5024
rect 12348 5040 12400 5092
rect 12532 5083 12584 5092
rect 12532 5049 12541 5083
rect 12541 5049 12575 5083
rect 12575 5049 12584 5083
rect 12532 5040 12584 5049
rect 13176 5083 13228 5092
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 13176 5049 13185 5083
rect 13185 5049 13219 5083
rect 13219 5049 13228 5083
rect 13176 5040 13228 5049
rect 12716 4972 12768 5024
rect 13084 4972 13136 5024
rect 14740 5108 14792 5160
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 16580 5108 16632 5160
rect 19616 5108 19668 5160
rect 19984 5108 20036 5160
rect 15476 5040 15528 5092
rect 17132 5083 17184 5092
rect 17132 5049 17141 5083
rect 17141 5049 17175 5083
rect 17175 5049 17184 5083
rect 17132 5040 17184 5049
rect 19340 5040 19392 5092
rect 21548 5108 21600 5160
rect 22008 5151 22060 5160
rect 22008 5117 22017 5151
rect 22017 5117 22051 5151
rect 22051 5117 22060 5151
rect 22008 5108 22060 5117
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22284 5151 22336 5160
rect 22100 5108 22152 5117
rect 22284 5117 22293 5151
rect 22293 5117 22327 5151
rect 22327 5117 22336 5151
rect 22284 5108 22336 5117
rect 23664 5151 23716 5160
rect 23664 5117 23673 5151
rect 23673 5117 23707 5151
rect 23707 5117 23716 5151
rect 23664 5108 23716 5117
rect 23756 5151 23808 5160
rect 23756 5117 23765 5151
rect 23765 5117 23799 5151
rect 23799 5117 23808 5151
rect 23756 5108 23808 5117
rect 23480 5083 23532 5092
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 20812 5015 20864 5024
rect 20812 4981 20821 5015
rect 20821 4981 20855 5015
rect 20855 4981 20864 5015
rect 20812 4972 20864 4981
rect 23480 5049 23489 5083
rect 23489 5049 23523 5083
rect 23523 5049 23532 5083
rect 24032 5108 24084 5160
rect 23480 5040 23532 5049
rect 24860 5040 24912 5092
rect 25780 5083 25832 5092
rect 25780 5049 25789 5083
rect 25789 5049 25823 5083
rect 25823 5049 25832 5083
rect 25780 5040 25832 5049
rect 23664 4972 23716 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 7564 4768 7616 4820
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 8484 4768 8536 4820
rect 9772 4768 9824 4820
rect 11244 4768 11296 4820
rect 12532 4768 12584 4820
rect 14740 4768 14792 4820
rect 15752 4768 15804 4820
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 19524 4811 19576 4820
rect 19524 4777 19533 4811
rect 19533 4777 19567 4811
rect 19567 4777 19576 4811
rect 19524 4768 19576 4777
rect 19984 4811 20036 4820
rect 19984 4777 19993 4811
rect 19993 4777 20027 4811
rect 20027 4777 20036 4811
rect 19984 4768 20036 4777
rect 20444 4811 20496 4820
rect 20444 4777 20453 4811
rect 20453 4777 20487 4811
rect 20487 4777 20496 4811
rect 20444 4768 20496 4777
rect 22100 4768 22152 4820
rect 3608 4632 3660 4684
rect 5540 4632 5592 4684
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6828 4632 6880 4684
rect 6920 4632 6972 4684
rect 7104 4632 7156 4684
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 8208 4675 8260 4684
rect 8208 4641 8217 4675
rect 8217 4641 8251 4675
rect 8251 4641 8260 4675
rect 8208 4632 8260 4641
rect 8300 4632 8352 4684
rect 8392 4564 8444 4616
rect 7564 4496 7616 4548
rect 12256 4700 12308 4752
rect 13268 4743 13320 4752
rect 13268 4709 13277 4743
rect 13277 4709 13311 4743
rect 13311 4709 13320 4743
rect 13268 4700 13320 4709
rect 18512 4743 18564 4752
rect 18512 4709 18521 4743
rect 18521 4709 18555 4743
rect 18555 4709 18564 4743
rect 18512 4700 18564 4709
rect 9128 4564 9180 4616
rect 9312 4564 9364 4616
rect 11520 4632 11572 4684
rect 16764 4632 16816 4684
rect 19156 4675 19208 4684
rect 19156 4641 19165 4675
rect 19165 4641 19199 4675
rect 19199 4641 19208 4675
rect 19156 4632 19208 4641
rect 20812 4632 20864 4684
rect 22560 4632 22612 4684
rect 23480 4632 23532 4684
rect 23756 4675 23808 4684
rect 23756 4641 23765 4675
rect 23765 4641 23799 4675
rect 23799 4641 23808 4675
rect 24124 4700 24176 4752
rect 23756 4632 23808 4641
rect 24952 4632 25004 4684
rect 11244 4564 11296 4616
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13544 4607 13596 4616
rect 10876 4496 10928 4548
rect 13084 4496 13136 4548
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 15476 4564 15528 4616
rect 22284 4564 22336 4616
rect 24216 4564 24268 4616
rect 13452 4496 13504 4548
rect 18144 4539 18196 4548
rect 18144 4505 18153 4539
rect 18153 4505 18187 4539
rect 18187 4505 18196 4539
rect 18144 4496 18196 4505
rect 22744 4496 22796 4548
rect 8208 4428 8260 4480
rect 9128 4428 9180 4480
rect 11336 4428 11388 4480
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 16580 4471 16632 4480
rect 16580 4437 16589 4471
rect 16589 4437 16623 4471
rect 16623 4437 16632 4471
rect 16580 4428 16632 4437
rect 17960 4428 18012 4480
rect 18236 4428 18288 4480
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 3608 4267 3660 4276
rect 3608 4233 3617 4267
rect 3617 4233 3651 4267
rect 3651 4233 3660 4267
rect 3608 4224 3660 4233
rect 3976 4267 4028 4276
rect 3976 4233 3985 4267
rect 3985 4233 4019 4267
rect 4019 4233 4028 4267
rect 3976 4224 4028 4233
rect 5540 4267 5592 4276
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 8944 4224 8996 4276
rect 9128 4224 9180 4276
rect 10968 4224 11020 4276
rect 11704 4224 11756 4276
rect 12256 4224 12308 4276
rect 16212 4267 16264 4276
rect 5356 4156 5408 4208
rect 6000 4156 6052 4208
rect 6828 4156 6880 4208
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 5172 3884 5224 3936
rect 7012 4020 7064 4072
rect 8668 4156 8720 4208
rect 10048 4156 10100 4208
rect 14188 4156 14240 4208
rect 16212 4233 16221 4267
rect 16221 4233 16255 4267
rect 16255 4233 16264 4267
rect 16212 4224 16264 4233
rect 19156 4267 19208 4276
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 20812 4224 20864 4276
rect 21180 4224 21232 4276
rect 9128 4088 9180 4140
rect 8392 4020 8444 4072
rect 7104 3952 7156 4004
rect 8668 3952 8720 4004
rect 11244 4088 11296 4140
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 10876 3995 10928 4004
rect 6828 3884 6880 3936
rect 7656 3884 7708 3936
rect 10876 3961 10885 3995
rect 10885 3961 10919 3995
rect 10919 3961 10928 3995
rect 10876 3952 10928 3961
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 11336 3952 11388 4004
rect 11520 3995 11572 4004
rect 11520 3961 11529 3995
rect 11529 3961 11563 3995
rect 11563 3961 11572 3995
rect 11520 3952 11572 3961
rect 12532 3995 12584 4004
rect 12532 3961 12541 3995
rect 12541 3961 12575 3995
rect 12575 3961 12584 3995
rect 12532 3952 12584 3961
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 13268 3952 13320 4004
rect 14464 4156 14516 4208
rect 16580 4156 16632 4208
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 16764 4088 16816 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 20444 4156 20496 4208
rect 20076 4020 20128 4072
rect 20260 4020 20312 4072
rect 21456 4156 21508 4208
rect 25412 4267 25464 4276
rect 22560 4199 22612 4208
rect 22560 4165 22569 4199
rect 22569 4165 22603 4199
rect 22603 4165 22612 4199
rect 22560 4156 22612 4165
rect 25412 4233 25421 4267
rect 25421 4233 25455 4267
rect 25455 4233 25464 4267
rect 25412 4224 25464 4233
rect 23664 4156 23716 4208
rect 22928 4088 22980 4140
rect 21732 4063 21784 4072
rect 21732 4029 21741 4063
rect 21741 4029 21775 4063
rect 21775 4029 21784 4063
rect 21732 4020 21784 4029
rect 21824 4020 21876 4072
rect 16212 3952 16264 4004
rect 12164 3884 12216 3893
rect 13820 3884 13872 3936
rect 15752 3884 15804 3936
rect 17684 3952 17736 4004
rect 18512 3952 18564 4004
rect 22744 3952 22796 4004
rect 20076 3884 20128 3936
rect 21824 3884 21876 3936
rect 23020 3884 23072 3936
rect 24952 3884 25004 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 7012 3680 7064 3732
rect 7840 3723 7892 3732
rect 7840 3689 7849 3723
rect 7849 3689 7883 3723
rect 7883 3689 7892 3723
rect 7840 3680 7892 3689
rect 9772 3680 9824 3732
rect 11244 3680 11296 3732
rect 13544 3680 13596 3732
rect 15476 3723 15528 3732
rect 15476 3689 15485 3723
rect 15485 3689 15519 3723
rect 15519 3689 15528 3723
rect 15476 3680 15528 3689
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 4620 3544 4672 3596
rect 5356 3544 5408 3596
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 9404 3612 9456 3664
rect 10048 3612 10100 3664
rect 11704 3612 11756 3664
rect 13728 3612 13780 3664
rect 13820 3655 13872 3664
rect 13820 3621 13829 3655
rect 13829 3621 13863 3655
rect 13863 3621 13872 3655
rect 13820 3612 13872 3621
rect 9128 3544 9180 3596
rect 11980 3544 12032 3596
rect 6920 3476 6972 3528
rect 7196 3519 7248 3528
rect 7196 3485 7205 3519
rect 7205 3485 7239 3519
rect 7239 3485 7248 3519
rect 7196 3476 7248 3485
rect 8760 3519 8812 3528
rect 6000 3408 6052 3460
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 9312 3476 9364 3528
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 13912 3476 13964 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 16672 3680 16724 3732
rect 17132 3680 17184 3732
rect 18512 3723 18564 3732
rect 15936 3612 15988 3664
rect 16396 3612 16448 3664
rect 16580 3655 16632 3664
rect 16580 3621 16589 3655
rect 16589 3621 16623 3655
rect 16623 3621 16632 3655
rect 16580 3612 16632 3621
rect 18512 3689 18521 3723
rect 18521 3689 18555 3723
rect 18555 3689 18564 3723
rect 18512 3680 18564 3689
rect 23664 3723 23716 3732
rect 23664 3689 23673 3723
rect 23673 3689 23707 3723
rect 23707 3689 23716 3723
rect 23664 3680 23716 3689
rect 17684 3612 17736 3664
rect 18328 3544 18380 3596
rect 19340 3587 19392 3596
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 19340 3544 19392 3553
rect 21732 3544 21784 3596
rect 22284 3544 22336 3596
rect 23020 3544 23072 3596
rect 24676 3680 24728 3732
rect 24216 3612 24268 3664
rect 24124 3587 24176 3596
rect 24124 3553 24133 3587
rect 24133 3553 24167 3587
rect 24167 3553 24176 3587
rect 24124 3544 24176 3553
rect 14096 3476 14148 3485
rect 5448 3340 5500 3392
rect 6092 3340 6144 3392
rect 6184 3340 6236 3392
rect 12532 3408 12584 3460
rect 13452 3451 13504 3460
rect 13452 3417 13461 3451
rect 13461 3417 13495 3451
rect 13495 3417 13504 3451
rect 13452 3408 13504 3417
rect 20168 3476 20220 3528
rect 23112 3476 23164 3528
rect 16488 3408 16540 3460
rect 17316 3408 17368 3460
rect 22560 3451 22612 3460
rect 22560 3417 22569 3451
rect 22569 3417 22603 3451
rect 22603 3417 22612 3451
rect 22560 3408 22612 3417
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 10692 3340 10744 3392
rect 12624 3340 12676 3392
rect 14556 3340 14608 3392
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 20260 3340 20312 3392
rect 21364 3383 21416 3392
rect 21364 3349 21373 3383
rect 21373 3349 21407 3383
rect 21407 3349 21416 3383
rect 21364 3340 21416 3349
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3240 3136 3292 3188
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6460 3179 6512 3188
rect 6460 3145 6469 3179
rect 6469 3145 6503 3179
rect 6503 3145 6512 3179
rect 6460 3136 6512 3145
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 8668 3179 8720 3188
rect 8668 3145 8677 3179
rect 8677 3145 8711 3179
rect 8711 3145 8720 3179
rect 10048 3179 10100 3188
rect 8668 3136 8720 3145
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 11704 3136 11756 3188
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 15568 3136 15620 3145
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 17684 3179 17736 3188
rect 17684 3145 17693 3179
rect 17693 3145 17727 3179
rect 17727 3145 17736 3179
rect 17684 3136 17736 3145
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 20168 3179 20220 3188
rect 20168 3145 20177 3179
rect 20177 3145 20211 3179
rect 20211 3145 20220 3179
rect 20168 3136 20220 3145
rect 21732 3179 21784 3188
rect 21732 3145 21741 3179
rect 21741 3145 21775 3179
rect 21775 3145 21784 3179
rect 21732 3136 21784 3145
rect 23020 3136 23072 3188
rect 24124 3136 24176 3188
rect 2872 3000 2924 3052
rect 4896 3000 4948 3052
rect 5356 3000 5408 3052
rect 6276 3000 6328 3052
rect 7196 3000 7248 3052
rect 9404 3000 9456 3052
rect 2412 2975 2464 2984
rect 2412 2941 2456 2975
rect 2456 2941 2464 2975
rect 2412 2932 2464 2941
rect 5264 2932 5316 2984
rect 6092 2932 6144 2984
rect 6368 2932 6420 2984
rect 7288 2932 7340 2984
rect 7840 2975 7892 2984
rect 5080 2864 5132 2916
rect 7380 2864 7432 2916
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 8668 2864 8720 2916
rect 3700 2796 3752 2848
rect 3976 2796 4028 2848
rect 4160 2839 4212 2848
rect 4160 2805 4169 2839
rect 4169 2805 4203 2839
rect 4203 2805 4212 2839
rect 4160 2796 4212 2805
rect 4988 2796 5040 2848
rect 6644 2796 6696 2848
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 18604 3068 18656 3120
rect 22376 3111 22428 3120
rect 22376 3077 22385 3111
rect 22385 3077 22419 3111
rect 22419 3077 22428 3111
rect 22376 3068 22428 3077
rect 23848 3068 23900 3120
rect 10876 3000 10928 3052
rect 11520 3000 11572 3052
rect 16580 3043 16632 3052
rect 16580 3009 16589 3043
rect 16589 3009 16623 3043
rect 16623 3009 16632 3043
rect 16580 3000 16632 3009
rect 18880 3000 18932 3052
rect 21824 3000 21876 3052
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 22560 3000 22612 3052
rect 23388 3000 23440 3052
rect 24216 3000 24268 3052
rect 16948 2932 17000 2984
rect 20168 2932 20220 2984
rect 22192 2975 22244 2984
rect 10692 2864 10744 2916
rect 9680 2796 9732 2848
rect 9956 2796 10008 2848
rect 11888 2864 11940 2916
rect 12624 2907 12676 2916
rect 12624 2873 12633 2907
rect 12633 2873 12667 2907
rect 12667 2873 12676 2907
rect 14556 2907 14608 2916
rect 12624 2864 12676 2873
rect 14556 2873 14565 2907
rect 14565 2873 14599 2907
rect 14599 2873 14608 2907
rect 14556 2864 14608 2873
rect 13544 2796 13596 2848
rect 15752 2864 15804 2916
rect 16120 2907 16172 2916
rect 16120 2873 16129 2907
rect 16129 2873 16163 2907
rect 16163 2873 16172 2907
rect 16120 2864 16172 2873
rect 15568 2796 15620 2848
rect 18512 2864 18564 2916
rect 21180 2864 21232 2916
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 22284 2864 22336 2916
rect 24676 2864 24728 2916
rect 23020 2839 23072 2848
rect 23020 2805 23029 2839
rect 23029 2805 23063 2839
rect 23063 2805 23072 2839
rect 23020 2796 23072 2805
rect 25228 2839 25280 2848
rect 25228 2805 25237 2839
rect 25237 2805 25271 2839
rect 25271 2805 25280 2839
rect 25228 2796 25280 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3700 2592 3752 2644
rect 6644 2635 6696 2644
rect 3240 2567 3292 2576
rect 3240 2533 3249 2567
rect 3249 2533 3283 2567
rect 3283 2533 3292 2567
rect 3240 2524 3292 2533
rect 5080 2567 5132 2576
rect 5080 2533 5089 2567
rect 5089 2533 5123 2567
rect 5123 2533 5132 2567
rect 5080 2524 5132 2533
rect 6000 2524 6052 2576
rect 2044 2456 2096 2508
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 664 2388 716 2440
rect 2964 2320 3016 2372
rect 2044 2295 2096 2304
rect 2044 2261 2053 2295
rect 2053 2261 2087 2295
rect 2087 2261 2096 2295
rect 2044 2252 2096 2261
rect 6920 2456 6972 2508
rect 7840 2592 7892 2644
rect 9220 2524 9272 2576
rect 9680 2592 9732 2644
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 9956 2567 10008 2576
rect 9956 2533 9965 2567
rect 9965 2533 9999 2567
rect 9999 2533 10008 2567
rect 9956 2524 10008 2533
rect 10048 2524 10100 2576
rect 13544 2524 13596 2576
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 7104 2388 7156 2440
rect 8760 2363 8812 2372
rect 8760 2329 8769 2363
rect 8769 2329 8803 2363
rect 8803 2329 8812 2363
rect 16396 2592 16448 2644
rect 19524 2592 19576 2644
rect 20996 2592 21048 2644
rect 15936 2524 15988 2576
rect 18512 2567 18564 2576
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 18788 2524 18840 2576
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 22192 2524 22244 2576
rect 24676 2524 24728 2576
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 21364 2456 21416 2508
rect 22744 2499 22796 2508
rect 22744 2465 22753 2499
rect 22753 2465 22787 2499
rect 22787 2465 22796 2499
rect 22744 2456 22796 2465
rect 8760 2320 8812 2329
rect 13912 2388 13964 2440
rect 15752 2388 15804 2440
rect 14004 2320 14056 2372
rect 16212 2320 16264 2372
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 21272 2431 21324 2440
rect 21272 2397 21281 2431
rect 21281 2397 21315 2431
rect 21315 2397 21324 2431
rect 21272 2388 21324 2397
rect 22100 2388 22152 2440
rect 19248 2320 19300 2372
rect 21640 2320 21692 2372
rect 26148 2456 26200 2508
rect 5540 2252 5592 2304
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 14464 2252 14516 2304
rect 16488 2295 16540 2304
rect 16488 2261 16497 2295
rect 16497 2261 16531 2295
rect 16531 2261 16540 2295
rect 16488 2252 16540 2261
rect 17132 2252 17184 2304
rect 22928 2295 22980 2304
rect 22928 2261 22937 2295
rect 22937 2261 22971 2295
rect 22971 2261 22980 2295
rect 22928 2252 22980 2261
rect 26148 2295 26200 2304
rect 26148 2261 26157 2295
rect 26157 2261 26191 2295
rect 26191 2261 26200 2295
rect 26148 2252 26200 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 4252 2048 4304 2100
rect 12532 2048 12584 2100
rect 7196 76 7248 128
rect 13544 76 13596 128
rect 9680 8 9732 60
rect 10784 8 10836 60
<< metal2 >>
rect 478 27520 534 28000
rect 1490 27520 1546 28000
rect 2594 27554 2650 28000
rect 3698 27554 3754 28000
rect 2594 27526 2912 27554
rect 2594 27520 2650 27526
rect 492 23662 520 27520
rect 1504 23798 1532 27520
rect 2884 23866 2912 27526
rect 3698 27526 3924 27554
rect 3698 27520 3754 27526
rect 3896 23866 3924 27526
rect 4710 27520 4766 28000
rect 5814 27554 5870 28000
rect 5814 27526 6224 27554
rect 5814 27520 5870 27526
rect 4724 24274 4752 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 1492 23792 1544 23798
rect 1492 23734 1544 23740
rect 2884 23662 2912 23802
rect 3896 23662 3924 23802
rect 6196 23798 6224 27526
rect 6918 27520 6974 28000
rect 7930 27520 7986 28000
rect 8300 27532 8352 27538
rect 6932 24818 6960 27520
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6184 23792 6236 23798
rect 6184 23734 6236 23740
rect 7944 23662 7972 27520
rect 9034 27532 9090 28000
rect 9034 27520 9036 27532
rect 8300 27474 8352 27480
rect 9088 27520 9090 27532
rect 9692 27526 10088 27554
rect 9036 27474 9088 27480
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 8024 24064 8076 24070
rect 8024 24006 8076 24012
rect 480 23656 532 23662
rect 480 23598 532 23604
rect 2872 23656 2924 23662
rect 2872 23598 2924 23604
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 2412 23520 2464 23526
rect 2412 23462 2464 23468
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2424 19961 2452 23462
rect 2410 19952 2466 19961
rect 2410 19887 2466 19896
rect 2700 17241 2728 23462
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 2686 17232 2742 17241
rect 2686 17167 2742 17176
rect 6748 16522 6776 23530
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6840 16726 6868 23462
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 7484 14890 7512 16118
rect 7852 15706 7880 23530
rect 8036 16114 8064 24006
rect 8128 23866 8156 24210
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8312 17746 8340 27474
rect 9048 27443 9076 27474
rect 8850 20496 8906 20505
rect 8850 20431 8906 20440
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8128 16250 8156 16662
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8220 16182 8248 16662
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8772 15978 8800 16526
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7392 14414 7420 14826
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 3974 13424 4030 13433
rect 3974 13359 4030 13368
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5030 1440 5714
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 664 2440 716 2446
rect 664 2382 716 2388
rect 386 82 442 480
rect 676 82 704 2382
rect 386 54 704 82
rect 1122 82 1178 480
rect 1412 82 1440 4966
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3620 4282 3648 4626
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3712 4154 3740 4966
rect 3988 4282 4016 13359
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5354 11112 5410 11121
rect 5354 11047 5410 11056
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5184 6798 5212 9318
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 4710 6488 4766 6497
rect 4710 6423 4766 6432
rect 4724 6390 4752 6423
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 5184 6322 5212 6734
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5276 5302 5304 5782
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5078 5128 5134 5137
rect 5078 5063 5134 5072
rect 5092 5030 5120 5063
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 5368 4214 5396 11047
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6458 10568 6514 10577
rect 6458 10503 6514 10512
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9178 6132 9318
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5460 8362 5488 8978
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 7188 5580 7890
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7449 6040 8366
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 5998 7440 6054 7449
rect 5998 7375 6054 7384
rect 5632 7200 5684 7206
rect 5552 7160 5632 7188
rect 5632 7142 5684 7148
rect 5644 6769 5672 7142
rect 6104 6905 6132 8298
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6380 7585 6408 8230
rect 6366 7576 6422 7585
rect 6472 7546 6500 10503
rect 6564 9042 6592 10610
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9654 6684 10066
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8294 6592 8978
rect 6748 8974 6776 13806
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6932 12442 6960 12650
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7484 11626 7512 14826
rect 8220 14822 8248 15574
rect 8772 15502 8800 15914
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8864 14482 8892 20431
rect 9692 18358 9720 27526
rect 10060 27520 10088 27526
rect 10138 27520 10194 28000
rect 11150 27520 11206 28000
rect 12254 27520 12310 28000
rect 13358 27520 13414 28000
rect 14462 27520 14518 28000
rect 15474 27554 15530 28000
rect 16578 27554 16634 28000
rect 15474 27526 15792 27554
rect 15474 27520 15530 27526
rect 10060 27492 10180 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 11164 21078 11192 27520
rect 12072 23588 12124 23594
rect 12072 23530 12124 23536
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10874 18728 10930 18737
rect 10874 18663 10930 18672
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 16017 9168 17682
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8956 14618 8984 14826
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9048 14550 9076 14826
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 13870 7972 14214
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 8864 13734 8892 14418
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7852 12646 7880 12854
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7194 11248 7250 11257
rect 7012 11212 7064 11218
rect 7194 11183 7250 11192
rect 7012 11154 7064 11160
rect 7024 10849 7052 11154
rect 7010 10840 7066 10849
rect 7010 10775 7012 10784
rect 7064 10775 7066 10784
rect 7012 10746 7064 10752
rect 7024 10715 7052 10746
rect 7102 10160 7158 10169
rect 7102 10095 7104 10104
rect 7156 10095 7158 10104
rect 7104 10066 7156 10072
rect 7116 9722 7144 10066
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8430 6776 8910
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6366 7511 6422 7520
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 5630 6760 5686 6769
rect 5630 6695 5686 6704
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5998 6488 6054 6497
rect 5998 6423 6054 6432
rect 6012 6322 6040 6423
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6288 6225 6316 7142
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6274 6216 6330 6225
rect 6274 6151 6330 6160
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 5817 6316 6054
rect 6274 5808 6330 5817
rect 6000 5772 6052 5778
rect 6274 5743 6330 5752
rect 6000 5714 6052 5720
rect 6012 5681 6040 5714
rect 5998 5672 6054 5681
rect 5998 5607 6054 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 3620 4126 3740 4154
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2884 3058 2912 3538
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2056 2310 2084 2450
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1122 54 1440 82
rect 1858 82 1914 480
rect 2056 82 2084 2246
rect 1858 54 2084 82
rect 2424 82 2452 2926
rect 3252 2582 3280 3130
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3054 2408 3110 2417
rect 2964 2372 3016 2378
rect 3016 2352 3054 2360
rect 3016 2343 3110 2352
rect 3016 2332 3096 2343
rect 2964 2314 3016 2320
rect 2686 82 2742 480
rect 2424 54 2742 82
rect 386 0 442 54
rect 1122 0 1178 54
rect 1858 0 1914 54
rect 2686 0 2742 54
rect 3422 82 3478 480
rect 3620 82 3648 4126
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3712 2650 3740 2790
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3988 1873 4016 2790
rect 3974 1864 4030 1873
rect 3974 1799 4030 1808
rect 3422 54 3648 82
rect 4172 82 4200 2790
rect 4264 2106 4292 3878
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4632 3194 4660 3538
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4632 3097 4660 3130
rect 4618 3088 4674 3097
rect 4618 3023 4674 3032
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 4250 82 4306 480
rect 4172 54 4306 82
rect 4908 82 4936 2994
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5000 2689 5028 2790
rect 4986 2680 5042 2689
rect 4986 2615 5042 2624
rect 5092 2582 5120 2858
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5184 785 5212 3878
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5276 3194 5304 3703
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5276 2990 5304 3130
rect 5368 3058 5396 3538
rect 5460 3482 5488 4966
rect 6012 4690 6040 5607
rect 6472 5574 6500 6734
rect 6564 6322 6592 6870
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6276 5568 6328 5574
rect 6460 5568 6512 5574
rect 6328 5545 6408 5556
rect 6328 5536 6422 5545
rect 6328 5528 6366 5536
rect 6276 5510 6328 5516
rect 6460 5510 6512 5516
rect 6366 5471 6422 5480
rect 6366 5400 6422 5409
rect 6472 5370 6500 5510
rect 6366 5335 6422 5344
rect 6460 5364 6512 5370
rect 6380 5302 6408 5335
rect 6460 5306 6512 5312
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5552 4282 5580 4626
rect 5998 4448 6054 4457
rect 5622 4380 5918 4400
rect 5998 4383 6054 4392
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 6012 4214 6040 4383
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5460 3454 5580 3482
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5460 1329 5488 3334
rect 5552 2553 5580 3454
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2582 6040 3402
rect 6196 3398 6224 5102
rect 6472 3602 6500 5170
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6104 2990 6132 3334
rect 6472 3194 6500 3538
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6000 2576 6052 2582
rect 5538 2544 5594 2553
rect 6000 2518 6052 2524
rect 5538 2479 5594 2488
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5446 1320 5502 1329
rect 5446 1255 5502 1264
rect 5170 776 5226 785
rect 5170 711 5226 720
rect 4986 82 5042 480
rect 4908 54 5042 82
rect 5552 82 5580 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6288 1193 6316 2994
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6380 1737 6408 2926
rect 6366 1728 6422 1737
rect 6366 1663 6422 1672
rect 6274 1184 6330 1193
rect 6274 1119 6330 1128
rect 6564 626 6592 5306
rect 6656 5030 6684 5714
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4593 6684 4966
rect 6642 4584 6698 4593
rect 6642 4519 6698 4528
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2650 6684 2790
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6748 2009 6776 5578
rect 6840 4690 6868 8230
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 7024 7886 7052 7919
rect 7012 7880 7064 7886
rect 6918 7848 6974 7857
rect 7012 7822 7064 7828
rect 6918 7783 6974 7792
rect 6932 7750 6960 7783
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7024 7546 7052 7822
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6932 5914 6960 6122
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7116 5166 7144 6394
rect 7208 5370 7236 11183
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7380 9036 7432 9042
rect 7432 8996 7512 9024
rect 7380 8978 7432 8984
rect 7484 8430 7512 8996
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 4690 7144 5102
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6840 4214 6868 4626
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6932 4060 6960 4626
rect 7012 4072 7064 4078
rect 6932 4032 7012 4060
rect 7012 4014 7064 4020
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6734 2000 6790 2009
rect 6734 1935 6790 1944
rect 6840 649 6868 3878
rect 7024 3738 7052 4014
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3369 6960 3470
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 7024 3194 7052 3674
rect 7116 3505 7144 3946
rect 7196 3528 7248 3534
rect 7102 3496 7158 3505
rect 7196 3470 7248 3476
rect 7102 3431 7158 3440
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7208 3058 7236 3470
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7300 2990 7328 8366
rect 7484 8090 7512 8366
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7576 7868 7604 10406
rect 7852 8022 7880 12582
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11558 8064 12242
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10674 7972 11154
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8036 10130 8064 11494
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8036 9382 8064 10066
rect 8128 9722 8156 13466
rect 8496 13394 8524 13670
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 11830 8340 12786
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12442 8432 12718
rect 8496 12714 8524 13330
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8496 12306 8524 12650
rect 8772 12306 8800 13262
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8496 11898 8524 12242
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8496 11218 8524 11834
rect 8588 11762 8616 12174
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8588 11354 8616 11698
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10606 8616 10950
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8588 10130 8616 10542
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8128 9518 8156 9658
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 9042 8064 9318
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8294 8064 8978
rect 8128 8838 8156 9454
rect 8588 9110 8616 9454
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7484 7840 7604 7868
rect 7656 7880 7708 7886
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 5574 7420 6258
rect 7484 5817 7512 7840
rect 7656 7822 7708 7828
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 6798 7604 7686
rect 7668 7546 7696 7822
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7760 7002 7788 7958
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7748 6792 7800 6798
rect 7800 6752 7880 6780
rect 7748 6734 7800 6740
rect 7576 6322 7604 6734
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7470 5808 7526 5817
rect 7470 5743 7526 5752
rect 7576 5642 7604 6258
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7668 5846 7696 6122
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7380 5568 7432 5574
rect 7656 5568 7708 5574
rect 7380 5510 7432 5516
rect 7576 5516 7656 5522
rect 7576 5510 7708 5516
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7392 2922 7420 5510
rect 7576 5494 7696 5510
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7484 5098 7512 5238
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7484 4690 7512 5034
rect 7576 4826 7604 5494
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 4049 7604 4490
rect 7562 4040 7618 4049
rect 7562 3975 7618 3984
rect 7668 3942 7696 5034
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 6920 2508 6972 2514
rect 6972 2468 7052 2496
rect 6920 2450 6972 2456
rect 7024 2428 7052 2468
rect 7104 2440 7156 2446
rect 7024 2400 7104 2428
rect 7104 2382 7156 2388
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 6472 598 6592 626
rect 6826 640 6882 649
rect 5814 82 5870 480
rect 5552 54 5870 82
rect 6472 82 6500 598
rect 6826 575 6882 584
rect 6550 82 6606 480
rect 7208 134 7236 2246
rect 6472 54 6606 82
rect 7196 128 7248 134
rect 7196 70 7248 76
rect 7378 82 7434 480
rect 7760 82 7788 6598
rect 7852 6458 7880 6752
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 4826 7880 5646
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 8036 4672 8064 8230
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 7721 8156 7754
rect 8114 7712 8170 7721
rect 8114 7647 8170 7656
rect 8220 7410 8248 8298
rect 8496 8022 8524 8978
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8498 8616 8910
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8588 8090 8616 8434
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8128 7002 8156 7210
rect 8116 6996 8168 7002
rect 8220 6984 8248 7346
rect 8300 6996 8352 7002
rect 8220 6956 8300 6984
rect 8116 6938 8168 6944
rect 8300 6938 8352 6944
rect 8128 6322 8156 6938
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8404 6322 8432 6870
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8128 5370 8156 6258
rect 8404 5846 8432 6258
rect 8680 6254 8708 9318
rect 8772 8974 8800 9386
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8864 6662 8892 13670
rect 9048 13462 9076 14486
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 9048 12986 9076 13398
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9140 8956 9168 15943
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15162 9628 15506
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13938 9536 14214
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9692 13814 9720 18294
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10782 17232 10838 17241
rect 10782 17167 10838 17176
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16114 9812 16390
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9784 15706 9812 16050
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9692 13786 9812 13814
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9692 12646 9720 13194
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9232 10470 9260 11494
rect 9600 11286 9628 11494
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9324 10266 9352 10950
rect 9416 10810 9444 11154
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 10266 9536 10474
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9232 9518 9260 9658
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9220 9512 9272 9518
rect 9324 9489 9352 9522
rect 9220 9454 9272 9460
rect 9310 9480 9366 9489
rect 9048 8928 9168 8956
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8128 5098 8156 5306
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8312 4690 8340 5102
rect 8496 4826 8524 5102
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8208 4684 8260 4690
rect 8036 4644 8208 4672
rect 8208 4626 8260 4632
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8220 4486 8248 4626
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8404 4078 8432 4558
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7852 2990 7880 3674
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 8390 2952 8446 2961
rect 7852 2650 7880 2926
rect 8390 2887 8446 2896
rect 8404 2854 8432 2887
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 3422 0 3478 54
rect 4250 0 4306 54
rect 4986 0 5042 54
rect 5814 0 5870 54
rect 6550 0 6606 54
rect 7378 54 7788 82
rect 8114 82 8170 480
rect 8588 82 8616 6054
rect 8956 5846 8984 8842
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8680 4214 8708 5034
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8680 3194 8708 3946
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8680 2922 8708 3130
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8772 2378 8800 3470
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 8114 54 8616 82
rect 8850 82 8906 480
rect 8956 82 8984 4218
rect 9048 3210 9076 8928
rect 9232 8362 9260 9454
rect 9310 9415 9366 9424
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 5846 9168 7142
rect 9416 6866 9444 8230
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7206 9536 7890
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9402 6352 9458 6361
rect 9402 6287 9458 6296
rect 9416 6186 9444 6287
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 4622 9168 5510
rect 9508 5234 9536 7142
rect 9600 6254 9628 8502
rect 9692 7750 9720 12582
rect 9784 9217 9812 13786
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9968 12442 9996 13262
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 10060 11830 10088 15914
rect 10152 15706 10180 16118
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10152 15026 10180 15642
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14074 10732 14758
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 12442 10180 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10152 11898 10180 12378
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10060 11286 10088 11766
rect 10152 11626 10180 11834
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11354 10732 12242
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10796 11286 10824 17167
rect 10888 15162 10916 18663
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 13814 10916 15098
rect 10980 14618 11008 15438
rect 11072 15162 11100 15574
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11164 14482 11192 16730
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11348 16114 11376 16594
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11256 15502 11284 15914
rect 11808 15910 11836 16594
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 14890 11284 15438
rect 11348 14958 11376 15846
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11164 14074 11192 14418
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10888 13786 11008 13814
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12714 10916 13126
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10060 10810 10088 11222
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10244 10742 10272 11086
rect 10796 10810 10824 11222
rect 10888 11150 10916 12650
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10198 9996 10678
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 10033 9904 10066
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 9876 9722 9904 9959
rect 9968 9722 9996 10134
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10152 9926 10180 10066
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9770 9208 9826 9217
rect 10152 9178 10180 9862
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10244 9518 10272 9658
rect 10428 9586 10456 9930
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9770 9143 9826 9152
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9784 8634 9812 9046
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9876 8294 9904 9046
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8498 10364 8842
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9784 6458 9812 8026
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9876 6390 9904 6598
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5370 9720 6122
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9968 5302 9996 7686
rect 10152 7546 10180 7890
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10704 7290 10732 10678
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10796 8906 10824 9386
rect 10980 9024 11008 13786
rect 11256 12850 11284 14826
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11440 13802 11468 14554
rect 11808 14006 11836 15846
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11992 14618 12020 15098
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12442 11468 12582
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9178 11100 9522
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10888 8996 11008 9024
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10796 7410 10824 8026
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10704 7262 10824 7290
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10152 5914 10180 6666
rect 10520 6390 10548 6734
rect 10704 6458 10732 6870
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10060 5370 10088 5782
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10140 5704 10192 5710
rect 10428 5681 10456 5714
rect 10140 5646 10192 5652
rect 10414 5672 10470 5681
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4282 9168 4422
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 3602 9168 4082
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9126 3224 9182 3233
rect 9048 3182 9126 3210
rect 9126 3159 9182 3168
rect 9232 2582 9260 4966
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9324 3534 9352 4558
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3670 9444 3878
rect 9784 3738 9812 4762
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 10060 3670 10088 4150
rect 9404 3664 9456 3670
rect 9402 3632 9404 3641
rect 10048 3664 10100 3670
rect 9456 3632 9458 3641
rect 10048 3606 10100 3612
rect 9402 3567 9458 3576
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3058 9444 3334
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9692 2854 9720 3470
rect 10060 3194 10088 3606
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9692 2650 9720 2790
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9968 2582 9996 2790
rect 10046 2680 10102 2689
rect 10046 2615 10102 2624
rect 10060 2582 10088 2615
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 8850 54 8984 82
rect 9678 60 9734 480
rect 7378 0 7434 54
rect 8114 0 8170 54
rect 8850 0 8906 54
rect 9678 8 9680 60
rect 9732 8 9734 60
rect 10152 82 10180 5646
rect 10414 5607 10470 5616
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 2922 10732 3334
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10414 82 10470 480
rect 10152 54 10470 82
rect 10796 66 10824 7262
rect 10888 5710 10916 8996
rect 11164 8906 11192 10066
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 7546 11008 8298
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10980 5001 11008 5102
rect 10966 4992 11022 5001
rect 10966 4927 11022 4936
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10888 4010 10916 4490
rect 10980 4282 11008 4927
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10888 3058 10916 3946
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11072 82 11100 8774
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7478 11192 8298
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11164 5778 11192 7414
rect 11256 6118 11284 10542
rect 11440 10198 11468 11018
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10266 11560 10610
rect 11808 10606 11836 13194
rect 11900 12306 11928 13738
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12753 12020 13330
rect 11978 12744 12034 12753
rect 11978 12679 12034 12688
rect 11992 12646 12020 12679
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11992 9654 12020 12582
rect 12084 10674 12112 23530
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12176 17202 12204 23462
rect 12268 18222 12296 27520
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12360 23662 12388 24754
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 13372 20058 13400 27520
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12268 13802 12296 16050
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12268 10810 12296 11222
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12072 10668 12124 10674
rect 12360 10656 12388 11290
rect 12452 10742 12480 15098
rect 12544 11121 12572 19994
rect 13082 19952 13138 19961
rect 13082 19887 13138 19896
rect 13358 19952 13414 19961
rect 13358 19887 13414 19896
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 15473 12756 15506
rect 12714 15464 12770 15473
rect 12714 15399 12770 15408
rect 12728 15162 12756 15399
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 14618 12756 14758
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12728 13870 12756 14554
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13376 12756 13806
rect 12820 13530 12848 18226
rect 13096 17814 13124 19887
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13096 17338 13124 17750
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13188 17270 13216 17750
rect 13176 17264 13228 17270
rect 13228 17224 13308 17252
rect 13176 17206 13228 17212
rect 13176 16720 13228 16726
rect 13176 16662 13228 16668
rect 13188 15978 13216 16662
rect 13280 16250 13308 17224
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13372 16182 13400 19887
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13556 18154 13584 18294
rect 14476 18222 14504 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 14844 20913 14872 21014
rect 14830 20904 14886 20913
rect 14830 20839 14886 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14384 17610 14412 18022
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 13648 17270 13676 17546
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13648 16522 13676 17206
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13464 16182 13492 16458
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 14016 16114 14044 16390
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 14108 15978 14136 16186
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13096 15026 13124 15302
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13096 14006 13124 14962
rect 13372 14482 13400 15642
rect 13832 15638 13860 15914
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14550 13676 14826
rect 13924 14822 13952 15098
rect 14016 14958 14044 15574
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12808 13388 12860 13394
rect 12728 13348 12808 13376
rect 12992 13388 13044 13394
rect 12860 13348 12940 13376
rect 12808 13330 12860 13336
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12820 11898 12848 12650
rect 12912 12646 12940 13348
rect 12992 13330 13044 13336
rect 13004 12918 13032 13330
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 12102 12940 12582
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11626 12848 11834
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12820 11354 12848 11562
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12808 11144 12860 11150
rect 12530 11112 12586 11121
rect 12808 11086 12860 11092
rect 12530 11047 12586 11056
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12820 10674 12848 11086
rect 12072 10610 12124 10616
rect 12268 10628 12388 10656
rect 12532 10668 12584 10674
rect 12268 10198 12296 10628
rect 12532 10610 12584 10616
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 10198 12388 10474
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12268 9722 12296 10134
rect 12544 10130 12572 10610
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12268 9450 12296 9658
rect 12452 9586 12480 9998
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11348 8090 11376 9114
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8090 11468 8978
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11440 7750 11468 8026
rect 11624 8022 11652 9318
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11900 8294 11928 8978
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11532 6662 11560 7822
rect 11624 7546 11652 7958
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11808 7410 11836 7822
rect 11900 7818 11928 8230
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 6798 11836 7346
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 6497 11652 6598
rect 11610 6488 11666 6497
rect 11610 6423 11666 6432
rect 11900 6322 11928 7754
rect 12164 7268 12216 7274
rect 12268 7256 12296 9386
rect 12452 9178 12480 9522
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12636 9110 12664 10202
rect 12820 10062 12848 10610
rect 12912 10538 12940 12038
rect 13004 11082 13032 12174
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12912 9926 12940 10474
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 13096 9217 13124 13806
rect 13372 13530 13400 14418
rect 13648 13802 13676 14486
rect 14016 13814 14044 14894
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13924 13786 14044 13814
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13188 12850 13216 13262
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13280 10742 13308 12854
rect 13648 12714 13676 13738
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12986 13860 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13648 12374 13676 12650
rect 13924 12442 13952 13786
rect 14108 12986 14136 15914
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 14074 14320 14214
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14292 13802 14320 14010
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14384 13530 14412 13942
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11354 13768 11630
rect 13924 11354 13952 12378
rect 14108 11898 14136 12922
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13372 10470 13400 10610
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13082 9208 13138 9217
rect 13082 9143 13138 9152
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12636 8634 12664 9046
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12216 7228 12296 7256
rect 12164 7210 12216 7216
rect 12268 7002 12296 7228
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 7002 12940 7142
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12268 6458 12296 6938
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4826 11284 5102
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11256 4146 11284 4558
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11256 3738 11284 4082
rect 11348 4010 11376 4422
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11440 2514 11468 5510
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4010 11560 4626
rect 11808 4457 11836 5646
rect 11900 5030 11928 5782
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11794 4448 11850 4457
rect 11794 4383 11850 4392
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11532 3058 11560 3946
rect 11716 3670 11744 4218
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11716 3194 11744 3606
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11900 2922 11928 4966
rect 12268 4758 12296 6394
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5914 12480 6190
rect 12544 6118 12572 6734
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 13096 5914 13124 9143
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8090 13216 8910
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12438 5536 12494 5545
rect 12438 5471 12494 5480
rect 12348 5092 12400 5098
rect 12452 5080 12480 5471
rect 12544 5234 12572 5578
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12532 5092 12584 5098
rect 12452 5052 12532 5080
rect 12348 5034 12400 5040
rect 12532 5034 12584 5040
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12268 4282 12296 4694
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12176 3641 12204 3878
rect 12162 3632 12218 3641
rect 11980 3596 12032 3602
rect 12162 3567 12218 3576
rect 11980 3538 12032 3544
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11992 2650 12020 3538
rect 12360 2650 12388 5034
rect 12544 4826 12572 5034
rect 13096 5030 13124 5850
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 4457 12572 4558
rect 12530 4448 12586 4457
rect 12530 4383 12586 4392
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 3466 12572 3946
rect 12728 3641 12756 4966
rect 13084 4548 13136 4554
rect 13188 4536 13216 5034
rect 13372 5001 13400 10406
rect 13648 10198 13676 10746
rect 13740 10538 13768 11154
rect 13924 10674 13952 11154
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13556 9654 13584 10134
rect 13648 9722 13676 10134
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13464 8294 13492 8434
rect 13556 8362 13584 8570
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13648 8022 13676 9658
rect 14108 9586 14136 9930
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14108 9110 14136 9522
rect 14200 9450 14228 13262
rect 14476 12345 14504 18158
rect 15384 18080 15436 18086
rect 15436 18040 15516 18068
rect 15384 18022 15436 18028
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14660 15638 14688 15914
rect 14752 15638 14780 16934
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14660 15026 14688 15574
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14660 13938 14688 14962
rect 14752 14822 14780 15574
rect 14844 15094 14872 15846
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14752 13814 14780 14758
rect 14936 14618 14964 14826
rect 15304 14618 15332 16050
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15396 15162 15424 15506
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14568 13786 14780 13814
rect 14568 13190 14596 13786
rect 15396 13734 15424 14418
rect 15488 14414 15516 18040
rect 15580 17338 15608 23598
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15580 16114 15608 16458
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 15094 15700 15438
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 14074 15516 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15764 13814 15792 27526
rect 16578 27526 16988 27554
rect 16578 27520 16634 27526
rect 15936 19916 15988 19922
rect 15988 19876 16068 19904
rect 15936 19858 15988 19864
rect 16040 19446 16068 19876
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 17338 15884 18022
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15948 15978 15976 17070
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15672 13786 15792 13814
rect 15948 13802 15976 15914
rect 16040 13814 16068 19382
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16132 18290 16160 18770
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16132 18193 16160 18226
rect 16118 18184 16174 18193
rect 16118 18119 16174 18128
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16132 15910 16160 16594
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16224 14074 16252 16526
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16316 13938 16344 19654
rect 16960 19514 16988 27526
rect 17682 27520 17738 28000
rect 18694 27554 18750 28000
rect 19798 27554 19854 28000
rect 18524 27526 18750 27554
rect 17696 24274 17724 27520
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 18524 23798 18552 27526
rect 18694 27520 18750 27526
rect 19536 27526 19854 27554
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16960 19310 16988 19450
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16500 18902 16528 19110
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17144 17882 17172 18838
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 17066 16528 17478
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16960 16794 16988 17614
rect 17236 17202 17264 18702
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 14890 16528 15302
rect 16684 14890 16712 15846
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17144 15026 17172 15438
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16304 13932 16356 13938
rect 16224 13892 16304 13920
rect 15936 13796 15988 13802
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14462 12336 14518 12345
rect 14462 12271 14518 12280
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14476 11558 14504 12174
rect 14568 11898 14596 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12442 15240 12786
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15212 12170 15240 12378
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 10470 14504 11494
rect 15396 11257 15424 13670
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12850 15516 13262
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15488 11830 15516 12786
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15382 11248 15438 11257
rect 15382 11183 15438 11192
rect 15488 11150 15516 11766
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14554 10840 14610 10849
rect 14554 10775 14610 10784
rect 14568 10674 14596 10775
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13648 7546 13676 7958
rect 13740 7886 13768 8502
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 8022 14136 8298
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7546 13768 7822
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 14200 7274 14228 8842
rect 14292 8090 14320 9862
rect 14660 9722 14688 10950
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 9926 14872 10542
rect 15580 10130 15608 11018
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 15476 9172 15528 9178
rect 15580 9160 15608 10066
rect 15672 9722 15700 13786
rect 16040 13786 16160 13814
rect 15936 13738 15988 13744
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15764 12986 15792 13398
rect 15948 13326 15976 13738
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15764 12442 15792 12922
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15764 10810 15792 11222
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 9178 15700 9318
rect 15528 9132 15608 9160
rect 15660 9172 15712 9178
rect 15476 9114 15528 9120
rect 15660 9114 15712 9120
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8634 15332 8978
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15672 8430 15700 9114
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15028 8294 15056 8366
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 8129 15056 8230
rect 15014 8120 15070 8129
rect 14280 8084 14332 8090
rect 15014 8055 15070 8064
rect 14280 8026 14332 8032
rect 14646 7848 14702 7857
rect 14702 7818 14872 7834
rect 14702 7812 14884 7818
rect 14702 7806 14832 7812
rect 14646 7783 14702 7792
rect 14832 7754 14884 7760
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14646 7576 14702 7585
rect 14646 7511 14702 7520
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14016 6633 14044 6802
rect 14002 6624 14058 6633
rect 14002 6559 14058 6568
rect 14016 6458 14044 6559
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14004 5772 14056 5778
rect 14108 5760 14136 6394
rect 14476 6322 14504 7142
rect 14660 6916 14688 7511
rect 14752 7342 14780 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 15672 7002 15700 8366
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7478 15792 7890
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 14740 6928 14792 6934
rect 14660 6888 14740 6916
rect 14740 6870 14792 6876
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14056 5732 14136 5760
rect 14004 5714 14056 5720
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13358 4992 13414 5001
rect 13358 4927 13414 4936
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13136 4508 13216 4536
rect 13084 4490 13136 4496
rect 13188 4146 13216 4508
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13280 4010 13308 4694
rect 13556 4622 13584 5646
rect 14016 5030 14044 5714
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 12714 3632 12770 3641
rect 12714 3567 12770 3576
rect 13464 3466 13492 4490
rect 13556 3738 13584 4558
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 12624 3392 12676 3398
rect 13464 3369 13492 3402
rect 12624 3334 12676 3340
rect 13450 3360 13506 3369
rect 12636 2922 12664 3334
rect 13450 3295 13506 3304
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 13556 2854 13584 3674
rect 13832 3670 13860 3878
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13740 3194 13768 3606
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13544 2848 13596 2854
rect 13924 2836 13952 3470
rect 14016 2961 14044 4966
rect 14200 4214 14228 5646
rect 14752 5302 14780 5782
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 14752 5166 14780 5238
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14752 4826 14780 5102
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14188 4208 14240 4214
rect 14464 4208 14516 4214
rect 14240 4168 14464 4196
rect 14188 4150 14240 4156
rect 14464 4150 14516 4156
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14002 2952 14058 2961
rect 14002 2887 14058 2896
rect 13924 2808 14044 2836
rect 13544 2790 13596 2796
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 13556 2582 13584 2790
rect 13544 2576 13596 2582
rect 12070 2544 12126 2553
rect 11428 2508 11480 2514
rect 13544 2518 13596 2524
rect 12070 2479 12126 2488
rect 11428 2450 11480 2456
rect 11242 82 11298 480
rect 9678 0 9734 8
rect 10414 0 10470 54
rect 10784 60 10836 66
rect 11072 54 11298 82
rect 10784 2 10836 8
rect 11242 0 11298 54
rect 11978 82 12034 480
rect 12084 82 12112 2479
rect 13912 2440 13964 2446
rect 13832 2417 13912 2428
rect 13818 2408 13912 2417
rect 13874 2400 13912 2408
rect 13912 2382 13964 2388
rect 14016 2378 14044 2808
rect 13818 2343 13874 2352
rect 14004 2372 14056 2378
rect 14004 2314 14056 2320
rect 12532 2100 12584 2106
rect 12532 2042 12584 2048
rect 11978 54 12112 82
rect 12544 82 12572 2042
rect 14108 1737 14136 3470
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 2922 14596 3334
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14200 2417 14228 2450
rect 14186 2408 14242 2417
rect 14186 2343 14242 2352
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14094 1728 14150 1737
rect 14094 1663 14150 1672
rect 12806 82 12862 480
rect 12544 54 12862 82
rect 11978 0 12034 54
rect 12806 0 12862 54
rect 13542 128 13598 480
rect 13542 76 13544 128
rect 13596 76 13598 128
rect 13542 0 13598 76
rect 14370 82 14426 480
rect 14476 82 14504 2246
rect 14568 1873 14596 2858
rect 14554 1864 14610 1873
rect 14554 1799 14610 1808
rect 14370 54 14504 82
rect 14844 82 14872 6666
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 5642 15332 6734
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15382 5944 15438 5953
rect 15382 5879 15438 5888
rect 15396 5778 15424 5879
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 5370 15424 5714
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15396 4593 15424 5306
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15488 4622 15516 5034
rect 15476 4616 15528 4622
rect 15382 4584 15438 4593
rect 15476 4558 15528 4564
rect 15382 4519 15438 4528
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15488 3738 15516 4558
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15580 3194 15608 6190
rect 15672 6186 15700 6938
rect 15856 6390 15884 12106
rect 15948 11830 15976 12310
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15948 10198 15976 11766
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15948 6662 15976 9658
rect 16040 7954 16068 13262
rect 16132 13258 16160 13786
rect 16224 13530 16252 13892
rect 16304 13874 16356 13880
rect 16408 13814 16436 14010
rect 16316 13802 16436 13814
rect 16304 13796 16436 13802
rect 16356 13786 16436 13796
rect 16304 13738 16356 13744
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16500 13433 16528 14826
rect 16684 14550 16712 14826
rect 17328 14618 17356 23598
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17512 19446 17540 23530
rect 18892 20058 18920 24006
rect 19168 23798 19196 24210
rect 19536 23866 19564 27526
rect 19798 27520 19854 27526
rect 20902 27520 20958 28000
rect 21914 27520 21970 28000
rect 23018 27554 23074 28000
rect 22756 27526 23074 27554
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20916 24410 20944 27520
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19996 23526 20024 24210
rect 21928 23866 21956 27520
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 22756 23798 22784 27526
rect 23018 27520 23074 27526
rect 24122 27520 24178 28000
rect 25134 27554 25190 28000
rect 24872 27526 25190 27554
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20812 23588 20864 23594
rect 20812 23530 20864 23536
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19996 20505 20024 23462
rect 20732 20992 20760 23462
rect 20824 21146 20852 23530
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20812 21004 20864 21010
rect 20732 20964 20812 20992
rect 20812 20946 20864 20952
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 19514 19104 19790
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 17500 19440 17552 19446
rect 19076 19417 19104 19450
rect 17500 19382 17552 19388
rect 19062 19408 19118 19417
rect 19062 19343 19118 19352
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17420 18086 17448 18838
rect 18432 18630 18460 19246
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18156 18290 18184 18566
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17420 17814 17448 18022
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 17338 17448 17750
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17972 17066 18000 18022
rect 18156 17882 18184 18226
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16794 18000 17002
rect 18432 16998 18460 18566
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18524 17678 18552 18226
rect 18616 17814 18644 19110
rect 19260 18970 19288 19654
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 17202 18552 17478
rect 18616 17338 18644 17750
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19168 17649 19196 17682
rect 19154 17640 19210 17649
rect 19154 17575 19210 17584
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 19168 17202 19196 17575
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18616 16794 18644 17002
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 19156 16720 19208 16726
rect 19260 16708 19288 17138
rect 19208 16680 19288 16708
rect 19156 16662 19208 16668
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 15978 17540 16526
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17788 15910 17816 16662
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17512 14890 17540 15574
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 16486 13424 16542 13433
rect 16486 13359 16542 13368
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16684 13190 16712 14486
rect 17236 13938 17264 14486
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17328 13870 17356 14554
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17420 13734 17448 14350
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16684 12442 16712 13126
rect 17420 12850 17448 13670
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12986 17540 13330
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 17316 12368 17368 12374
rect 16762 12336 16818 12345
rect 17316 12310 17368 12316
rect 16762 12271 16818 12280
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16224 10588 16252 10950
rect 16396 10600 16448 10606
rect 16224 10560 16396 10588
rect 16224 10033 16252 10560
rect 16396 10542 16448 10548
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16210 10024 16266 10033
rect 16210 9959 16266 9968
rect 16118 9752 16174 9761
rect 16118 9687 16174 9696
rect 16132 8294 16160 9687
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16224 9178 16252 9386
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16316 9042 16344 10406
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16408 8362 16436 9114
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16408 8090 16436 8298
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16040 7546 16068 7890
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15580 2854 15608 3130
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15106 82 15162 480
rect 14844 54 15162 82
rect 15672 82 15700 5510
rect 15948 5302 15976 6598
rect 16040 5914 16068 7482
rect 16132 7002 16160 7822
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7274 16436 7686
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16132 6322 16160 6938
rect 16408 6662 16436 7210
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15764 3942 15792 4762
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4282 16252 4422
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16224 4010 16252 4218
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 16408 3670 16436 6598
rect 16500 5166 16528 10474
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 8498 16620 8774
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16592 5166 16620 5850
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 16396 3664 16448 3670
rect 16500 3641 16528 5102
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16592 4214 16620 4422
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16592 3670 16620 4150
rect 16684 4146 16712 5578
rect 16776 4690 16804 12271
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17052 11898 17080 12174
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17328 11830 17356 12310
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 10985 17080 11494
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 11014 17356 11086
rect 17696 11014 17724 15030
rect 18156 14890 18184 16390
rect 18616 16114 18644 16526
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15706 18644 16050
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18708 15638 18736 16390
rect 19168 16182 19196 16662
rect 19156 16176 19208 16182
rect 18878 16144 18934 16153
rect 18788 16108 18840 16114
rect 19156 16118 19208 16124
rect 18878 16079 18934 16088
rect 18788 16050 18840 16056
rect 18800 16017 18828 16050
rect 18786 16008 18842 16017
rect 18786 15943 18842 15952
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18892 15502 18920 16079
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 15026 18920 15438
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 17960 14884 18012 14890
rect 18144 14884 18196 14890
rect 18012 14844 18092 14872
rect 17960 14826 18012 14832
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14618 17908 14758
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17316 11008 17368 11014
rect 17038 10976 17094 10985
rect 17316 10950 17368 10956
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17038 10911 17094 10920
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9586 17080 9862
rect 17236 9722 17264 10202
rect 17328 10198 17356 10950
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8634 17264 9046
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17144 7546 17172 7958
rect 17328 7886 17356 10134
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16960 6662 16988 7346
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 17236 6254 17264 6870
rect 17420 6798 17448 7210
rect 17512 6798 17540 10950
rect 17880 10742 17908 11222
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17788 10470 17816 10542
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 9110 17816 10406
rect 17972 9466 18000 13670
rect 18064 11762 18092 14844
rect 18144 14826 18196 14832
rect 18156 14550 18184 14826
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 13326 18184 14214
rect 18248 14074 18276 14486
rect 18432 14414 18460 14962
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18156 11694 18184 13126
rect 18800 12850 18828 13398
rect 18892 13190 18920 14758
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18984 14006 19012 14282
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18984 13002 19012 13262
rect 18892 12974 19012 13002
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18156 11354 18184 11630
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18616 11121 18644 11630
rect 18418 11112 18474 11121
rect 18328 11076 18380 11082
rect 18418 11047 18474 11056
rect 18602 11112 18658 11121
rect 18602 11047 18658 11056
rect 18328 11018 18380 11024
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18064 10266 18092 10542
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18340 10062 18368 11018
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18432 9602 18460 11047
rect 18708 10577 18736 12038
rect 18800 11626 18828 12786
rect 18892 12646 18920 12974
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18694 10568 18750 10577
rect 18800 10538 18828 11562
rect 18892 10810 18920 12582
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18694 10503 18750 10512
rect 18788 10532 18840 10538
rect 18708 9994 18736 10503
rect 18788 10474 18840 10480
rect 18984 10266 19012 12718
rect 19076 12306 19104 14826
rect 19352 14074 19380 20334
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19444 18154 19472 18838
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19536 16726 19564 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19996 19854 20024 20431
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20088 19378 20116 19994
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20180 18290 20208 20742
rect 20824 20262 20852 20946
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20180 17882 20208 18226
rect 20272 18154 20300 19314
rect 20456 18902 20484 20198
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20732 18766 20760 19178
rect 20720 18760 20772 18766
rect 20824 18737 20852 20198
rect 20916 19961 20944 23598
rect 23124 23526 23152 24210
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 20902 19952 20958 19961
rect 20902 19887 20958 19896
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21008 19378 21036 19858
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21192 19242 21220 19654
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21192 18902 21220 19178
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 20720 18702 20772 18708
rect 20810 18728 20866 18737
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16720 19576 16726
rect 19444 16680 19524 16708
rect 19444 15570 19472 16680
rect 19524 16662 19576 16668
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 19996 16046 20024 16662
rect 20180 16046 20208 16934
rect 20272 16794 20300 18090
rect 20732 17678 20760 18702
rect 20810 18663 20866 18672
rect 21008 17882 21036 18838
rect 21192 18426 21220 18838
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21468 18290 21496 18702
rect 21560 18426 21588 19178
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21560 18086 21588 18362
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 21652 17814 21680 19246
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 21652 17338 21680 17750
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20548 16046 20576 17002
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19536 15706 19564 15914
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 20180 15638 20208 15982
rect 20548 15706 20576 15982
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 20444 15632 20496 15638
rect 20444 15574 20496 15580
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19444 15162 19472 15506
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20180 15162 20208 15370
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20180 14958 20208 15098
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20364 14822 20392 15438
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 12782 19196 13874
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13394 19380 13670
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 12442 19196 12718
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19076 11354 19104 12242
rect 19352 11898 19380 12582
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19064 11348 19116 11354
rect 19116 11308 19196 11336
rect 19064 11290 19116 11296
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18788 10056 18840 10062
rect 18786 10024 18788 10033
rect 18840 10024 18842 10033
rect 18696 9988 18748 9994
rect 18786 9959 18842 9968
rect 18696 9930 18748 9936
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18340 9574 18460 9602
rect 18800 9586 18828 9959
rect 19076 9722 19104 10066
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18788 9580 18840 9586
rect 17880 9438 18000 9466
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17696 8294 17724 8910
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 8090 17724 8230
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17788 6905 17816 8910
rect 17774 6896 17830 6905
rect 17774 6831 17830 6840
rect 17408 6792 17460 6798
rect 17328 6752 17408 6780
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16960 4826 16988 5850
rect 17052 5846 17080 6054
rect 17328 5914 17356 6752
rect 17408 6734 17460 6740
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17774 6760 17830 6769
rect 17512 6458 17540 6734
rect 17774 6695 17776 6704
rect 17828 6695 17830 6704
rect 17776 6666 17828 6672
rect 17788 6458 17816 6666
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17420 5370 17448 5782
rect 17880 5370 17908 9438
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9178 18000 9318
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18248 8838 18276 9522
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8362 18276 8774
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7546 18000 7890
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17972 5273 18000 5510
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16776 4146 16804 4626
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16684 3738 16712 4082
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16580 3664 16632 3670
rect 16396 3606 16448 3612
rect 16486 3632 16542 3641
rect 15948 3194 15976 3606
rect 16580 3606 16632 3612
rect 16486 3567 16542 3576
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15764 2446 15792 2858
rect 15948 2582 15976 3130
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16132 2360 16160 2858
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16212 2372 16264 2378
rect 16132 2332 16212 2360
rect 16132 785 16160 2332
rect 16212 2314 16264 2320
rect 16118 776 16174 785
rect 16118 711 16174 720
rect 15842 82 15898 480
rect 15672 54 15898 82
rect 16408 82 16436 2586
rect 16500 2310 16528 3402
rect 16592 3058 16620 3606
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16500 1329 16528 2246
rect 16486 1320 16542 1329
rect 16486 1255 16542 1264
rect 16776 1193 16804 4082
rect 16960 2990 16988 4762
rect 17144 3738 17172 5034
rect 18064 4729 18092 6598
rect 18050 4720 18106 4729
rect 18050 4655 18106 4664
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17696 3670 17724 3946
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17144 2310 17172 2450
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17144 2009 17172 2246
rect 17130 2000 17186 2009
rect 17130 1935 17186 1944
rect 16762 1184 16818 1193
rect 16762 1119 16818 1128
rect 16670 82 16726 480
rect 16408 54 16726 82
rect 17328 82 17356 3402
rect 17696 3194 17724 3606
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17406 82 17462 480
rect 17328 54 17462 82
rect 17972 82 18000 4422
rect 18156 4146 18184 4490
rect 18248 4486 18276 7142
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18340 3602 18368 9574
rect 18788 9522 18840 9528
rect 19076 9217 19104 9658
rect 19062 9208 19118 9217
rect 19062 9143 19118 9152
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18432 2961 18460 8230
rect 18984 7954 19012 9046
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18984 7546 19012 7890
rect 19062 7848 19118 7857
rect 19062 7783 19118 7792
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 19076 7478 19104 7783
rect 19064 7472 19116 7478
rect 18694 7440 18750 7449
rect 19064 7414 19116 7420
rect 18694 7375 18696 7384
rect 18748 7375 18750 7384
rect 18696 7346 18748 7352
rect 18708 7002 18736 7346
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18984 6458 19012 6870
rect 19076 6633 19104 7142
rect 19062 6624 19118 6633
rect 19062 6559 19118 6568
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18604 5840 18656 5846
rect 18524 5800 18604 5828
rect 18524 5030 18552 5800
rect 18604 5782 18656 5788
rect 18708 5409 18736 6054
rect 18694 5400 18750 5409
rect 19076 5370 19104 6559
rect 19168 6322 19196 11308
rect 19340 11212 19392 11218
rect 19260 11172 19340 11200
rect 19260 10470 19288 11172
rect 19340 11154 19392 11160
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10130 19288 10406
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19444 7410 19472 14418
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19536 13852 19564 14010
rect 20088 13870 20116 14282
rect 20364 13870 20392 14758
rect 20456 14006 20484 15574
rect 20548 14940 20576 15642
rect 20732 15094 20760 16390
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15570 20852 15846
rect 21008 15706 21036 17070
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21284 16726 21312 17002
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 20824 15366 20852 15506
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20824 15026 20852 15302
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20628 14952 20680 14958
rect 20548 14912 20628 14940
rect 20628 14894 20680 14900
rect 20824 14346 20852 14962
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 19616 13864 19668 13870
rect 19536 13824 19616 13852
rect 19536 13530 19564 13824
rect 19616 13806 19668 13812
rect 20076 13864 20128 13870
rect 20352 13864 20404 13870
rect 20076 13806 20128 13812
rect 20272 13812 20352 13814
rect 20272 13806 20404 13812
rect 20272 13786 20392 13806
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19536 12782 19564 13466
rect 20272 13190 20300 13786
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19536 12170 19564 12718
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19536 11762 19564 12106
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19536 10470 19564 10678
rect 20180 10606 20208 12242
rect 20272 12170 20300 13126
rect 20364 12782 20392 13126
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20364 12102 20392 12718
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11286 20392 12038
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19536 9586 19564 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 20088 9926 20116 10406
rect 20180 9926 20208 10542
rect 20456 10130 20484 13942
rect 20824 13938 20852 14282
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19536 8906 19564 9386
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19536 8090 19564 8842
rect 19720 8634 19748 8978
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19890 8528 19946 8537
rect 19890 8463 19946 8472
rect 19904 8430 19932 8463
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19996 8362 20024 9046
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8090 20024 8298
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19536 7993 19564 8026
rect 19522 7984 19578 7993
rect 19522 7919 19578 7928
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19168 5828 19196 6258
rect 19338 6216 19394 6225
rect 19338 6151 19394 6160
rect 19352 6118 19380 6151
rect 19444 6118 19472 6734
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19444 5914 19472 6054
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19248 5840 19300 5846
rect 19168 5800 19248 5828
rect 19248 5782 19300 5788
rect 18694 5335 18750 5344
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18602 4992 18658 5001
rect 18524 4758 18552 4966
rect 18602 4927 18658 4936
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18524 3738 18552 3946
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18418 2952 18474 2961
rect 18524 2922 18552 3674
rect 18616 3126 18644 4927
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18418 2887 18474 2896
rect 18512 2916 18564 2922
rect 18432 2632 18460 2887
rect 18512 2858 18564 2864
rect 18340 2604 18460 2632
rect 18340 649 18368 2604
rect 18524 2582 18552 2858
rect 18800 2582 18828 5238
rect 19340 5092 19392 5098
rect 19536 5080 19564 6598
rect 19812 6254 19840 6802
rect 19996 6254 20024 7414
rect 20088 7274 20116 9862
rect 20456 9178 20484 10066
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20548 7342 20576 12582
rect 20640 12374 20668 12786
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20640 11830 20668 12310
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20916 11694 20944 13942
rect 21008 13190 21036 14894
rect 21100 14618 21128 15370
rect 21744 14890 21772 15506
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21836 14822 21864 15506
rect 21928 15094 21956 16118
rect 22020 15473 22048 21082
rect 22560 19916 22612 19922
rect 22560 19858 22612 19864
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22204 17814 22232 18226
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 17338 22232 17614
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22112 16114 22140 16730
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22204 16250 22232 16526
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22006 15464 22062 15473
rect 22006 15399 22062 15408
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21100 14414 21128 14554
rect 21836 14550 21864 14758
rect 21824 14544 21876 14550
rect 21824 14486 21876 14492
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21100 14074 21128 14350
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 13530 21128 14010
rect 21744 13734 21772 14418
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21560 13326 21588 13670
rect 21744 13394 21772 13670
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21560 12646 21588 13262
rect 21744 13190 21772 13330
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21928 12374 21956 15030
rect 22020 13870 22048 15399
rect 22204 15162 22232 15914
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22204 14482 22232 14758
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 12714 22140 13670
rect 22388 13394 22416 14418
rect 22480 13814 22508 19654
rect 22572 19514 22600 19858
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 18290 23060 18770
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 23492 18193 23520 24686
rect 24136 23866 24164 27520
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 25327
rect 24872 24138 24900 27526
rect 25134 27520 25190 27526
rect 26238 27520 26294 28000
rect 27342 27520 27398 28000
rect 25226 27024 25282 27033
rect 25226 26959 25282 26968
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24858 24032 24914 24041
rect 24858 23967 24914 23976
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24872 23474 24900 23967
rect 25148 23866 25176 24210
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25148 23474 25176 23802
rect 24780 23446 24900 23474
rect 25056 23446 25176 23474
rect 24780 23322 24808 23446
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23860 19174 23888 19858
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23478 18184 23534 18193
rect 23112 18148 23164 18154
rect 23478 18119 23534 18128
rect 23112 18090 23164 18096
rect 23124 17814 23152 18090
rect 23112 17808 23164 17814
rect 23112 17750 23164 17756
rect 23124 17338 23152 17750
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23388 17604 23440 17610
rect 23388 17546 23440 17552
rect 23400 17338 23428 17546
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23020 17060 23072 17066
rect 23020 17002 23072 17008
rect 23032 16726 23060 17002
rect 23584 16726 23612 17614
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23032 16250 23060 16662
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23860 16153 23888 19110
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 17066 24072 18022
rect 24136 17882 24164 22374
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22607
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24766 21312 24822 21321
rect 24766 21247 24822 21256
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24780 20602 24808 21247
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24596 20058 24624 20334
rect 24766 20088 24822 20097
rect 24584 20052 24636 20058
rect 24766 20023 24822 20032
rect 24584 19994 24636 20000
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24780 19514 24808 20023
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24228 18222 24256 18566
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24136 17202 24164 17818
rect 24596 17649 24624 18022
rect 24688 17746 24716 18566
rect 24780 18086 24808 18770
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24582 17640 24638 17649
rect 24582 17575 24638 17584
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17338 24716 17682
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 24044 16794 24072 17002
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23846 16144 23902 16153
rect 23846 16079 23902 16088
rect 24044 15706 24072 16730
rect 24504 16726 24532 16934
rect 24492 16720 24544 16726
rect 24544 16680 24716 16708
rect 24492 16662 24544 16668
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24308 16108 24360 16114
rect 24228 16068 24308 16096
rect 24228 15978 24256 16068
rect 24308 16050 24360 16056
rect 24216 15972 24268 15978
rect 24216 15914 24268 15920
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23388 15632 23440 15638
rect 23388 15574 23440 15580
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22848 14074 22876 14418
rect 22940 14278 22968 15438
rect 23400 15094 23428 15574
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23112 14884 23164 14890
rect 23112 14826 23164 14832
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22480 13786 22600 13814
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22112 12442 22140 12650
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21192 11694 21220 12174
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 20916 11218 20944 11630
rect 21192 11218 21220 11630
rect 21376 11354 21404 12174
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 22020 11694 22048 12106
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21744 11218 21772 11494
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 20916 10742 20944 11154
rect 21192 10810 21220 11154
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20640 9178 20668 9930
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20640 8498 20668 9114
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20824 8430 20852 8978
rect 20916 8634 20944 10678
rect 21744 10470 21772 11154
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 21008 9450 21036 9930
rect 21376 9926 21404 10066
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 21376 9382 21404 9862
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 21284 8430 21312 8978
rect 21376 8566 21404 9318
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 8022 20668 8230
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20640 7478 20668 7958
rect 20824 7936 20852 8366
rect 21284 8022 21312 8366
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 20996 7948 21048 7954
rect 20824 7908 20996 7936
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5914 20024 6190
rect 20088 5914 20116 7210
rect 20548 7002 20576 7278
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20824 6866 20852 7908
rect 20996 7890 21048 7896
rect 20996 7812 21048 7818
rect 21048 7772 21128 7800
rect 20996 7754 21048 7760
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20272 5778 20300 6802
rect 21008 6497 21036 7142
rect 20994 6488 21050 6497
rect 20994 6423 21050 6432
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19628 5273 19656 5646
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19614 5264 19670 5273
rect 19614 5199 19670 5208
rect 19628 5166 19656 5199
rect 19996 5166 20024 5306
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19392 5052 19564 5080
rect 19340 5034 19392 5040
rect 19536 4826 19564 5052
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4826 20024 5102
rect 20456 4826 20484 5238
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19168 4282 19196 4626
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19996 4154 20024 4762
rect 20456 4214 20484 4762
rect 20824 4690 20852 4966
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4282 20852 4626
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20444 4208 20496 4214
rect 19996 4126 20116 4154
rect 20444 4150 20496 4156
rect 20088 4078 20116 4126
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20088 3942 20116 4014
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 18878 3496 18934 3505
rect 18878 3431 18934 3440
rect 18892 3398 18920 3431
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3058 18920 3334
rect 19352 3194 19380 3538
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20180 3194 20208 3470
rect 20272 3398 20300 4014
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 20180 2990 20208 3130
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 18512 2576 18564 2582
rect 18418 2544 18474 2553
rect 18512 2518 18564 2524
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18418 2479 18474 2488
rect 18432 2446 18460 2479
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 18326 640 18382 649
rect 18326 575 18382 584
rect 18234 82 18290 480
rect 17972 54 18290 82
rect 14370 0 14426 54
rect 15106 0 15162 54
rect 15842 0 15898 54
rect 16670 0 16726 54
rect 17406 0 17462 54
rect 18234 0 18290 54
rect 18970 82 19026 480
rect 19260 82 19288 2314
rect 18970 54 19288 82
rect 19536 82 19564 2586
rect 19798 82 19854 480
rect 19536 54 19854 82
rect 18970 0 19026 54
rect 19798 0 19854 54
rect 20534 82 20590 480
rect 20916 82 20944 6326
rect 21100 4154 21128 7772
rect 21284 6866 21312 7958
rect 21376 7410 21404 8502
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21192 4282 21220 6122
rect 21468 5846 21496 9386
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21652 7750 21680 8910
rect 21928 8430 21956 8978
rect 22020 8974 22048 11630
rect 22296 10810 22324 12650
rect 22480 12646 22508 13126
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21744 7954 21772 8230
rect 21928 8090 21956 8366
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 21744 6866 21772 7414
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21836 6866 21864 7210
rect 22204 6866 22232 9590
rect 22296 9586 22324 9862
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22296 8498 22324 9522
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22480 8294 22508 12582
rect 22572 8430 22600 13786
rect 22940 13462 22968 14214
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22664 11354 22692 12242
rect 22756 11762 22784 12650
rect 23020 12368 23072 12374
rect 22940 12328 23020 12356
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22940 11558 22968 12328
rect 23020 12310 23072 12316
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 11626 23060 12174
rect 23020 11620 23072 11626
rect 23020 11562 23072 11568
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22664 10606 22692 11290
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22848 9489 22876 9998
rect 22834 9480 22890 9489
rect 22940 9450 22968 11494
rect 23032 11354 23060 11562
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22834 9415 22890 9424
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22480 7750 22508 7890
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 21744 6322 21772 6802
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 22020 6254 22048 6598
rect 22480 6322 22508 7686
rect 22940 7206 22968 7822
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21376 5370 21404 5714
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21008 4126 21128 4154
rect 21008 2650 21036 4126
rect 21192 2922 21220 4218
rect 21376 4154 21404 5306
rect 21468 4214 21496 5510
rect 22020 5166 22048 6190
rect 22112 5574 22140 6190
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22112 5166 22140 5510
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 21560 4486 21588 5102
rect 22112 4826 22140 5102
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22296 4622 22324 5102
rect 22388 4672 22416 6190
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22480 5370 22508 5714
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22572 5234 22600 7142
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22560 4684 22612 4690
rect 22388 4644 22560 4672
rect 22560 4626 22612 4632
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21284 4126 21404 4154
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21180 2916 21232 2922
rect 21180 2858 21232 2864
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21192 2514 21220 2858
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21284 2446 21312 4126
rect 21560 4060 21588 4422
rect 22572 4214 22600 4626
rect 22756 4554 22784 5510
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 22940 4146 22968 7142
rect 23032 6662 23060 7822
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23032 5137 23060 6598
rect 23018 5128 23074 5137
rect 23018 5063 23074 5072
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 21732 4072 21784 4078
rect 21560 4032 21732 4060
rect 21732 4014 21784 4020
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21744 3602 21772 4014
rect 21836 3942 21864 4014
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21376 2514 21404 3334
rect 21744 3194 21772 3538
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21836 3058 21864 3878
rect 22374 3632 22430 3641
rect 22284 3596 22336 3602
rect 22374 3567 22430 3576
rect 22284 3538 22336 3544
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 21364 2508 21416 2514
rect 21364 2450 21416 2456
rect 22112 2446 22140 2994
rect 22204 2990 22232 3334
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22204 2582 22232 2926
rect 22296 2922 22324 3538
rect 22388 3126 22416 3567
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22572 3058 22600 3402
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 21640 2372 21692 2378
rect 21640 2314 21692 2320
rect 20534 54 20944 82
rect 21362 82 21418 480
rect 21652 82 21680 2314
rect 21362 54 21680 82
rect 22098 82 22154 480
rect 22296 82 22324 2858
rect 22756 2514 22784 3946
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23032 3602 23060 3878
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 22926 3360 22982 3369
rect 22926 3295 22982 3304
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22940 2310 22968 3295
rect 23032 3194 23060 3538
rect 23124 3534 23152 14826
rect 23676 14618 23704 14894
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23952 14482 23980 15098
rect 24030 14648 24086 14657
rect 24136 14618 24164 15846
rect 24228 14958 24256 15914
rect 24688 15638 24716 16680
rect 24780 16590 24808 17002
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24780 16182 24808 16526
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24780 15706 24808 16118
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24030 14583 24086 14592
rect 24124 14612 24176 14618
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23952 14074 23980 14418
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 24044 13814 24072 14583
rect 24124 14554 24176 14560
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24872 14074 24900 19246
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24964 15162 24992 15506
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 23952 13786 24072 13814
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23768 11762 23796 12106
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23216 10470 23244 11154
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23216 10198 23244 10406
rect 23492 10198 23520 10610
rect 23204 10192 23256 10198
rect 23480 10192 23532 10198
rect 23204 10134 23256 10140
rect 23400 10140 23480 10146
rect 23400 10134 23532 10140
rect 23216 9382 23244 10134
rect 23400 10118 23520 10134
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23216 8004 23244 9318
rect 23308 8634 23336 9862
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23400 8498 23428 10118
rect 23572 9988 23624 9994
rect 23572 9930 23624 9936
rect 23584 9722 23612 9930
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23584 9110 23612 9386
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23584 8294 23612 9046
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23860 8362 23888 8570
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23296 8016 23348 8022
rect 23216 7976 23296 8004
rect 23296 7958 23348 7964
rect 23308 7546 23336 7958
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23584 7002 23612 8230
rect 23768 8090 23796 8298
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23308 5914 23336 6734
rect 23584 6118 23612 6938
rect 23756 6180 23808 6186
rect 23756 6122 23808 6128
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23768 5710 23796 6122
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23676 5166 23704 5646
rect 23768 5273 23796 5646
rect 23860 5302 23888 5782
rect 23848 5296 23900 5302
rect 23754 5264 23810 5273
rect 23848 5238 23900 5244
rect 23754 5199 23810 5208
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 23492 4690 23520 5034
rect 23676 5030 23704 5102
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23768 4690 23796 5102
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23664 4208 23716 4214
rect 23664 4150 23716 4156
rect 23952 4154 23980 13786
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12714 24072 13126
rect 24032 12708 24084 12714
rect 24032 12650 24084 12656
rect 24136 12442 24164 13330
rect 24228 12850 24256 13670
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24030 12200 24086 12209
rect 24030 12135 24086 12144
rect 24044 10985 24072 12135
rect 24136 11626 24164 12378
rect 24228 11762 24256 12786
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11830 24716 12174
rect 24780 11898 24808 12310
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24124 11620 24176 11626
rect 24124 11562 24176 11568
rect 24136 11354 24164 11562
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24030 10976 24086 10985
rect 24030 10911 24086 10920
rect 24030 10704 24086 10713
rect 24030 10639 24086 10648
rect 24044 9761 24072 10639
rect 24228 10198 24256 11086
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10674 24716 10950
rect 24964 10674 24992 13806
rect 25056 11354 25084 23446
rect 25240 22778 25268 26959
rect 26252 24954 26280 27520
rect 26240 24948 26292 24954
rect 26240 24890 26292 24896
rect 27356 24410 27384 27520
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25608 22438 25636 23122
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25410 18728 25466 18737
rect 25410 18663 25466 18672
rect 25424 18426 25452 18663
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 25148 16726 25176 18090
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 25148 16250 25176 16662
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25134 16008 25190 16017
rect 25134 15943 25190 15952
rect 25148 15706 25176 15943
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25424 14006 25452 14418
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25516 13870 25544 21286
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25608 13530 25636 22374
rect 27618 17912 27674 17921
rect 27540 17882 27618 17898
rect 27528 17876 27618 17882
rect 27580 17870 27618 17876
rect 27618 17847 27674 17856
rect 27528 17818 27580 17824
rect 27618 13968 27674 13977
rect 27618 13903 27674 13912
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25792 12646 25820 13330
rect 27632 12889 27660 13903
rect 27618 12880 27674 12889
rect 27618 12815 27674 12824
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 24030 9752 24086 9761
rect 24030 9687 24086 9696
rect 24136 9586 24164 9930
rect 24228 9926 24256 10134
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24216 9920 24268 9926
rect 24216 9862 24268 9868
rect 24228 9722 24256 9862
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24044 8634 24072 8910
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 24136 7954 24164 9522
rect 24676 9444 24728 9450
rect 24676 9386 24728 9392
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24228 8022 24256 8910
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8022 24716 9386
rect 24780 9178 24808 9998
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24872 8838 24900 10406
rect 24964 9586 24992 10610
rect 25148 10470 25176 11154
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25148 10033 25176 10406
rect 25240 10062 25268 11494
rect 25228 10056 25280 10062
rect 25134 10024 25190 10033
rect 25228 9998 25280 10004
rect 25134 9959 25190 9968
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25042 8528 25098 8537
rect 25042 8463 25098 8472
rect 25056 8430 25084 8463
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 25042 7984 25098 7993
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24228 7410 24256 7958
rect 25240 7954 25268 8774
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25042 7919 25098 7928
rect 25228 7948 25280 7954
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24032 7268 24084 7274
rect 24032 7210 24084 7216
rect 24676 7268 24728 7274
rect 24676 7210 24728 7216
rect 24044 5914 24072 7210
rect 24216 6656 24268 6662
rect 24216 6598 24268 6604
rect 24228 6186 24256 6598
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6390 24716 7210
rect 25056 6866 25084 7919
rect 25228 7890 25280 7896
rect 25240 7546 25268 7890
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24124 5840 24176 5846
rect 24124 5782 24176 5788
rect 24136 5409 24164 5782
rect 24228 5778 24256 6122
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24122 5400 24178 5409
rect 24228 5370 24256 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24122 5335 24178 5344
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 23676 3738 23704 4150
rect 23860 4126 23980 4154
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23032 2854 23060 3130
rect 23860 3126 23888 4126
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22098 54 22324 82
rect 22834 82 22890 480
rect 23032 82 23060 2790
rect 22834 54 23060 82
rect 23400 82 23428 2994
rect 23662 82 23718 480
rect 23400 54 23718 82
rect 24044 82 24072 5102
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 24136 3602 24164 4694
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24228 3670 24256 4558
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 3738 24716 4966
rect 24780 4729 24808 6598
rect 25056 6458 25084 6802
rect 25332 6769 25360 7142
rect 25318 6760 25374 6769
rect 25318 6695 25374 6704
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24766 4720 24822 4729
rect 24766 4655 24822 4664
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24136 3194 24164 3538
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24228 3058 24256 3606
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 24688 2922 24716 3674
rect 24676 2916 24728 2922
rect 24676 2858 24728 2864
rect 24688 2582 24716 2858
rect 24676 2576 24728 2582
rect 24872 2553 24900 5034
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24964 3942 24992 4626
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24676 2518 24728 2524
rect 24858 2544 24914 2553
rect 24858 2479 24914 2488
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24398 82 24454 480
rect 24044 54 24454 82
rect 24964 82 24992 3878
rect 25056 3505 25084 6054
rect 25424 4282 25452 6666
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25700 4154 25728 8230
rect 25792 7274 25820 12582
rect 25870 12200 25926 12209
rect 25870 12135 25926 12144
rect 25884 7546 25912 12135
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25884 7342 25912 7482
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 27618 7304 27674 7313
rect 25780 7268 25832 7274
rect 27618 7239 27674 7248
rect 25780 7210 25832 7216
rect 27632 6361 27660 7239
rect 27618 6352 27674 6361
rect 27618 6287 27674 6296
rect 27252 6180 27304 6186
rect 27252 6122 27304 6128
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 25792 5098 25820 5714
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 25780 5092 25832 5098
rect 25780 5034 25832 5040
rect 25792 5001 25820 5034
rect 25778 4992 25834 5001
rect 25778 4927 25834 4936
rect 25700 4126 25820 4154
rect 25042 3496 25098 3505
rect 25042 3431 25098 3440
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25240 2417 25268 2790
rect 25226 2408 25282 2417
rect 25226 2343 25282 2352
rect 25226 82 25282 480
rect 24964 54 25282 82
rect 25792 82 25820 4126
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 26160 2310 26188 2450
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26160 1193 26188 2246
rect 26146 1184 26202 1193
rect 26146 1119 26202 1128
rect 25962 82 26018 480
rect 25792 54 26018 82
rect 26528 82 26556 5238
rect 26790 82 26846 480
rect 26528 54 26846 82
rect 27264 82 27292 6122
rect 27526 82 27582 480
rect 27264 54 27582 82
rect 20534 0 20590 54
rect 21362 0 21418 54
rect 22098 0 22154 54
rect 22834 0 22890 54
rect 23662 0 23718 54
rect 24398 0 24454 54
rect 25226 0 25282 54
rect 25962 0 26018 54
rect 26790 0 26846 54
rect 27526 0 27582 54
<< via2 >>
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 2410 19896 2466 19952
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 2686 17176 2742 17232
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 8850 20440 8906 20496
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 3974 13368 4030 13424
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5354 11056 5410 11112
rect 4710 6432 4766 6488
rect 5078 5072 5134 5128
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6458 10512 6514 10568
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5998 7384 6054 7440
rect 6366 7520 6422 7576
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10874 18672 10930 18728
rect 9126 15952 9182 16008
rect 7194 11192 7250 11248
rect 7010 10804 7066 10840
rect 7010 10784 7012 10804
rect 7012 10784 7064 10804
rect 7064 10784 7066 10804
rect 7102 10124 7158 10160
rect 7102 10104 7104 10124
rect 7104 10104 7156 10124
rect 7156 10104 7158 10124
rect 6090 6840 6146 6896
rect 5630 6704 5686 6760
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5998 6432 6054 6488
rect 6274 6160 6330 6216
rect 6274 5752 6330 5808
rect 5998 5616 6054 5672
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 3054 2352 3110 2408
rect 3974 1808 4030 1864
rect 4618 3032 4674 3088
rect 4986 2624 5042 2680
rect 5262 3712 5318 3768
rect 6366 5480 6422 5536
rect 6366 5344 6422 5400
rect 5998 4392 6054 4448
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5538 2488 5594 2544
rect 5446 1264 5502 1320
rect 5170 720 5226 776
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6366 1672 6422 1728
rect 6274 1128 6330 1184
rect 6642 4528 6698 4584
rect 7010 7928 7066 7984
rect 6918 7792 6974 7848
rect 6734 1944 6790 2000
rect 6918 3304 6974 3360
rect 7102 3440 7158 3496
rect 7470 5752 7526 5808
rect 7562 3984 7618 4040
rect 6826 584 6882 640
rect 8114 7656 8170 7712
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10782 17176 10838 17232
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 8390 2896 8446 2952
rect 9310 9424 9366 9480
rect 9402 6296 9458 6352
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9862 9968 9918 10024
rect 9770 9152 9826 9208
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 9126 3168 9182 3224
rect 9402 3612 9404 3632
rect 9404 3612 9456 3632
rect 9456 3612 9458 3632
rect 9402 3576 9458 3612
rect 10046 2624 10102 2680
rect 10414 5616 10470 5672
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10966 4936 11022 4992
rect 11978 12688 12034 12744
rect 13082 19896 13138 19952
rect 13358 19896 13414 19952
rect 12714 15408 12770 15464
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14830 20848 14886 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 12530 11056 12586 11112
rect 11610 6432 11666 6488
rect 13082 9152 13138 9208
rect 11794 4392 11850 4448
rect 12438 5480 12494 5536
rect 12162 3576 12218 3632
rect 12530 4392 12586 4448
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 16118 18128 16174 18184
rect 14462 12280 14518 12336
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15382 11192 15438 11248
rect 14554 10784 14610 10840
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15014 8064 15070 8120
rect 14646 7792 14702 7848
rect 14646 7520 14702 7576
rect 14002 6568 14058 6624
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 13358 4936 13414 4992
rect 12714 3576 12770 3632
rect 13450 3304 13506 3360
rect 14002 2896 14058 2952
rect 12070 2488 12126 2544
rect 13818 2352 13874 2408
rect 14186 2352 14242 2408
rect 14094 1672 14150 1728
rect 14554 1808 14610 1864
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 5888 15438 5944
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15382 4528 15438 4584
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19982 20440 20038 20496
rect 19062 19352 19118 19408
rect 19154 17584 19210 17640
rect 16486 13368 16542 13424
rect 16762 12280 16818 12336
rect 16210 9968 16266 10024
rect 16118 9696 16174 9752
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 18878 16088 18934 16144
rect 18786 15952 18842 16008
rect 17038 10920 17094 10976
rect 18418 11056 18474 11112
rect 18602 11056 18658 11112
rect 18694 10512 18750 10568
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20902 19896 20958 19952
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20810 18672 20866 18728
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 18786 10004 18788 10024
rect 18788 10004 18840 10024
rect 18840 10004 18842 10024
rect 18786 9968 18842 10004
rect 17774 6840 17830 6896
rect 17774 6724 17830 6760
rect 17774 6704 17776 6724
rect 17776 6704 17828 6724
rect 17828 6704 17830 6724
rect 17958 5208 18014 5264
rect 16486 3576 16542 3632
rect 16118 720 16174 776
rect 16486 1264 16542 1320
rect 18050 4664 18106 4720
rect 17130 1944 17186 2000
rect 16762 1128 16818 1184
rect 19062 9152 19118 9208
rect 19062 7792 19118 7848
rect 18694 7404 18750 7440
rect 18694 7384 18696 7404
rect 18696 7384 18748 7404
rect 18748 7384 18750 7404
rect 19062 6568 19118 6624
rect 18694 5344 18750 5400
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19890 8472 19946 8528
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19522 7928 19578 7984
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19338 6160 19394 6216
rect 18602 4936 18658 4992
rect 18418 2896 18474 2952
rect 22006 15408 22062 15464
rect 24766 25336 24822 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 25226 26968 25282 27024
rect 24858 23976 24914 24032
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22616 24822 22672
rect 23478 18128 23534 18184
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 21256 24822 21312
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20032 24822 20088
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24582 17584 24638 17640
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 23846 16088 23902 16144
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20994 6432 21050 6488
rect 19614 5208 19670 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 18878 3440 18934 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 18418 2488 18474 2544
rect 18326 584 18382 640
rect 22834 9424 22890 9480
rect 23018 5072 23074 5128
rect 22374 3576 22430 3632
rect 22926 3304 22982 3360
rect 24030 14592 24086 14648
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 23754 5208 23810 5264
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24030 12144 24086 12200
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24030 10920 24086 10976
rect 24030 10648 24086 10704
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 25410 18672 25466 18728
rect 25134 15952 25190 16008
rect 27618 17856 27674 17912
rect 27618 13912 27674 13968
rect 27618 12824 27674 12880
rect 24030 9696 24086 9752
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 25134 9968 25190 10024
rect 25042 8472 25098 8528
rect 25042 7928 25098 7984
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24122 5344 24178 5400
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25318 6704 25374 6760
rect 24766 4664 24822 4720
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24858 2488 24914 2544
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25870 12144 25926 12200
rect 27618 7248 27674 7304
rect 27618 6296 27674 6352
rect 25778 4936 25834 4992
rect 25042 3440 25098 3496
rect 25226 2352 25282 2408
rect 26146 1128 26202 1184
<< metal3 >>
rect 27520 27208 28000 27328
rect 25221 27026 25287 27029
rect 27662 27026 27722 27208
rect 25221 27024 27722 27026
rect 25221 26968 25226 27024
rect 25282 26968 27722 27024
rect 25221 26966 27722 26968
rect 25221 26963 25287 26966
rect 27520 25848 28000 25968
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25394 24827 25397
rect 27662 25394 27722 25848
rect 24761 25392 27722 25394
rect 24761 25336 24766 25392
rect 24822 25336 27722 25392
rect 24761 25334 27722 25336
rect 24761 25331 24827 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24608
rect 19610 24447 19930 24448
rect 24853 24034 24919 24037
rect 27662 24034 27722 24488
rect 24853 24032 27722 24034
rect 24853 23976 24858 24032
rect 24914 23976 27722 24032
rect 24853 23974 27722 23976
rect 24853 23971 24919 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 27520 23128 28000 23248
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 24761 22674 24827 22677
rect 27662 22674 27722 23128
rect 24761 22672 27722 22674
rect 24761 22616 24766 22672
rect 24822 22616 27722 22672
rect 24761 22614 27722 22616
rect 24761 22611 24827 22614
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21888
rect 24277 21727 24597 21728
rect 24761 21314 24827 21317
rect 27662 21314 27722 21768
rect 24761 21312 27722 21314
rect 24761 21256 24766 21312
rect 24822 21256 27722 21312
rect 24761 21254 27722 21256
rect 24761 21251 24827 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 14825 20906 14891 20909
rect 15510 20906 15516 20908
rect 14825 20904 15516 20906
rect 14825 20848 14830 20904
rect 14886 20848 15516 20904
rect 14825 20846 15516 20848
rect 14825 20843 14891 20846
rect 15510 20844 15516 20846
rect 15580 20844 15586 20908
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 27520 20544 28000 20664
rect 8845 20498 8911 20501
rect 19977 20498 20043 20501
rect 8845 20496 20043 20498
rect 8845 20440 8850 20496
rect 8906 20440 19982 20496
rect 20038 20440 20043 20496
rect 8845 20438 20043 20440
rect 8845 20435 8911 20438
rect 19977 20435 20043 20438
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 24761 20090 24827 20093
rect 27662 20090 27722 20544
rect 24761 20088 27722 20090
rect 24761 20032 24766 20088
rect 24822 20032 27722 20088
rect 24761 20030 27722 20032
rect 24761 20027 24827 20030
rect 2405 19954 2471 19957
rect 13077 19954 13143 19957
rect 2405 19952 13143 19954
rect 2405 19896 2410 19952
rect 2466 19896 13082 19952
rect 13138 19896 13143 19952
rect 2405 19894 13143 19896
rect 2405 19891 2471 19894
rect 13077 19891 13143 19894
rect 13353 19954 13419 19957
rect 20897 19954 20963 19957
rect 13353 19952 20963 19954
rect 13353 19896 13358 19952
rect 13414 19896 20902 19952
rect 20958 19896 20963 19952
rect 13353 19894 20963 19896
rect 13353 19891 13419 19894
rect 20897 19891 20963 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 15510 19348 15516 19412
rect 15580 19410 15586 19412
rect 19057 19410 19123 19413
rect 15580 19408 19123 19410
rect 15580 19352 19062 19408
rect 19118 19352 19123 19408
rect 15580 19350 19123 19352
rect 15580 19348 15586 19350
rect 19057 19347 19123 19350
rect 27520 19184 28000 19304
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 10869 18730 10935 18733
rect 20805 18730 20871 18733
rect 10869 18728 20871 18730
rect 10869 18672 10874 18728
rect 10930 18672 20810 18728
rect 20866 18672 20871 18728
rect 10869 18670 20871 18672
rect 10869 18667 10935 18670
rect 20805 18667 20871 18670
rect 25405 18730 25471 18733
rect 27662 18730 27722 19184
rect 25405 18728 27722 18730
rect 25405 18672 25410 18728
rect 25466 18672 27722 18728
rect 25405 18670 27722 18672
rect 25405 18667 25471 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 16113 18186 16179 18189
rect 23473 18186 23539 18189
rect 16113 18184 23539 18186
rect 16113 18128 16118 18184
rect 16174 18128 23478 18184
rect 23534 18128 23539 18184
rect 16113 18126 23539 18128
rect 16113 18123 16179 18126
rect 23473 18123 23539 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 27520 17912 28000 17944
rect 27520 17856 27618 17912
rect 27674 17856 28000 17912
rect 27520 17824 28000 17856
rect 19149 17642 19215 17645
rect 24577 17642 24643 17645
rect 19149 17640 24643 17642
rect 19149 17584 19154 17640
rect 19210 17584 24582 17640
rect 24638 17584 24643 17640
rect 19149 17582 24643 17584
rect 19149 17579 19215 17582
rect 24577 17579 24643 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 2681 17234 2747 17237
rect 10777 17234 10843 17237
rect 2681 17232 10843 17234
rect 2681 17176 2686 17232
rect 2742 17176 10782 17232
rect 10838 17176 10843 17232
rect 2681 17174 10843 17176
rect 2681 17171 2747 17174
rect 10777 17171 10843 17174
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 27520 16464 28000 16584
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 18873 16146 18939 16149
rect 23841 16146 23907 16149
rect 18873 16144 23907 16146
rect 18873 16088 18878 16144
rect 18934 16088 23846 16144
rect 23902 16088 23907 16144
rect 18873 16086 23907 16088
rect 18873 16083 18939 16086
rect 23841 16083 23907 16086
rect 9121 16010 9187 16013
rect 18781 16010 18847 16013
rect 9121 16008 18847 16010
rect 9121 15952 9126 16008
rect 9182 15952 18786 16008
rect 18842 15952 18847 16008
rect 9121 15950 18847 15952
rect 9121 15947 9187 15950
rect 18781 15947 18847 15950
rect 25129 16010 25195 16013
rect 27662 16010 27722 16464
rect 25129 16008 27722 16010
rect 25129 15952 25134 16008
rect 25190 15952 27722 16008
rect 25129 15950 27722 15952
rect 25129 15947 25195 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 12709 15466 12775 15469
rect 22001 15466 22067 15469
rect 12709 15464 22067 15466
rect 12709 15408 12714 15464
rect 12770 15408 22006 15464
rect 22062 15408 22067 15464
rect 12709 15406 22067 15408
rect 12709 15403 12775 15406
rect 22001 15403 22067 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 15104 28000 15224
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 24025 14650 24091 14653
rect 27662 14650 27722 15104
rect 24025 14648 27722 14650
rect 24025 14592 24030 14648
rect 24086 14592 27722 14648
rect 24025 14590 27722 14592
rect 24025 14587 24091 14590
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13968 28000 14000
rect 27520 13912 27618 13968
rect 27674 13912 28000 13968
rect 27520 13880 28000 13912
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3969 13426 4035 13429
rect 16481 13426 16547 13429
rect 3969 13424 16547 13426
rect 3969 13368 3974 13424
rect 4030 13368 16486 13424
rect 16542 13368 16547 13424
rect 3969 13366 16547 13368
rect 3969 13363 4035 13366
rect 16481 13363 16547 13366
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 27613 12882 27679 12885
rect 19290 12880 27679 12882
rect 19290 12824 27618 12880
rect 27674 12824 27679 12880
rect 19290 12822 27679 12824
rect 11973 12746 12039 12749
rect 19290 12746 19350 12822
rect 27613 12819 27679 12822
rect 11973 12744 19350 12746
rect 11973 12688 11978 12744
rect 12034 12688 19350 12744
rect 11973 12686 19350 12688
rect 11973 12683 12039 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12640
rect 19610 12479 19930 12480
rect 14457 12338 14523 12341
rect 16757 12338 16823 12341
rect 14457 12336 16823 12338
rect 14457 12280 14462 12336
rect 14518 12280 16762 12336
rect 16818 12280 16823 12336
rect 14457 12278 16823 12280
rect 14457 12275 14523 12278
rect 16757 12275 16823 12278
rect 24025 12202 24091 12205
rect 25865 12202 25931 12205
rect 27662 12202 27722 12520
rect 24025 12200 27722 12202
rect 24025 12144 24030 12200
rect 24086 12144 25870 12200
rect 25926 12144 27722 12200
rect 24025 12142 27722 12144
rect 24025 12139 24091 12142
rect 25865 12139 25931 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 7189 11250 7255 11253
rect 15377 11250 15443 11253
rect 7189 11248 15443 11250
rect 7189 11192 7194 11248
rect 7250 11192 15382 11248
rect 15438 11192 15443 11248
rect 7189 11190 15443 11192
rect 7189 11187 7255 11190
rect 15377 11187 15443 11190
rect 27520 11160 28000 11280
rect 5349 11114 5415 11117
rect 12525 11114 12591 11117
rect 18413 11114 18479 11117
rect 18597 11114 18663 11117
rect 5349 11112 18663 11114
rect 5349 11056 5354 11112
rect 5410 11056 12530 11112
rect 12586 11056 18418 11112
rect 18474 11056 18602 11112
rect 18658 11056 18663 11112
rect 5349 11054 18663 11056
rect 5349 11051 5415 11054
rect 12525 11051 12591 11054
rect 18413 11051 18479 11054
rect 18597 11051 18663 11054
rect 17033 10978 17099 10981
rect 24025 10978 24091 10981
rect 17033 10976 24091 10978
rect 17033 10920 17038 10976
rect 17094 10920 24030 10976
rect 24086 10920 24091 10976
rect 17033 10918 24091 10920
rect 17033 10915 17099 10918
rect 24025 10915 24091 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 7005 10842 7071 10845
rect 14549 10842 14615 10845
rect 7005 10840 14615 10842
rect 7005 10784 7010 10840
rect 7066 10784 14554 10840
rect 14610 10784 14615 10840
rect 7005 10782 14615 10784
rect 7005 10779 7071 10782
rect 14549 10779 14615 10782
rect 24025 10706 24091 10709
rect 27662 10706 27722 11160
rect 24025 10704 27722 10706
rect 24025 10648 24030 10704
rect 24086 10648 27722 10704
rect 24025 10646 27722 10648
rect 24025 10643 24091 10646
rect 6453 10570 6519 10573
rect 18689 10570 18755 10573
rect 6453 10568 18755 10570
rect 6453 10512 6458 10568
rect 6514 10512 18694 10568
rect 18750 10512 18755 10568
rect 6453 10510 18755 10512
rect 6453 10507 6519 10510
rect 18689 10507 18755 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 7097 10162 7163 10165
rect 7097 10160 27722 10162
rect 7097 10104 7102 10160
rect 7158 10104 27722 10160
rect 7097 10102 27722 10104
rect 7097 10099 7163 10102
rect 9857 10026 9923 10029
rect 16205 10026 16271 10029
rect 9857 10024 16271 10026
rect 9857 9968 9862 10024
rect 9918 9968 16210 10024
rect 16266 9968 16271 10024
rect 9857 9966 16271 9968
rect 9857 9963 9923 9966
rect 16205 9963 16271 9966
rect 18781 10026 18847 10029
rect 25129 10026 25195 10029
rect 18781 10024 25195 10026
rect 18781 9968 18786 10024
rect 18842 9968 25134 10024
rect 25190 9968 25195 10024
rect 18781 9966 25195 9968
rect 18781 9963 18847 9966
rect 25129 9963 25195 9966
rect 27662 9920 27722 10102
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 16113 9754 16179 9757
rect 24025 9754 24091 9757
rect 16113 9752 24091 9754
rect 16113 9696 16118 9752
rect 16174 9696 24030 9752
rect 24086 9696 24091 9752
rect 16113 9694 24091 9696
rect 16113 9691 16179 9694
rect 24025 9691 24091 9694
rect 9305 9482 9371 9485
rect 22829 9482 22895 9485
rect 9305 9480 22895 9482
rect 9305 9424 9310 9480
rect 9366 9424 22834 9480
rect 22890 9424 22895 9480
rect 9305 9422 22895 9424
rect 9305 9419 9371 9422
rect 22829 9419 22895 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 9765 9208 9831 9213
rect 9765 9152 9770 9208
rect 9826 9152 9831 9208
rect 9765 9147 9831 9152
rect 13077 9210 13143 9213
rect 19057 9210 19123 9213
rect 13077 9208 19123 9210
rect 13077 9152 13082 9208
rect 13138 9152 19062 9208
rect 19118 9152 19123 9208
rect 13077 9150 19123 9152
rect 13077 9147 13143 9150
rect 19057 9147 19123 9150
rect 9768 9076 9828 9147
rect 9768 9014 9812 9076
rect 9806 9012 9812 9014
rect 9876 9012 9882 9076
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 19885 8530 19951 8533
rect 25037 8530 25103 8533
rect 19885 8528 25103 8530
rect 19885 8472 19890 8528
rect 19946 8472 25042 8528
rect 25098 8472 25103 8528
rect 19885 8470 25103 8472
rect 19885 8467 19951 8470
rect 25037 8467 25103 8470
rect 27520 8440 28000 8560
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 14590 8060 14596 8124
rect 14660 8122 14666 8124
rect 15009 8122 15075 8125
rect 14660 8120 15075 8122
rect 14660 8064 15014 8120
rect 15070 8064 15075 8120
rect 14660 8062 15075 8064
rect 14660 8060 14666 8062
rect 15009 8059 15075 8062
rect 7005 7986 7071 7989
rect 19517 7986 19583 7989
rect 7005 7984 19583 7986
rect 7005 7928 7010 7984
rect 7066 7928 19522 7984
rect 19578 7928 19583 7984
rect 7005 7926 19583 7928
rect 7005 7923 7071 7926
rect 19517 7923 19583 7926
rect 25037 7986 25103 7989
rect 27662 7986 27722 8440
rect 25037 7984 27722 7986
rect 25037 7928 25042 7984
rect 25098 7928 27722 7984
rect 25037 7926 27722 7928
rect 25037 7923 25103 7926
rect 6913 7850 6979 7853
rect 14641 7850 14707 7853
rect 19057 7850 19123 7853
rect 6913 7848 14707 7850
rect 6913 7792 6918 7848
rect 6974 7792 14646 7848
rect 14702 7792 14707 7848
rect 6913 7790 14707 7792
rect 6913 7787 6979 7790
rect 14641 7787 14707 7790
rect 14782 7848 19123 7850
rect 14782 7792 19062 7848
rect 19118 7792 19123 7848
rect 14782 7790 19123 7792
rect 8109 7714 8175 7717
rect 14782 7714 14842 7790
rect 19057 7787 19123 7790
rect 8109 7712 14842 7714
rect 8109 7656 8114 7712
rect 8170 7656 14842 7712
rect 8109 7654 14842 7656
rect 8109 7651 8175 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6361 7578 6427 7581
rect 14641 7578 14707 7581
rect 6361 7576 14707 7578
rect 6361 7520 6366 7576
rect 6422 7520 14646 7576
rect 14702 7520 14707 7576
rect 6361 7518 14707 7520
rect 6361 7515 6427 7518
rect 14641 7515 14707 7518
rect 5993 7442 6059 7445
rect 18689 7442 18755 7445
rect 5993 7440 18755 7442
rect 5993 7384 5998 7440
rect 6054 7384 18694 7440
rect 18750 7384 18755 7440
rect 5993 7382 18755 7384
rect 5993 7379 6059 7382
rect 18689 7379 18755 7382
rect 27520 7304 28000 7336
rect 27520 7248 27618 7304
rect 27674 7248 28000 7304
rect 27520 7216 28000 7248
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 6085 6898 6151 6901
rect 17769 6898 17835 6901
rect 6085 6896 17835 6898
rect 6085 6840 6090 6896
rect 6146 6840 17774 6896
rect 17830 6840 17835 6896
rect 6085 6838 17835 6840
rect 6085 6835 6151 6838
rect 17769 6835 17835 6838
rect 5625 6762 5691 6765
rect 17769 6762 17835 6765
rect 25313 6762 25379 6765
rect 5625 6760 17602 6762
rect 5625 6704 5630 6760
rect 5686 6704 17602 6760
rect 5625 6702 17602 6704
rect 5625 6699 5691 6702
rect 9806 6564 9812 6628
rect 9876 6626 9882 6628
rect 13997 6626 14063 6629
rect 9876 6624 14063 6626
rect 9876 6568 14002 6624
rect 14058 6568 14063 6624
rect 9876 6566 14063 6568
rect 17542 6626 17602 6702
rect 17769 6760 25379 6762
rect 17769 6704 17774 6760
rect 17830 6704 25318 6760
rect 25374 6704 25379 6760
rect 17769 6702 25379 6704
rect 17769 6699 17835 6702
rect 25313 6699 25379 6702
rect 19057 6626 19123 6629
rect 17542 6624 19123 6626
rect 17542 6568 19062 6624
rect 19118 6568 19123 6624
rect 17542 6566 19123 6568
rect 9876 6564 9882 6566
rect 13997 6563 14063 6566
rect 19057 6563 19123 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 4705 6490 4771 6493
rect 4838 6490 4844 6492
rect 4705 6488 4844 6490
rect 4705 6432 4710 6488
rect 4766 6432 4844 6488
rect 4705 6430 4844 6432
rect 4705 6427 4771 6430
rect 4838 6428 4844 6430
rect 4908 6428 4914 6492
rect 5993 6490 6059 6493
rect 11605 6490 11671 6493
rect 5993 6488 11671 6490
rect 5993 6432 5998 6488
rect 6054 6432 11610 6488
rect 11666 6432 11671 6488
rect 5993 6430 11671 6432
rect 5993 6427 6059 6430
rect 11605 6427 11671 6430
rect 17350 6428 17356 6492
rect 17420 6490 17426 6492
rect 20989 6490 21055 6493
rect 17420 6488 21055 6490
rect 17420 6432 20994 6488
rect 21050 6432 21055 6488
rect 17420 6430 21055 6432
rect 17420 6428 17426 6430
rect 20989 6427 21055 6430
rect 9397 6354 9463 6357
rect 27613 6354 27679 6357
rect 9397 6352 27679 6354
rect 9397 6296 9402 6352
rect 9458 6296 27618 6352
rect 27674 6296 27679 6352
rect 9397 6294 27679 6296
rect 9397 6291 9463 6294
rect 27613 6291 27679 6294
rect 6269 6218 6335 6221
rect 19333 6218 19399 6221
rect 6269 6216 19399 6218
rect 6269 6160 6274 6216
rect 6330 6160 19338 6216
rect 19394 6160 19399 6216
rect 6269 6158 19399 6160
rect 6269 6155 6335 6158
rect 19333 6155 19399 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 15377 5946 15443 5949
rect 27520 5948 28000 5976
rect 15510 5946 15516 5948
rect 15377 5944 15516 5946
rect 15377 5888 15382 5944
rect 15438 5888 15516 5944
rect 15377 5886 15516 5888
rect 15377 5883 15443 5886
rect 15510 5884 15516 5886
rect 15580 5884 15586 5948
rect 27520 5884 27660 5948
rect 27724 5884 28000 5948
rect 27520 5856 28000 5884
rect 6269 5810 6335 5813
rect 7465 5810 7531 5813
rect 6269 5808 19350 5810
rect 6269 5752 6274 5808
rect 6330 5752 7470 5808
rect 7526 5752 19350 5808
rect 6269 5750 19350 5752
rect 6269 5747 6335 5750
rect 7465 5747 7531 5750
rect 5993 5674 6059 5677
rect 10409 5674 10475 5677
rect 5993 5672 10475 5674
rect 5993 5616 5998 5672
rect 6054 5616 10414 5672
rect 10470 5616 10475 5672
rect 5993 5614 10475 5616
rect 19290 5674 19350 5750
rect 27654 5674 27660 5676
rect 19290 5614 27660 5674
rect 5993 5611 6059 5614
rect 10409 5611 10475 5614
rect 27654 5612 27660 5614
rect 27724 5612 27730 5676
rect 6361 5538 6427 5541
rect 12433 5538 12499 5541
rect 6361 5536 12499 5538
rect 6361 5480 6366 5536
rect 6422 5480 12438 5536
rect 12494 5480 12499 5536
rect 6361 5478 12499 5480
rect 6361 5475 6427 5478
rect 12433 5475 12499 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 6361 5402 6427 5405
rect 6494 5402 6500 5404
rect 6361 5400 6500 5402
rect 6361 5344 6366 5400
rect 6422 5344 6500 5400
rect 6361 5342 6500 5344
rect 6361 5339 6427 5342
rect 6494 5340 6500 5342
rect 6564 5340 6570 5404
rect 18689 5402 18755 5405
rect 24117 5402 24183 5405
rect 18689 5400 24183 5402
rect 18689 5344 18694 5400
rect 18750 5344 24122 5400
rect 24178 5344 24183 5400
rect 18689 5342 24183 5344
rect 18689 5339 18755 5342
rect 24117 5339 24183 5342
rect 9622 5204 9628 5268
rect 9692 5266 9698 5268
rect 17953 5266 18019 5269
rect 9692 5264 18019 5266
rect 9692 5208 17958 5264
rect 18014 5208 18019 5264
rect 9692 5206 18019 5208
rect 9692 5204 9698 5206
rect 17953 5203 18019 5206
rect 19609 5266 19675 5269
rect 23749 5266 23815 5269
rect 19609 5264 23815 5266
rect 19609 5208 19614 5264
rect 19670 5208 23754 5264
rect 23810 5208 23815 5264
rect 19609 5206 23815 5208
rect 19609 5203 19675 5206
rect 23749 5203 23815 5206
rect 5073 5130 5139 5133
rect 23013 5130 23079 5133
rect 5073 5128 23079 5130
rect 5073 5072 5078 5128
rect 5134 5072 23018 5128
rect 23074 5072 23079 5128
rect 5073 5070 23079 5072
rect 5073 5067 5139 5070
rect 23013 5067 23079 5070
rect 10961 4994 11027 4997
rect 13353 4994 13419 4997
rect 18597 4994 18663 4997
rect 10961 4992 18663 4994
rect 10961 4936 10966 4992
rect 11022 4936 13358 4992
rect 13414 4936 18602 4992
rect 18658 4936 18663 4992
rect 10961 4934 18663 4936
rect 10961 4931 11027 4934
rect 13353 4931 13419 4934
rect 18597 4931 18663 4934
rect 25773 4994 25839 4997
rect 25773 4992 27722 4994
rect 25773 4936 25778 4992
rect 25834 4936 27722 4992
rect 25773 4934 27722 4936
rect 25773 4931 25839 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 18045 4722 18111 4725
rect 24761 4722 24827 4725
rect 18045 4720 24827 4722
rect 18045 4664 18050 4720
rect 18106 4664 24766 4720
rect 24822 4664 24827 4720
rect 18045 4662 24827 4664
rect 18045 4659 18111 4662
rect 24761 4659 24827 4662
rect 27662 4616 27722 4934
rect 6637 4586 6703 4589
rect 15377 4586 15443 4589
rect 6637 4584 15443 4586
rect 6637 4528 6642 4584
rect 6698 4528 15382 4584
rect 15438 4528 15443 4584
rect 6637 4526 15443 4528
rect 6637 4523 6703 4526
rect 15377 4523 15443 4526
rect 27520 4496 28000 4616
rect 5993 4450 6059 4453
rect 11789 4450 11855 4453
rect 12525 4450 12591 4453
rect 5993 4448 12591 4450
rect 5993 4392 5998 4448
rect 6054 4392 11794 4448
rect 11850 4392 12530 4448
rect 12586 4392 12591 4448
rect 5993 4390 12591 4392
rect 5993 4387 6059 4390
rect 11789 4387 11855 4390
rect 12525 4387 12591 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7557 4042 7623 4045
rect 9622 4042 9628 4044
rect 7557 4040 9628 4042
rect 7557 3984 7562 4040
rect 7618 3984 9628 4040
rect 7557 3982 9628 3984
rect 7557 3979 7623 3982
rect 9622 3980 9628 3982
rect 9692 3980 9698 4044
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 5257 3770 5323 3773
rect 9806 3770 9812 3772
rect 5257 3768 9812 3770
rect 5257 3712 5262 3768
rect 5318 3712 9812 3768
rect 5257 3710 9812 3712
rect 5257 3707 5323 3710
rect 9806 3708 9812 3710
rect 9876 3708 9882 3772
rect 9397 3634 9463 3637
rect 12157 3634 12223 3637
rect 9397 3632 12223 3634
rect 9397 3576 9402 3632
rect 9458 3576 12162 3632
rect 12218 3576 12223 3632
rect 9397 3574 12223 3576
rect 9397 3571 9463 3574
rect 12157 3571 12223 3574
rect 12709 3634 12775 3637
rect 16481 3634 16547 3637
rect 22369 3634 22435 3637
rect 12709 3632 13830 3634
rect 12709 3576 12714 3632
rect 12770 3576 13830 3632
rect 12709 3574 13830 3576
rect 12709 3571 12775 3574
rect 7097 3498 7163 3501
rect 12712 3498 12772 3571
rect 7097 3496 12772 3498
rect 7097 3440 7102 3496
rect 7158 3440 12772 3496
rect 7097 3438 12772 3440
rect 13770 3498 13830 3574
rect 16481 3632 22435 3634
rect 16481 3576 16486 3632
rect 16542 3576 22374 3632
rect 22430 3576 22435 3632
rect 16481 3574 22435 3576
rect 16481 3571 16547 3574
rect 22369 3571 22435 3574
rect 18873 3498 18939 3501
rect 25037 3498 25103 3501
rect 13770 3438 18706 3498
rect 7097 3435 7163 3438
rect 6913 3362 6979 3365
rect 13445 3362 13511 3365
rect 6913 3360 13511 3362
rect 6913 3304 6918 3360
rect 6974 3304 13450 3360
rect 13506 3304 13511 3360
rect 6913 3302 13511 3304
rect 18646 3362 18706 3438
rect 18873 3496 25103 3498
rect 18873 3440 18878 3496
rect 18934 3440 25042 3496
rect 25098 3440 25103 3496
rect 18873 3438 25103 3440
rect 18873 3435 18939 3438
rect 25037 3435 25103 3438
rect 22921 3362 22987 3365
rect 18646 3360 22987 3362
rect 18646 3304 22926 3360
rect 22982 3304 22987 3360
rect 18646 3302 22987 3304
rect 6913 3299 6979 3302
rect 13445 3299 13511 3302
rect 22921 3299 22987 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 9121 3226 9187 3229
rect 9254 3226 9260 3228
rect 7974 3224 9260 3226
rect 7974 3168 9126 3224
rect 9182 3168 9260 3224
rect 7974 3166 9260 3168
rect 4613 3090 4679 3093
rect 7974 3090 8034 3166
rect 9121 3163 9187 3166
rect 9254 3164 9260 3166
rect 9324 3164 9330 3228
rect 27520 3136 28000 3256
rect 4613 3088 8034 3090
rect 4613 3032 4618 3088
rect 4674 3032 8034 3088
rect 4613 3030 8034 3032
rect 4613 3027 4679 3030
rect 8385 2954 8451 2957
rect 13997 2954 14063 2957
rect 8385 2952 14063 2954
rect 8385 2896 8390 2952
rect 8446 2896 14002 2952
rect 14058 2896 14063 2952
rect 8385 2894 14063 2896
rect 8385 2891 8451 2894
rect 13997 2891 14063 2894
rect 18413 2954 18479 2957
rect 27662 2954 27722 3136
rect 18413 2952 27722 2954
rect 18413 2896 18418 2952
rect 18474 2896 27722 2952
rect 18413 2894 27722 2896
rect 18413 2891 18479 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4981 2682 5047 2685
rect 10041 2682 10107 2685
rect 4981 2680 10107 2682
rect 4981 2624 4986 2680
rect 5042 2624 10046 2680
rect 10102 2624 10107 2680
rect 4981 2622 10107 2624
rect 4981 2619 5047 2622
rect 10041 2619 10107 2622
rect 5533 2546 5599 2549
rect 12065 2546 12131 2549
rect 5533 2544 12131 2546
rect 5533 2488 5538 2544
rect 5594 2488 12070 2544
rect 12126 2488 12131 2544
rect 5533 2486 12131 2488
rect 5533 2483 5599 2486
rect 12065 2483 12131 2486
rect 18413 2546 18479 2549
rect 24853 2546 24919 2549
rect 18413 2544 24919 2546
rect 18413 2488 18418 2544
rect 18474 2488 24858 2544
rect 24914 2488 24919 2544
rect 18413 2486 24919 2488
rect 18413 2483 18479 2486
rect 24853 2483 24919 2486
rect 3049 2410 3115 2413
rect 13813 2410 13879 2413
rect 3049 2408 13879 2410
rect 3049 2352 3054 2408
rect 3110 2352 13818 2408
rect 13874 2352 13879 2408
rect 3049 2350 13879 2352
rect 3049 2347 3115 2350
rect 13813 2347 13879 2350
rect 14038 2348 14044 2412
rect 14108 2410 14114 2412
rect 14181 2410 14247 2413
rect 14108 2408 14247 2410
rect 14108 2352 14186 2408
rect 14242 2352 14247 2408
rect 14108 2350 14247 2352
rect 14108 2348 14114 2350
rect 14181 2347 14247 2350
rect 25221 2410 25287 2413
rect 25221 2408 27722 2410
rect 25221 2352 25226 2408
rect 25282 2352 27722 2408
rect 25221 2350 27722 2352
rect 25221 2347 25287 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6729 2002 6795 2005
rect 17125 2002 17191 2005
rect 6729 2000 17191 2002
rect 6729 1944 6734 2000
rect 6790 1944 17130 2000
rect 17186 1944 17191 2000
rect 6729 1942 17191 1944
rect 6729 1939 6795 1942
rect 17125 1939 17191 1942
rect 27662 1896 27722 2350
rect 3969 1866 4035 1869
rect 14549 1866 14615 1869
rect 3969 1864 14615 1866
rect 3969 1808 3974 1864
rect 4030 1808 14554 1864
rect 14610 1808 14615 1864
rect 3969 1806 14615 1808
rect 3969 1803 4035 1806
rect 14549 1803 14615 1806
rect 27520 1776 28000 1896
rect 6361 1730 6427 1733
rect 14089 1730 14155 1733
rect 6361 1728 14155 1730
rect 6361 1672 6366 1728
rect 6422 1672 14094 1728
rect 14150 1672 14155 1728
rect 6361 1670 14155 1672
rect 6361 1667 6427 1670
rect 14089 1667 14155 1670
rect 5441 1322 5507 1325
rect 16481 1322 16547 1325
rect 5441 1320 16547 1322
rect 5441 1264 5446 1320
rect 5502 1264 16486 1320
rect 16542 1264 16547 1320
rect 5441 1262 16547 1264
rect 5441 1259 5507 1262
rect 16481 1259 16547 1262
rect 6269 1186 6335 1189
rect 16757 1186 16823 1189
rect 6269 1184 16823 1186
rect 6269 1128 6274 1184
rect 6330 1128 16762 1184
rect 16818 1128 16823 1184
rect 6269 1126 16823 1128
rect 6269 1123 6335 1126
rect 16757 1123 16823 1126
rect 26141 1186 26207 1189
rect 26141 1184 27722 1186
rect 26141 1128 26146 1184
rect 26202 1128 27722 1184
rect 26141 1126 27722 1128
rect 26141 1123 26207 1126
rect 5165 778 5231 781
rect 16113 778 16179 781
rect 5165 776 16179 778
rect 5165 720 5170 776
rect 5226 720 16118 776
rect 16174 720 16179 776
rect 5165 718 16179 720
rect 5165 715 5231 718
rect 16113 715 16179 718
rect 27662 672 27722 1126
rect 6821 642 6887 645
rect 18321 642 18387 645
rect 6821 640 18387 642
rect 6821 584 6826 640
rect 6882 584 18326 640
rect 18382 584 18387 640
rect 6821 582 18387 584
rect 6821 579 6887 582
rect 18321 579 18387 582
rect 27520 552 28000 672
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 15516 20844 15580 20908
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 15516 19348 15580 19412
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 9812 9012 9876 9076
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 14596 8060 14660 8124
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 9812 6564 9876 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 4844 6428 4908 6492
rect 17356 6428 17420 6492
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 15516 5884 15580 5948
rect 27660 5884 27724 5948
rect 27660 5612 27724 5676
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 6500 5340 6564 5404
rect 9628 5204 9692 5268
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 9628 3980 9692 4044
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 9812 3708 9876 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 9260 3164 9324 3228
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 14044 2348 14108 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 9811 9076 9877 9077
rect 9811 9012 9812 9076
rect 9876 9012 9877 9076
rect 9811 9011 9877 9012
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 9814 6629 9874 9011
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 15515 20908 15581 20909
rect 15515 20844 15516 20908
rect 15580 20844 15581 20908
rect 15515 20843 15581 20844
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 15518 19413 15578 20843
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 15515 19412 15581 19413
rect 15515 19348 15516 19412
rect 15580 19348 15581 19412
rect 15515 19347 15581 19348
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14595 8124 14661 8125
rect 14595 8060 14596 8124
rect 14660 8060 14661 8124
rect 14595 8059 14661 8060
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 9811 6628 9877 6629
rect 9811 6564 9812 6628
rect 9876 6564 9877 6628
rect 9811 6563 9877 6564
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 6499 5404 6565 5405
rect 6499 5340 6500 5404
rect 6564 5340 6565 5404
rect 6499 5339 6565 5340
rect 6502 5218 6562 5339
rect 9627 5268 9693 5269
rect 9627 5204 9628 5268
rect 9692 5204 9693 5268
rect 9627 5203 9693 5204
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 9630 4045 9690 5203
rect 9627 4044 9693 4045
rect 9627 3980 9628 4044
rect 9692 3980 9693 4044
rect 9627 3979 9693 3980
rect 9814 3773 9874 6563
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 14598 5218 14658 8059
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 15518 5949 15578 19347
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 15515 5948 15581 5949
rect 15515 5884 15516 5948
rect 15580 5884 15581 5948
rect 15515 5883 15581 5884
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 9811 3772 9877 3773
rect 9811 3708 9812 3772
rect 9876 3708 9877 3772
rect 9811 3707 9877 3708
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 9259 3228 9325 3229
rect 9259 3164 9260 3228
rect 9324 3164 9325 3228
rect 9259 3163 9325 3164
rect 9262 2498 9322 3163
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2128 10597 2688
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 27659 5948 27725 5949
rect 27659 5884 27660 5948
rect 27724 5884 27725 5948
rect 27659 5883 27725 5884
rect 27662 5677 27722 5883
rect 27659 5676 27725 5677
rect 27659 5612 27660 5676
rect 27724 5612 27725 5676
rect 27659 5611 27725 5612
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 4758 6492 4994 6578
rect 4758 6428 4844 6492
rect 4844 6428 4908 6492
rect 4908 6428 4994 6492
rect 4758 6342 4994 6428
rect 6414 4982 6650 5218
rect 17270 6492 17506 6578
rect 17270 6428 17356 6492
rect 17356 6428 17420 6492
rect 17420 6428 17506 6492
rect 17270 6342 17506 6428
rect 14510 4982 14746 5218
rect 9174 2262 9410 2498
rect 13958 2412 14194 2498
rect 13958 2348 14044 2412
rect 14044 2348 14108 2412
rect 14108 2348 14194 2412
rect 13958 2262 14194 2348
<< metal5 >>
rect 4716 6578 17548 6620
rect 4716 6342 4758 6578
rect 4994 6342 17270 6578
rect 17506 6342 17548 6578
rect 4716 6300 17548 6342
rect 6372 5218 14788 5260
rect 6372 4982 6414 5218
rect 6650 4982 14510 5218
rect 14746 4982 14788 5218
rect 6372 4940 14788 4982
rect 9132 2498 14236 2540
rect 9132 2262 9174 2498
rect 9410 2262 13958 2498
rect 14194 2262 14236 2498
rect 9132 2220 14236 2262
use scs8hd_decap_8  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_17
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_12
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_22 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_46
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use scs8hd_conb_1  _189_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_60
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _217_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 -1 2720
box -38 -48 406 592
use scs8hd_nor2_4  _139_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _216_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_177
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_173
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_181
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_200
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_1  _100_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _076_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_or3_4  _093_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_263 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_231
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 130 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use scs8hd_or3_4  _135_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_247
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_49
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6900 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_72
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_213
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _077_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 406 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_265
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_103
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_169
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_177
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_240
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_244
timestamp 1586364061
transform 1 0 23552 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_25
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_29
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_37
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_76
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_91
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_155
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 130 592
use scs8hd_or3_4  _096_
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__C
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_205
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_222
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 314 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_18
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_40
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_124
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _214_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_185
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_198
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_nor4_4  _172_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 1602 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_or3_4  _081_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_229
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_235
timestamp 1586364061
transform 1 0 22724 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_242
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_243
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 23552 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_257
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_253
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_265
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_261
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_264
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_48
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _215_
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_169
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_nor4_4  _171_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_255
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_262
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 406 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_190
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_256
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_267
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_271
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_121
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 15364 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_146
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_164
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_185
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_198
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _082_
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 22356 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_222
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_229
timestamp 1586364061
transform 1 0 22172 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_6  FILLER_10_233
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_248
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_252
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_45
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_72
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_76
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_129
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 406 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 866 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_206
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_1  _147_
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_or3_4  _146_
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_188
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _167_
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23368 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 25116 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_257
timestamp 1586364061
transform 1 0 24748 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_264
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_126
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_150
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_184
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _125_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 1050 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_244
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_249
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_262
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _117_
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_212
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 314 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_242
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_260
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _118_
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_118
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 590 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1602 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23000 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_232
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_249
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_253
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_260
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_272
timestamp 1586364061
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_76
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 406 592
use scs8hd_nor4_4  _169_
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 1602 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_238
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_265
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_165
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_250
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_254
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 590 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 866 592
use scs8hd_conb_1  _198_
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_189
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_205
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_209
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__D
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__D
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 1602 592
use scs8hd_nor4_4  _159_
timestamp 1586364061
transform 1 0 21436 0 -1 13600
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_238
timestamp 1586364061
transform 1 0 23000 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _196_
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_255
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_255
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_70
timestamp 1586364061
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_133
timestamp 1586364061
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_188
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_192
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 314 592
use scs8hd_nor4_4  _165_
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 1602 592
use scs8hd_decap_4  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_224
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_231
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_235
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_249
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_265
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_273
timestamp 1586364061
transform 1 0 26220 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_73
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_76
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _199_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_148
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_151
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_176
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_193
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 19596 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _157_
timestamp 1586364061
transform 1 0 21528 0 -1 14688
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_243
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _160_
timestamp 1586364061
transform 1 0 25392 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_256
timestamp 1586364061
transform 1 0 24656 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_267
timestamp 1586364061
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 314 592
use scs8hd_nor4_4  _164_
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_230
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_256
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_261
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_267
timestamp 1586364061
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_271
timestamp 1586364061
transform 1 0 26036 0 1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_72
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_96
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_100
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_103
timestamp 1586364061
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _161_
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_181
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_24_232
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_255
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_70
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 774 592
use scs8hd_conb_1  _197_
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_131
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_169
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_190
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_194
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _162_
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_223
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_146
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_201
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__D
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_203
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_207
timestamp 1586364061
transform 1 0 20148 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_211
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_226
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_230
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_230
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_245
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 866 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 25484 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_250
timestamp 1586364061
transform 1 0 24104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_262
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_261
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_268
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_209
timestamp 1586364061
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_230
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 406 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_164
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16008 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_182
timestamp 1586364061
transform 1 0 17848 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_189
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23184 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_243
timestamp 1586364061
transform 1 0 23460 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_266
timestamp 1586364061
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_200
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_218
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_231
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_235
timestamp 1586364061
transform 1 0 22724 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_243
timestamp 1586364061
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_249
timestamp 1586364061
transform 1 0 24012 0 1 19040
box -38 -48 590 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_259
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_263
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_275
timestamp 1586364061
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_165
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_177
timestamp 1586364061
transform 1 0 17388 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_189
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_197
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_6  FILLER_32_207
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_224
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_235
timestamp 1586364061
transform 1 0 22724 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_243
timestamp 1586364061
transform 1 0 23460 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_247
timestamp 1586364061
transform 1 0 23828 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_259
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 314 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_213
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_229
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_218
timestamp 1586364061
transform 1 0 21160 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_230
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_241
timestamp 1586364061
transform 1 0 23276 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_242
timestamp 1586364061
transform 1 0 23368 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_259
timestamp 1586364061
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_263
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_254
timestamp 1586364061
transform 1 0 24472 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_266
timestamp 1586364061
transform 1 0 25576 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_275
timestamp 1586364061
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25392 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_262
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_17
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_28
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_44
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_60
timestamp 1586364061
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_56
timestamp 1586364061
transform 1 0 6256 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_71
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_81
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_85
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_83
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_126
timestamp 1586364061
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_186
timestamp 1586364061
transform 1 0 18216 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 18216 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_194
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_190
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_198
timestamp 1586364061
transform 1 0 19320 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_212
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_224
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_243
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _218_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 590 592
use scs8hd_buf_2  _219_
timestamp 1586364061
transform 1 0 24288 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_251
timestamp 1586364061
transform 1 0 24196 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_256
timestamp 1586364061
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_260
timestamp 1586364061
transform 1 0 25024 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_41_272
timestamp 1586364061
transform 1 0 26128 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_276
timestamp 1586364061
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 22098 0 22154 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 22834 0 22890 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 23662 0 23718 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 24398 0 24454 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 25226 0 25282 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 25962 0 26018 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 26790 0 26846 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 4250 0 4306 480 6 bottom_left_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 4986 0 5042 480 6 bottom_left_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 5814 0 5870 480 6 bottom_left_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 386 0 442 480 6 bottom_left_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 1858 0 1914 480 6 bottom_left_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 2686 0 2742 480 6 bottom_left_grid_pin_7_
port 13 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_9_
port 14 nsew default input
rlabel metal2 s 20534 0 20590 480 6 bottom_right_grid_pin_11_
port 15 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[0]
port 16 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal3 s 27520 5856 28000 5976 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal3 s 27520 16464 28000 16584 6 chanx_right_out[1]
port 26 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chanx_right_out[2]
port 27 nsew default tristate
rlabel metal3 s 27520 19184 28000 19304 6 chanx_right_out[3]
port 28 nsew default tristate
rlabel metal3 s 27520 20544 28000 20664 6 chanx_right_out[4]
port 29 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[5]
port 30 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[6]
port 31 nsew default tristate
rlabel metal3 s 27520 24488 28000 24608 6 chanx_right_out[7]
port 32 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[8]
port 33 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 14462 27520 14518 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 15474 27520 15530 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 17682 27520 17738 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 19798 27520 19854 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 25134 27520 25190 28000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 26238 27520 26294 28000 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 27342 27520 27398 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 data_in
port 70 nsew default input
rlabel metal2 s 21362 0 21418 480 6 enable
port 71 nsew default input
rlabel metal3 s 27520 27208 28000 27328 6 right_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 27520 1776 28000 1896 6 right_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 5814 27520 5870 28000 6 top_left_grid_pin_11_
port 74 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 top_left_grid_pin_13_
port 75 nsew default input
rlabel metal2 s 7930 27520 7986 28000 6 top_left_grid_pin_15_
port 76 nsew default input
rlabel metal2 s 478 27520 534 28000 6 top_left_grid_pin_1_
port 77 nsew default input
rlabel metal2 s 1490 27520 1546 28000 6 top_left_grid_pin_3_
port 78 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_5_
port 79 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_7_
port 80 nsew default input
rlabel metal2 s 4710 27520 4766 28000 6 top_left_grid_pin_9_
port 81 nsew default input
rlabel metal3 s 27520 552 28000 672 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
