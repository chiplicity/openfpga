VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_left
  CLASS BLOCK ;
  FOREIGN grid_io_left ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 139.440 80.000 140.040 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 197.600 20.150 200.000 ;
    END
  END ccff_tail
  PIN gfpga_pad_GPIO_A
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 197.600 60.170 200.000 ;
    END
  END gfpga_pad_GPIO_A
  PIN gfpga_pad_GPIO_IE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 179.560 80.000 180.160 ;
    END
  END gfpga_pad_GPIO_IE
  PIN gfpga_pad_GPIO_OE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END gfpga_pad_GPIO_OE
  PIN gfpga_pad_GPIO_Y
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END gfpga_pad_GPIO_Y
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 19.760 80.000 20.360 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 59.200 80.000 59.800 ;
    END
  END right_width_0_height_0__pin_1_lower
  PIN right_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 99.320 80.000 99.920 ;
    END
  END right_width_0_height_0__pin_1_upper
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 74.060 187.920 ;
      LAYER met2 ;
        RECT 13.890 197.320 19.590 197.610 ;
        RECT 20.430 197.320 59.610 197.610 ;
        RECT 60.450 197.320 72.925 197.610 ;
        RECT 13.890 2.680 72.925 197.320 ;
        RECT 13.890 2.400 19.590 2.680 ;
        RECT 20.430 2.400 59.610 2.680 ;
        RECT 60.450 2.400 72.925 2.680 ;
      LAYER met3 ;
        RECT 2.400 180.560 77.600 187.845 ;
        RECT 2.400 179.160 77.200 180.560 ;
        RECT 2.400 140.440 77.600 179.160 ;
        RECT 2.400 139.040 77.200 140.440 ;
        RECT 2.400 101.000 77.600 139.040 ;
        RECT 2.800 100.320 77.600 101.000 ;
        RECT 2.800 99.600 77.200 100.320 ;
        RECT 2.400 98.920 77.200 99.600 ;
        RECT 2.400 60.200 77.600 98.920 ;
        RECT 2.400 58.800 77.200 60.200 ;
        RECT 2.400 20.760 77.600 58.800 ;
        RECT 2.400 19.360 77.200 20.760 ;
        RECT 2.400 10.715 77.600 19.360 ;
      LAYER met4 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END grid_io_left
END LIBRARY

