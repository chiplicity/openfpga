magic
tech EFS8A
magscale 1 2
timestamp 1602096022
<< locali >>
rect 29 17459 63 22457
rect 29 11339 63 17289
rect 121 13719 155 18309
rect 121 9027 155 13345
rect 213 10387 247 17017
rect 121 8993 247 9027
rect 121 119 155 8925
rect 213 6851 247 8993
rect 305 6647 339 17493
rect 397 10523 431 16541
rect 489 14467 523 22389
rect 581 14739 615 23205
rect 673 16779 707 19193
rect 397 9843 431 10353
rect 489 9843 523 13549
rect 581 9843 615 14569
rect 673 9911 707 15929
rect 765 13515 799 19125
rect 857 16031 891 21641
rect 949 17867 983 23069
rect 6101 22423 6135 22525
rect 5089 21879 5123 22389
rect 6193 22287 6227 22525
rect 6285 22287 6319 22593
rect 7389 22151 7423 23001
rect 7757 22015 7791 23069
rect 8033 22083 8067 22865
rect 8861 22627 8895 23205
rect 8953 22899 8987 23545
rect 9045 22219 9079 22933
rect 11069 22151 11103 22321
rect 2145 21471 2179 21641
rect 1443 21437 1478 21471
rect 6871 21437 6951 21471
rect 16681 21335 16715 21641
rect 8585 20927 8619 20961
rect 8401 20893 8619 20927
rect 8769 19873 8953 19907
rect 6009 19227 6043 19397
rect 6285 19159 6319 19397
rect 9229 19295 9263 19465
rect 13645 19363 13679 19465
rect 12265 19261 12449 19295
rect 7665 19159 7699 19261
rect 11529 19159 11563 19261
rect 8803 19125 8987 19159
rect 13737 19023 13771 19261
rect 14749 19193 14875 19227
rect 14841 19159 14875 19193
rect 13737 18989 13863 19023
rect 9597 18411 9631 18785
rect 13829 18615 13863 18989
rect 18371 18785 18498 18819
rect 19475 18785 19510 18819
rect 13829 18581 13921 18615
rect 5641 18207 5675 18377
rect 14841 18207 14875 18377
rect 6469 18071 6503 18173
rect 16405 18071 16439 18173
rect 6285 17527 6319 17833
rect 14105 17527 14139 17629
rect 18245 17595 18279 17697
rect 3341 17051 3375 17289
rect 4445 16983 4479 17289
rect 9965 16983 9999 17289
rect 13645 16983 13679 17153
rect 13737 17119 13771 17289
rect 16773 17051 16807 17289
rect 857 13583 891 15589
rect 397 9809 707 9843
rect 397 4157 431 9741
rect 489 4471 523 9809
rect 581 8483 615 9809
rect 673 6715 707 9809
rect 765 5559 799 13209
rect 857 5015 891 13413
rect 949 12427 983 16677
rect 3433 15351 3467 16201
rect 3525 15895 3559 16201
rect 15209 15895 15243 16133
rect 4491 15657 4629 15691
rect 5457 15487 5491 15657
rect 6193 15521 6411 15555
rect 6193 15419 6227 15521
rect 2145 13719 2179 15113
rect 12725 14807 12759 15521
rect 14933 15419 14967 15657
rect 14749 14807 14783 15113
rect 16313 14943 16347 15113
rect 16405 14875 16439 15113
rect 12811 14569 12817 14603
rect 3617 14263 3651 14433
rect 3893 14331 3927 14569
rect 12811 14501 12845 14569
rect 4077 14467 4111 14501
rect 4077 14433 4330 14467
rect 3614 14229 3651 14263
rect 3614 14059 3648 14229
rect 3614 14025 3651 14059
rect 3617 13787 3651 14025
rect 4445 13719 4479 13957
rect 6377 13719 6411 14501
rect 6469 13719 6503 13957
rect 9597 13719 9631 14025
rect 16399 13515 16433 13787
rect 16399 13481 16439 13515
rect 1041 13175 1075 13481
rect 16405 13447 16439 13481
rect 16037 13175 16071 13413
rect 16589 12937 16681 12971
rect 1547 12801 1685 12835
rect 10517 12427 10551 12597
rect 10511 12393 10551 12427
rect 949 10591 983 12393
rect 10511 12325 10545 12393
rect 6929 12257 7113 12291
rect 14473 12087 14507 12257
rect 8217 11543 8251 11577
rect 8211 11509 8251 11543
rect 7113 10999 7147 11305
rect 8211 11237 8245 11509
rect 16123 11305 16129 11339
rect 16123 11237 16157 11305
rect 14139 11169 14174 11203
rect 17543 11169 17578 11203
rect 5175 10455 5209 10523
rect 5175 10421 5181 10455
rect 7751 10421 7883 10455
rect 1777 10251 1811 10421
rect 7751 10251 7785 10421
rect 1771 10217 1777 10251
rect 1771 10168 1811 10217
rect 1771 10149 1805 10168
rect 4169 9503 4203 10217
rect 7751 10149 7785 10217
rect 6101 9367 6135 9605
rect 7665 9367 7699 9673
rect 4203 9333 4295 9367
rect 8401 9367 8435 10557
rect 9631 10081 9758 10115
rect 10333 9979 10367 10149
rect 10735 10081 10770 10115
rect 11529 9367 11563 9469
rect 11989 9367 12023 10081
rect 17831 9877 17969 9911
rect 15393 9503 15427 9605
rect 14743 9367 14777 9435
rect 14743 9333 14749 9367
rect 4260 9299 4294 9333
rect 4260 9265 4295 9299
rect 4261 9231 4295 9265
rect 4260 9197 4295 9231
rect 4260 9163 4294 9197
rect 4169 9129 4294 9163
rect 397 4123 615 4157
rect 581 2635 615 4123
rect 949 3179 983 8857
rect 4169 8823 4203 9129
rect 5031 9061 5076 9095
rect 6101 8823 6135 9333
rect 8401 8823 8435 9333
rect 10425 8823 10459 9129
rect 11247 9129 11253 9163
rect 11247 9061 11281 9129
rect 19751 8993 19786 9027
rect 8401 8789 8769 8823
rect 6101 8619 6135 8789
rect 1443 8381 1478 8415
rect 3433 8279 3467 8585
rect 5089 8075 5123 8517
rect 7941 8279 7975 8381
rect 9137 8075 9171 8381
rect 5083 8041 5123 8075
rect 9137 8041 9263 8075
rect 5083 8007 5117 8041
rect 9137 7735 9171 8041
rect 13093 7735 13127 7973
rect 17509 7871 17543 7973
rect 1547 7701 1639 7735
rect 6193 7667 6227 7701
rect 6193 7633 6319 7667
rect 5583 7497 5675 7531
rect 2605 7191 2639 7497
rect 5641 7259 5675 7497
rect 6285 7191 6319 7633
rect 8309 7327 8343 7497
rect 9597 7327 9631 7497
rect 10241 7191 10275 7497
rect 13921 7327 13955 7497
rect 8211 6953 8217 6987
rect 12167 6953 12173 6987
rect 4077 6647 4111 6953
rect 8211 6885 8245 6953
rect 12167 6885 12201 6953
rect 6745 6715 6779 6885
rect 9321 6647 9355 6817
rect 1719 6205 1754 6239
rect 12817 6171 12851 6409
rect 19257 6103 19291 6341
rect 3283 5729 3318 5763
rect 8619 5729 8654 5763
rect 9229 5695 9263 5865
rect 9321 5559 9355 5797
rect 14013 5151 14047 5321
rect 15519 5117 15611 5151
rect 16899 5117 16934 5151
rect 1771 5015 1805 5083
rect 2783 5015 2817 5083
rect 8211 5015 8245 5083
rect 14013 5015 14047 5117
rect 1771 4981 1811 5015
rect 2783 4981 2789 5015
rect 8211 4981 8217 5015
rect 15577 5015 15611 5117
rect 1777 4811 1811 4981
rect 18337 4811 18371 5049
rect 1771 4777 1777 4811
rect 18331 4777 18371 4811
rect 1771 4709 1805 4777
rect 3571 4709 3652 4743
rect 18331 4709 18365 4777
rect 3467 4641 3502 4675
rect 16037 4471 16071 4573
rect 21741 4471 21775 4641
rect 6135 4233 6181 4267
rect 4905 3995 4939 4233
rect 19257 3995 19291 4165
rect 1863 3927 1897 3995
rect 5359 3927 5393 3995
rect 1863 3893 1869 3927
rect 5359 3893 5365 3927
rect 1771 3689 1777 3723
rect 4531 3689 4537 3723
rect 10787 3689 10793 3723
rect 1771 3621 1805 3689
rect 4531 3621 4565 3689
rect 10787 3621 10821 3689
rect 9171 3553 9206 3587
rect 16497 3519 16531 3621
rect 4077 3485 4199 3519
rect 4077 3451 4111 3485
rect 17877 3383 17911 3689
rect 6503 2941 6538 2975
rect 12115 2941 12150 2975
rect 1771 2839 1805 2907
rect 2783 2839 2817 2907
rect 5767 2873 5812 2907
rect 1771 2805 1777 2839
rect 2783 2805 2789 2839
rect 17049 2295 17083 2397
rect 14335 2261 14473 2295
rect 19533 2295 19567 2397
<< viali >>
rect 8953 23545 8987 23579
rect 581 23205 615 23239
rect 29 22457 63 22491
rect 489 22389 523 22423
rect 29 17425 63 17459
rect 121 18309 155 18343
rect 29 17289 63 17323
rect 305 17493 339 17527
rect 121 13685 155 13719
rect 213 17017 247 17051
rect 29 11305 63 11339
rect 121 13345 155 13379
rect 213 10353 247 10387
rect 121 8925 155 8959
rect 213 6817 247 6851
rect 397 16541 431 16575
rect 8861 23205 8895 23239
rect 949 23069 983 23103
rect 857 21641 891 21675
rect 673 19193 707 19227
rect 673 16745 707 16779
rect 765 19125 799 19159
rect 581 14705 615 14739
rect 673 15929 707 15963
rect 489 14433 523 14467
rect 581 14569 615 14603
rect 397 10489 431 10523
rect 489 13549 523 13583
rect 397 10353 431 10387
rect 7757 23069 7791 23103
rect 7389 23001 7423 23035
rect 6285 22593 6319 22627
rect 6101 22525 6135 22559
rect 5089 22389 5123 22423
rect 6101 22389 6135 22423
rect 6193 22525 6227 22559
rect 6193 22253 6227 22287
rect 6285 22253 6319 22287
rect 7389 22117 7423 22151
rect 8033 22865 8067 22899
rect 8953 22865 8987 22899
rect 9045 22933 9079 22967
rect 8861 22593 8895 22627
rect 9045 22185 9079 22219
rect 11069 22321 11103 22355
rect 11069 22117 11103 22151
rect 8033 22049 8067 22083
rect 7757 21981 7791 22015
rect 5089 21845 5123 21879
rect 2145 21641 2179 21675
rect 2237 21641 2271 21675
rect 3893 21641 3927 21675
rect 9597 21641 9631 21675
rect 13645 21641 13679 21675
rect 14473 21641 14507 21675
rect 16497 21641 16531 21675
rect 16681 21641 16715 21675
rect 18502 21641 18536 21675
rect 19349 21641 19383 21675
rect 1961 21505 1995 21539
rect 4242 21573 4276 21607
rect 4353 21573 4387 21607
rect 6377 21573 6411 21607
rect 11575 21573 11609 21607
rect 13277 21573 13311 21607
rect 16129 21573 16163 21607
rect 2513 21505 2547 21539
rect 4445 21505 4479 21539
rect 6745 21505 6779 21539
rect 7021 21505 7055 21539
rect 1409 21437 1443 21471
rect 2145 21437 2179 21471
rect 2421 21437 2455 21471
rect 2697 21437 2731 21471
rect 4077 21437 4111 21471
rect 5676 21437 5710 21471
rect 6837 21437 6871 21471
rect 7205 21437 7239 21471
rect 7665 21437 7699 21471
rect 8712 21437 8746 21471
rect 9137 21437 9171 21471
rect 10057 21437 10091 21471
rect 10333 21437 10367 21471
rect 11472 21437 11506 21471
rect 11897 21437 11931 21471
rect 14289 21437 14323 21471
rect 3157 21369 3191 21403
rect 8309 21369 8343 21403
rect 8815 21369 8849 21403
rect 12357 21369 12391 21403
rect 12725 21369 12759 21403
rect 12817 21369 12851 21403
rect 15209 21369 15243 21403
rect 15577 21369 15611 21403
rect 15669 21369 15703 21403
rect 18613 21573 18647 21607
rect 18705 21505 18739 21539
rect 21327 21505 21361 21539
rect 17084 21437 17118 21471
rect 17785 21437 17819 21471
rect 19936 21437 19970 21471
rect 20361 21437 20395 21471
rect 21224 21437 21258 21471
rect 21649 21437 21683 21471
rect 17187 21369 17221 21403
rect 18337 21369 18371 21403
rect 19717 21369 19751 21403
rect 1547 21301 1581 21335
rect 3433 21301 3467 21335
rect 4721 21301 4755 21335
rect 5089 21301 5123 21335
rect 5457 21301 5491 21335
rect 5779 21301 5813 21335
rect 8033 21301 8067 21335
rect 9873 21301 9907 21335
rect 10885 21301 10919 21335
rect 11345 21301 11379 21335
rect 14933 21301 14967 21335
rect 16681 21301 16715 21335
rect 16865 21301 16899 21335
rect 18153 21301 18187 21335
rect 18981 21301 19015 21335
rect 20039 21301 20073 21335
rect 2881 21097 2915 21131
rect 5917 21097 5951 21131
rect 7113 21097 7147 21131
rect 12265 21097 12299 21131
rect 14013 21097 14047 21131
rect 15025 21097 15059 21131
rect 2605 21029 2639 21063
rect 4537 21029 4571 21063
rect 5641 21029 5675 21063
rect 15393 21029 15427 21063
rect 15485 21029 15519 21063
rect 17049 21029 17083 21063
rect 18521 21029 18555 21063
rect 18613 21029 18647 21063
rect 21005 21029 21039 21063
rect 21097 21029 21131 21063
rect 1777 20961 1811 20995
rect 2053 20961 2087 20995
rect 3341 20961 3375 20995
rect 5273 20961 5307 20995
rect 6377 20961 6411 20995
rect 6561 20961 6595 20995
rect 7941 20961 7975 20995
rect 8217 20961 8251 20995
rect 8585 20961 8619 20995
rect 9689 20961 9723 20995
rect 9965 20961 9999 20995
rect 11253 20961 11287 20995
rect 11529 20961 11563 20995
rect 12909 20961 12943 20995
rect 13553 20961 13587 20995
rect 2237 20893 2271 20927
rect 4445 20893 4479 20927
rect 4905 20893 4939 20927
rect 6745 20893 6779 20927
rect 8309 20893 8343 20927
rect 10149 20893 10183 20927
rect 11345 20893 11379 20927
rect 11989 20893 12023 20927
rect 16957 20893 16991 20927
rect 17601 20893 17635 20927
rect 19165 20893 19199 20927
rect 3801 20825 3835 20859
rect 7481 20825 7515 20859
rect 9045 20825 9079 20859
rect 9781 20825 9815 20859
rect 15945 20825 15979 20859
rect 21557 20825 21591 20859
rect 4675 20757 4709 20791
rect 4813 20757 4847 20791
rect 8677 20757 8711 20791
rect 9413 20757 9447 20791
rect 10701 20757 10735 20791
rect 11161 20757 11195 20791
rect 12633 20757 12667 20791
rect 3065 20553 3099 20587
rect 4261 20553 4295 20587
rect 4629 20553 4663 20587
rect 5733 20553 5767 20587
rect 6101 20553 6135 20587
rect 9229 20553 9263 20587
rect 11437 20553 11471 20587
rect 19441 20553 19475 20587
rect 20821 20553 20855 20587
rect 21465 20553 21499 20587
rect 4491 20485 4525 20519
rect 8493 20485 8527 20519
rect 9597 20485 9631 20519
rect 10701 20485 10735 20519
rect 20177 20485 20211 20519
rect 2697 20417 2731 20451
rect 3157 20417 3191 20451
rect 3893 20417 3927 20451
rect 4721 20417 4755 20451
rect 13921 20417 13955 20451
rect 1409 20349 1443 20383
rect 2936 20349 2970 20383
rect 7205 20349 7239 20383
rect 7481 20349 7515 20383
rect 8712 20349 8746 20383
rect 9689 20349 9723 20383
rect 10241 20349 10275 20383
rect 11253 20349 11287 20383
rect 11897 20349 11931 20383
rect 12265 20349 12299 20383
rect 12449 20349 12483 20383
rect 12909 20349 12943 20383
rect 14289 20349 14323 20383
rect 14565 20349 14599 20383
rect 15025 20349 15059 20383
rect 15485 20349 15519 20383
rect 15853 20349 15887 20383
rect 16129 20349 16163 20383
rect 18337 20349 18371 20383
rect 18521 20349 18555 20383
rect 19692 20349 19726 20383
rect 20980 20349 21014 20383
rect 2789 20281 2823 20315
rect 4353 20281 4387 20315
rect 5089 20281 5123 20315
rect 6561 20281 6595 20315
rect 8033 20281 8067 20315
rect 8815 20281 8849 20315
rect 10425 20281 10459 20315
rect 16865 20281 16899 20315
rect 17877 20281 17911 20315
rect 21741 20281 21775 20315
rect 1593 20213 1627 20247
rect 2053 20213 2087 20247
rect 3433 20213 3467 20247
rect 5457 20213 5491 20247
rect 7021 20213 7055 20247
rect 11161 20213 11195 20247
rect 12541 20213 12575 20247
rect 13461 20213 13495 20247
rect 14105 20213 14139 20247
rect 15669 20213 15703 20247
rect 17233 20213 17267 20247
rect 18153 20213 18187 20247
rect 19073 20213 19107 20247
rect 19763 20213 19797 20247
rect 21051 20213 21085 20247
rect 1547 20009 1581 20043
rect 1869 20009 1903 20043
rect 5457 20009 5491 20043
rect 5917 20009 5951 20043
rect 6101 20009 6135 20043
rect 15393 20009 15427 20043
rect 16957 20009 16991 20043
rect 18521 20009 18555 20043
rect 21097 20009 21131 20043
rect 3893 19941 3927 19975
rect 7113 19941 7147 19975
rect 7665 19941 7699 19975
rect 10425 19941 10459 19975
rect 1476 19873 1510 19907
rect 2421 19873 2455 19907
rect 2697 19873 2731 19907
rect 4445 19873 4479 19907
rect 4675 19873 4709 19907
rect 6009 19873 6043 19907
rect 6469 19873 6503 19907
rect 8309 19873 8343 19907
rect 8493 19873 8527 19907
rect 8953 19873 8987 19907
rect 9689 19873 9723 19907
rect 10149 19873 10183 19907
rect 11253 19873 11287 19907
rect 11713 19873 11747 19907
rect 12817 19873 12851 19907
rect 12909 19873 12943 19907
rect 13093 19873 13127 19907
rect 15577 19873 15611 19907
rect 15761 19873 15795 19907
rect 16865 19873 16899 19907
rect 17417 19873 17451 19907
rect 18613 19873 18647 19907
rect 18889 19873 18923 19907
rect 19625 19873 19659 19907
rect 20913 19873 20947 19907
rect 3157 19805 3191 19839
rect 4261 19805 4295 19839
rect 4813 19805 4847 19839
rect 5181 19805 5215 19839
rect 11989 19805 12023 19839
rect 13277 19805 13311 19839
rect 14381 19805 14415 19839
rect 15117 19805 15151 19839
rect 2513 19737 2547 19771
rect 18061 19737 18095 19771
rect 2237 19669 2271 19703
rect 3433 19669 3467 19703
rect 4583 19669 4617 19703
rect 9045 19669 9079 19703
rect 9413 19669 9447 19703
rect 10793 19669 10827 19703
rect 11161 19669 11195 19703
rect 12541 19669 12575 19703
rect 14105 19669 14139 19703
rect 4997 19465 5031 19499
rect 9229 19465 9263 19499
rect 9321 19465 9355 19499
rect 10609 19465 10643 19499
rect 11253 19465 11287 19499
rect 13553 19465 13587 19499
rect 13645 19465 13679 19499
rect 14151 19465 14185 19499
rect 16865 19465 16899 19499
rect 21327 19465 21361 19499
rect 2513 19397 2547 19431
rect 2789 19397 2823 19431
rect 6009 19397 6043 19431
rect 5365 19329 5399 19363
rect 1409 19261 1443 19295
rect 1961 19261 1995 19295
rect 3008 19261 3042 19295
rect 3985 19261 4019 19295
rect 4445 19261 4479 19295
rect 5549 19261 5583 19295
rect 6285 19397 6319 19431
rect 7021 19397 7055 19431
rect 6101 19261 6135 19295
rect 3433 19193 3467 19227
rect 6009 19193 6043 19227
rect 14289 19397 14323 19431
rect 18705 19397 18739 19431
rect 13645 19329 13679 19363
rect 14381 19329 14415 19363
rect 20177 19329 20211 19363
rect 6837 19261 6871 19295
rect 7665 19261 7699 19295
rect 7941 19261 7975 19295
rect 8401 19261 8435 19295
rect 9229 19261 9263 19295
rect 9505 19261 9539 19295
rect 10057 19261 10091 19295
rect 11069 19261 11103 19295
rect 11529 19261 11563 19295
rect 12449 19261 12483 19295
rect 12909 19261 12943 19295
rect 13737 19261 13771 19295
rect 15577 19261 15611 19295
rect 16037 19261 16071 19295
rect 19625 19261 19659 19295
rect 20085 19261 20119 19295
rect 21224 19261 21258 19295
rect 21649 19261 21683 19295
rect 10241 19193 10275 19227
rect 1501 19125 1535 19159
rect 3111 19125 3145 19159
rect 3893 19125 3927 19159
rect 4261 19125 4295 19159
rect 5733 19125 5767 19159
rect 6285 19125 6319 19159
rect 6561 19125 6595 19159
rect 7389 19125 7423 19159
rect 7665 19125 7699 19159
rect 7757 19125 7791 19159
rect 8033 19125 8067 19159
rect 8769 19125 8803 19159
rect 10977 19125 11011 19159
rect 11529 19125 11563 19159
rect 11713 19125 11747 19159
rect 12541 19125 12575 19159
rect 14012 19193 14046 19227
rect 15393 19193 15427 19227
rect 18153 19193 18187 19227
rect 18245 19193 18279 19227
rect 13829 19125 13863 19159
rect 14841 19125 14875 19159
rect 15117 19125 15151 19159
rect 15669 19125 15703 19159
rect 17325 19125 17359 19159
rect 17785 19125 17819 19159
rect 19073 19125 19107 19159
rect 19533 19125 19567 19159
rect 20913 19125 20947 19159
rect 6745 18921 6779 18955
rect 8309 18921 8343 18955
rect 9919 18921 9953 18955
rect 10241 18853 10275 18887
rect 12081 18853 12115 18887
rect 12449 18853 12483 18887
rect 2053 18785 2087 18819
rect 2329 18785 2363 18819
rect 3341 18785 3375 18819
rect 4261 18785 4295 18819
rect 4491 18785 4525 18819
rect 5825 18785 5859 18819
rect 6193 18785 6227 18819
rect 7481 18785 7515 18819
rect 7665 18785 7699 18819
rect 9413 18785 9447 18819
rect 9597 18785 9631 18819
rect 9816 18785 9850 18819
rect 11069 18785 11103 18819
rect 11529 18785 11563 18819
rect 12909 18785 12943 18819
rect 13093 18785 13127 18819
rect 2513 18717 2547 18751
rect 4629 18717 4663 18751
rect 5457 18717 5491 18751
rect 6377 18717 6411 18751
rect 7941 18717 7975 18751
rect 8953 18717 8987 18751
rect 2881 18649 2915 18683
rect 3893 18649 3927 18683
rect 1685 18581 1719 18615
rect 5089 18581 5123 18615
rect 7021 18581 7055 18615
rect 8585 18581 8619 18615
rect 11805 18717 11839 18751
rect 13277 18717 13311 18751
rect 10609 18649 10643 18683
rect 14013 18921 14047 18955
rect 15117 18921 15151 18955
rect 16313 18921 16347 18955
rect 18889 18921 18923 18955
rect 16037 18853 16071 18887
rect 21097 18853 21131 18887
rect 14264 18785 14298 18819
rect 15393 18785 15427 18819
rect 16957 18785 16991 18819
rect 17325 18785 17359 18819
rect 18153 18785 18187 18819
rect 18337 18785 18371 18819
rect 19441 18785 19475 18819
rect 14657 18717 14691 18751
rect 17417 18717 17451 18751
rect 18567 18717 18601 18751
rect 21005 18717 21039 18751
rect 21373 18717 21407 18751
rect 13645 18581 13679 18615
rect 13921 18581 13955 18615
rect 14335 18581 14369 18615
rect 19579 18581 19613 18615
rect 2789 18377 2823 18411
rect 3414 18377 3448 18411
rect 3893 18377 3927 18411
rect 4353 18377 4387 18411
rect 5641 18377 5675 18411
rect 5917 18377 5951 18411
rect 6193 18377 6227 18411
rect 9597 18377 9631 18411
rect 9781 18377 9815 18411
rect 12265 18377 12299 18411
rect 14841 18377 14875 18411
rect 15393 18377 15427 18411
rect 16957 18377 16991 18411
rect 21327 18377 21361 18411
rect 3525 18309 3559 18343
rect 3157 18241 3191 18275
rect 3617 18241 3651 18275
rect 5365 18241 5399 18275
rect 11621 18241 11655 18275
rect 20913 18309 20947 18343
rect 19717 18241 19751 18275
rect 19993 18241 20027 18275
rect 1685 18173 1719 18207
rect 1961 18173 1995 18207
rect 4721 18173 4755 18207
rect 5089 18173 5123 18207
rect 5273 18173 5307 18207
rect 5641 18173 5675 18207
rect 6469 18173 6503 18207
rect 6837 18173 6871 18207
rect 7297 18173 7331 18207
rect 8401 18173 8435 18207
rect 8953 18173 8987 18207
rect 10333 18173 10367 18207
rect 10701 18173 10735 18207
rect 12633 18173 12667 18207
rect 12909 18173 12943 18207
rect 14289 18173 14323 18207
rect 14473 18173 14507 18207
rect 14841 18173 14875 18207
rect 15853 18173 15887 18207
rect 16129 18173 16163 18207
rect 16405 18173 16439 18207
rect 17877 18173 17911 18207
rect 18061 18173 18095 18207
rect 18521 18173 18555 18207
rect 21224 18173 21258 18207
rect 21649 18173 21683 18207
rect 3249 18105 3283 18139
rect 7573 18105 7607 18139
rect 9137 18105 9171 18139
rect 9505 18105 9539 18139
rect 13921 18105 13955 18139
rect 17325 18105 17359 18139
rect 19809 18105 19843 18139
rect 22017 18105 22051 18139
rect 1501 18037 1535 18071
rect 6469 18037 6503 18071
rect 6561 18037 6595 18071
rect 7849 18037 7883 18071
rect 8217 18037 8251 18071
rect 10333 18037 10367 18071
rect 11345 18037 11379 18071
rect 12541 18037 12575 18071
rect 13553 18037 13587 18071
rect 14105 18037 14139 18071
rect 15025 18037 15059 18071
rect 15669 18037 15703 18071
rect 16405 18037 16439 18071
rect 16681 18037 16715 18071
rect 18153 18037 18187 18071
rect 19073 18037 19107 18071
rect 19441 18037 19475 18071
rect 949 17833 983 17867
rect 1869 17833 1903 17867
rect 3893 17833 3927 17867
rect 6285 17833 6319 17867
rect 6653 17833 6687 17867
rect 8401 17833 8435 17867
rect 10149 17833 10183 17867
rect 11437 17833 11471 17867
rect 11713 17833 11747 17867
rect 15393 17833 15427 17867
rect 16313 17833 16347 17867
rect 18153 17833 18187 17867
rect 18521 17833 18555 17867
rect 19809 17833 19843 17867
rect 21005 17833 21039 17867
rect 4261 17765 4295 17799
rect 1476 17697 1510 17731
rect 2697 17697 2731 17731
rect 2973 17697 3007 17731
rect 4997 17697 5031 17731
rect 5457 17697 5491 17731
rect 3157 17629 3191 17663
rect 5641 17629 5675 17663
rect 2329 17561 2363 17595
rect 9045 17765 9079 17799
rect 13001 17765 13035 17799
rect 16865 17765 16899 17799
rect 6837 17697 6871 17731
rect 7021 17697 7055 17731
rect 8620 17697 8654 17731
rect 10057 17697 10091 17731
rect 10609 17697 10643 17731
rect 11621 17697 11655 17731
rect 12081 17697 12115 17731
rect 12633 17697 12667 17731
rect 13185 17697 13219 17731
rect 13645 17697 13679 17731
rect 14289 17697 14323 17731
rect 15485 17697 15519 17731
rect 15853 17697 15887 17731
rect 17509 17697 17543 17731
rect 18245 17697 18279 17731
rect 18429 17697 18463 17731
rect 18889 17697 18923 17731
rect 20913 17697 20947 17731
rect 21465 17697 21499 17731
rect 7941 17629 7975 17663
rect 13737 17629 13771 17663
rect 14105 17629 14139 17663
rect 6377 17561 6411 17595
rect 9873 17561 9907 17595
rect 14933 17561 14967 17595
rect 18245 17561 18279 17595
rect 1547 17493 1581 17527
rect 3525 17493 3559 17527
rect 4905 17493 4939 17527
rect 6009 17493 6043 17527
rect 6285 17493 6319 17527
rect 7665 17493 7699 17527
rect 8723 17493 8757 17527
rect 9413 17493 9447 17527
rect 11069 17493 11103 17527
rect 14105 17493 14139 17527
rect 14565 17493 14599 17527
rect 16773 17493 16807 17527
rect 19441 17493 19475 17527
rect 2513 17289 2547 17323
rect 2881 17289 2915 17323
rect 3341 17289 3375 17323
rect 1685 17085 1719 17119
rect 1961 17085 1995 17119
rect 4445 17289 4479 17323
rect 9413 17289 9447 17323
rect 9965 17289 9999 17323
rect 10057 17289 10091 17323
rect 13553 17289 13587 17323
rect 13737 17289 13771 17323
rect 13829 17289 13863 17323
rect 16773 17289 16807 17323
rect 16957 17289 16991 17323
rect 17785 17289 17819 17323
rect 19073 17289 19107 17323
rect 19441 17289 19475 17323
rect 21373 17289 21407 17323
rect 21741 17289 21775 17323
rect 3525 17153 3559 17187
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 3341 17017 3375 17051
rect 4353 17017 4387 17051
rect 6653 17221 6687 17255
rect 7481 17221 7515 17255
rect 5089 17153 5123 17187
rect 6929 17153 6963 17187
rect 8493 17153 8527 17187
rect 8769 17153 8803 17187
rect 5457 17085 5491 17119
rect 5733 17085 5767 17119
rect 4721 17017 4755 17051
rect 5917 17017 5951 17051
rect 7021 17017 7055 17051
rect 8585 17017 8619 17051
rect 10609 17221 10643 17255
rect 11805 17221 11839 17255
rect 13645 17153 13679 17187
rect 10977 17085 11011 17119
rect 11345 17085 11379 17119
rect 11529 17085 11563 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 13185 17017 13219 17051
rect 15485 17153 15519 17187
rect 13737 17085 13771 17119
rect 14013 17085 14047 17119
rect 14473 17085 14507 17119
rect 15577 17085 15611 17119
rect 16037 17085 16071 17119
rect 18061 17153 18095 17187
rect 17233 17085 17267 17119
rect 18153 17085 18187 17119
rect 19717 17085 19751 17119
rect 21189 17085 21223 17119
rect 22109 17085 22143 17119
rect 15117 17017 15151 17051
rect 16313 17017 16347 17051
rect 16773 17017 16807 17051
rect 19625 17017 19659 17051
rect 1501 16949 1535 16983
rect 4445 16949 4479 16983
rect 6193 16949 6227 16983
rect 7849 16949 7883 16983
rect 8309 16949 8343 16983
rect 9965 16949 9999 16983
rect 12173 16949 12207 16983
rect 13645 16949 13679 16983
rect 14105 16949 14139 16983
rect 20913 16949 20947 16983
rect 1593 16745 1627 16779
rect 2053 16745 2087 16779
rect 2421 16745 2455 16779
rect 2697 16745 2731 16779
rect 3709 16745 3743 16779
rect 9413 16745 9447 16779
rect 11345 16745 11379 16779
rect 12541 16745 12575 16779
rect 14105 16745 14139 16779
rect 15117 16745 15151 16779
rect 16957 16745 16991 16779
rect 18337 16745 18371 16779
rect 18889 16745 18923 16779
rect 857 15997 891 16031
rect 949 16677 983 16711
rect 5635 16677 5669 16711
rect 7481 16677 7515 16711
rect 8217 16677 8251 16711
rect 8769 16677 8803 16711
rect 9873 16677 9907 16711
rect 16681 16677 16715 16711
rect 19441 16677 19475 16711
rect 21097 16677 21131 16711
rect 857 15589 891 15623
rect 857 13549 891 13583
rect 765 13481 799 13515
rect 857 13413 891 13447
rect 673 9877 707 9911
rect 765 13209 799 13243
rect 305 6613 339 6647
rect 397 9741 431 9775
rect 581 8449 615 8483
rect 673 6681 707 6715
rect 765 5525 799 5559
rect 1409 16609 1443 16643
rect 3040 16609 3074 16643
rect 4328 16609 4362 16643
rect 5273 16609 5307 16643
rect 6469 16609 6503 16643
rect 11437 16609 11471 16643
rect 11713 16609 11747 16643
rect 12817 16609 12851 16643
rect 13277 16609 13311 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 16957 16609 16991 16643
rect 17325 16609 17359 16643
rect 18429 16609 18463 16643
rect 18705 16609 18739 16643
rect 7021 16541 7055 16575
rect 8125 16541 8159 16575
rect 9781 16541 9815 16575
rect 10425 16541 10459 16575
rect 13553 16541 13587 16575
rect 15853 16541 15887 16575
rect 21005 16541 21039 16575
rect 21281 16541 21315 16575
rect 3111 16473 3145 16507
rect 4399 16473 4433 16507
rect 14381 16473 14415 16507
rect 17877 16473 17911 16507
rect 18521 16473 18555 16507
rect 4721 16405 4755 16439
rect 5181 16405 5215 16439
rect 6193 16405 6227 16439
rect 6929 16405 6963 16439
rect 7849 16405 7883 16439
rect 9137 16405 9171 16439
rect 10701 16405 10735 16439
rect 11069 16405 11103 16439
rect 16405 16405 16439 16439
rect 2053 16201 2087 16235
rect 2513 16201 2547 16235
rect 3433 16201 3467 16235
rect 1593 16133 1627 16167
rect 2697 16065 2731 16099
rect 1409 15997 1443 16031
rect 2789 15929 2823 15963
rect 3341 15929 3375 15963
rect 1685 15657 1719 15691
rect 3249 15657 3283 15691
rect 2329 15589 2363 15623
rect 2421 15589 2455 15623
rect 2973 15589 3007 15623
rect 3525 16201 3559 16235
rect 4445 16201 4479 16235
rect 5181 16201 5215 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 11115 16201 11149 16235
rect 12173 16201 12207 16235
rect 15393 16201 15427 16235
rect 17233 16201 17267 16235
rect 19073 16201 19107 16235
rect 4307 16133 4341 16167
rect 4813 16133 4847 16167
rect 8493 16133 8527 16167
rect 10885 16133 10919 16167
rect 11805 16133 11839 16167
rect 15209 16133 15243 16167
rect 19441 16133 19475 16167
rect 4537 16065 4571 16099
rect 7941 16065 7975 16099
rect 9229 16065 9263 16099
rect 10425 16065 10459 16099
rect 11437 16065 11471 16099
rect 13921 16065 13955 16099
rect 10149 15997 10183 16031
rect 11044 15997 11078 16031
rect 12449 15997 12483 16031
rect 12909 15997 12943 16031
rect 14289 15997 14323 16031
rect 14565 15997 14599 16031
rect 4169 15929 4203 15963
rect 7665 15929 7699 15963
rect 8042 15929 8076 15963
rect 8861 15929 8895 15963
rect 9505 15929 9539 15963
rect 9597 15929 9631 15963
rect 16865 16065 16899 16099
rect 22017 16065 22051 16099
rect 15853 15997 15887 16031
rect 16037 15997 16071 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 19717 15997 19751 16031
rect 21240 15997 21274 16031
rect 21327 15997 21361 16031
rect 16313 15929 16347 15963
rect 18797 15929 18831 15963
rect 19625 15929 19659 15963
rect 3525 15861 3559 15895
rect 3617 15861 3651 15895
rect 3985 15861 4019 15895
rect 5549 15861 5583 15895
rect 5733 15861 5767 15895
rect 6837 15861 6871 15895
rect 7297 15861 7331 15895
rect 12725 15861 12759 15895
rect 13461 15861 13495 15895
rect 14105 15861 14139 15895
rect 15209 15861 15243 15895
rect 20913 15861 20947 15895
rect 21649 15861 21683 15895
rect 4629 15657 4663 15691
rect 5365 15657 5399 15691
rect 5457 15657 5491 15691
rect 8953 15657 8987 15691
rect 14933 15657 14967 15691
rect 15117 15657 15151 15691
rect 19441 15657 19475 15691
rect 3617 15521 3651 15555
rect 4388 15521 4422 15555
rect 5641 15589 5675 15623
rect 6469 15589 6503 15623
rect 8125 15589 8159 15623
rect 8677 15589 8711 15623
rect 9873 15589 9907 15623
rect 11437 15589 11471 15623
rect 11989 15589 12023 15623
rect 4813 15453 4847 15487
rect 5457 15453 5491 15487
rect 12725 15521 12759 15555
rect 12817 15521 12851 15555
rect 13277 15521 13311 15555
rect 7665 15453 7699 15487
rect 8033 15453 8067 15487
rect 9781 15453 9815 15487
rect 11345 15453 11379 15487
rect 6193 15385 6227 15419
rect 6929 15385 6963 15419
rect 10333 15385 10367 15419
rect 10793 15385 10827 15419
rect 2053 15317 2087 15351
rect 3433 15317 3467 15351
rect 6009 15317 6043 15351
rect 7297 15317 7331 15351
rect 9321 15317 9355 15351
rect 11069 15317 11103 15351
rect 12541 15317 12575 15351
rect 2145 15113 2179 15147
rect 4905 15113 4939 15147
rect 11253 15113 11287 15147
rect 12587 15113 12621 15147
rect 1593 15045 1627 15079
rect 1409 14909 1443 14943
rect 1961 14909 1995 14943
rect 1547 14569 1581 14603
rect 1444 14433 1478 14467
rect 1961 14297 1995 14331
rect 1593 14025 1627 14059
rect 1915 13957 1949 13991
rect 1828 13821 1862 13855
rect 8401 15045 8435 15079
rect 11989 15045 12023 15079
rect 2697 14977 2731 15011
rect 3709 14977 3743 15011
rect 5733 14977 5767 15011
rect 7941 14977 7975 15011
rect 8677 14977 8711 15011
rect 10517 14977 10551 15011
rect 12484 14909 12518 14943
rect 3157 14841 3191 14875
rect 3617 14841 3651 14875
rect 4071 14841 4105 14875
rect 6929 14841 6963 14875
rect 7021 14841 7055 14875
rect 7573 14841 7607 14875
rect 8769 14841 8803 14875
rect 9321 14841 9355 14875
rect 9781 14841 9815 14875
rect 10241 14841 10275 14875
rect 10333 14841 10367 14875
rect 11621 14841 11655 14875
rect 13461 15453 13495 15487
rect 20913 15589 20947 15623
rect 15301 15521 15335 15555
rect 15761 15521 15795 15555
rect 17141 15521 17175 15555
rect 17417 15521 17451 15555
rect 18429 15521 18463 15555
rect 18981 15521 19015 15555
rect 21005 15521 21039 15555
rect 15853 15453 15887 15487
rect 17601 15453 17635 15487
rect 19073 15453 19107 15487
rect 14381 15385 14415 15419
rect 14933 15385 14967 15419
rect 18061 15385 18095 15419
rect 19809 15385 19843 15419
rect 14105 15317 14139 15351
rect 16313 15317 16347 15351
rect 16681 15317 16715 15351
rect 20177 15317 20211 15351
rect 20545 15317 20579 15351
rect 14749 15113 14783 15147
rect 15025 15113 15059 15147
rect 16313 15113 16347 15147
rect 13737 14977 13771 15011
rect 14013 14977 14047 15011
rect 12909 14909 12943 14943
rect 14105 14841 14139 14875
rect 14657 14841 14691 14875
rect 15301 14909 15335 14943
rect 15761 14909 15795 14943
rect 16037 14909 16071 14943
rect 16221 14909 16255 14943
rect 16313 14909 16347 14943
rect 16405 15113 16439 15147
rect 16589 15113 16623 15147
rect 17325 15113 17359 15147
rect 17785 15113 17819 15147
rect 20913 15113 20947 15147
rect 21741 15113 21775 15147
rect 21327 14977 21361 15011
rect 22017 14977 22051 15011
rect 19073 14909 19107 14943
rect 19441 14909 19475 14943
rect 19625 14909 19659 14943
rect 20085 14909 20119 14943
rect 21240 14909 21274 14943
rect 16405 14841 16439 14875
rect 18153 14841 18187 14875
rect 18245 14841 18279 14875
rect 18797 14841 18831 14875
rect 2421 14773 2455 14807
rect 4629 14773 4663 14807
rect 5365 14773 5399 14807
rect 6285 14773 6319 14807
rect 12725 14773 12759 14807
rect 13277 14773 13311 14807
rect 14749 14773 14783 14807
rect 16865 14773 16899 14807
rect 19717 14773 19751 14807
rect 3801 14569 3835 14603
rect 3893 14569 3927 14603
rect 5181 14569 5215 14603
rect 8217 14569 8251 14603
rect 8677 14569 8711 14603
rect 10517 14569 10551 14603
rect 12817 14569 12851 14603
rect 13369 14569 13403 14603
rect 14013 14569 14047 14603
rect 14335 14569 14369 14603
rect 15853 14569 15887 14603
rect 20361 14569 20395 14603
rect 2605 14501 2639 14535
rect 3617 14433 3651 14467
rect 2513 14365 2547 14399
rect 3065 14297 3099 14331
rect 4077 14501 4111 14535
rect 5635 14501 5669 14535
rect 6377 14501 6411 14535
rect 7618 14501 7652 14535
rect 10149 14501 10183 14535
rect 11063 14501 11097 14535
rect 14749 14501 14783 14535
rect 16313 14501 16347 14535
rect 16957 14501 16991 14535
rect 18521 14501 18555 14535
rect 19625 14501 19659 14535
rect 4399 14433 4433 14467
rect 5273 14365 5307 14399
rect 3893 14297 3927 14331
rect 2237 14229 2271 14263
rect 4721 14229 4755 14263
rect 6193 14229 6227 14263
rect 2605 14025 2639 14059
rect 2237 13889 2271 13923
rect 2916 13821 2950 13855
rect 3341 13821 3375 13855
rect 4261 13957 4295 13991
rect 4445 13957 4479 13991
rect 4721 13957 4755 13991
rect 3617 13753 3651 13787
rect 4813 13821 4847 13855
rect 5273 13821 5307 13855
rect 5549 13821 5583 13855
rect 6193 13821 6227 13855
rect 7297 14433 7331 14467
rect 9724 14433 9758 14467
rect 9827 14433 9861 14467
rect 14264 14433 14298 14467
rect 15669 14433 15703 14467
rect 20913 14433 20947 14467
rect 21189 14433 21223 14467
rect 10701 14365 10735 14399
rect 12449 14365 12483 14399
rect 16865 14365 16899 14399
rect 17325 14365 17359 14399
rect 18429 14365 18463 14399
rect 18797 14365 18831 14399
rect 21373 14365 21407 14399
rect 9321 14297 9355 14331
rect 11621 14297 11655 14331
rect 15577 14297 15611 14331
rect 19993 14297 20027 14331
rect 21005 14297 21039 14331
rect 22293 14297 22327 14331
rect 6561 14229 6595 14263
rect 6837 14229 6871 14263
rect 8953 14229 8987 14263
rect 11989 14229 12023 14263
rect 12265 14229 12299 14263
rect 15025 14229 15059 14263
rect 16589 14229 16623 14263
rect 18153 14229 18187 14263
rect 22017 14229 22051 14263
rect 8401 14025 8435 14059
rect 9597 14025 9631 14059
rect 11161 14025 11195 14059
rect 12265 14025 12299 14059
rect 14105 14025 14139 14059
rect 14473 14025 14507 14059
rect 14841 14025 14875 14059
rect 15071 14025 15105 14059
rect 16957 14025 16991 14059
rect 17785 14025 17819 14059
rect 19165 14025 19199 14059
rect 20913 14025 20947 14059
rect 22201 14025 22235 14059
rect 2145 13685 2179 13719
rect 3019 13685 3053 13719
rect 3709 13685 3743 13719
rect 4445 13685 4479 13719
rect 5825 13685 5859 13719
rect 6377 13685 6411 13719
rect 6469 13957 6503 13991
rect 8677 13957 8711 13991
rect 6653 13889 6687 13923
rect 7481 13889 7515 13923
rect 9045 13889 9079 13923
rect 9367 13889 9401 13923
rect 9264 13821 9298 13855
rect 7802 13753 7836 13787
rect 21373 13957 21407 13991
rect 10241 13889 10275 13923
rect 13185 13889 13219 13923
rect 18429 13889 18463 13923
rect 9781 13821 9815 13855
rect 14968 13821 15002 13855
rect 15393 13821 15427 13855
rect 16037 13821 16071 13855
rect 19533 13821 19567 13855
rect 19809 13821 19843 13855
rect 20177 13821 20211 13855
rect 21189 13821 21223 13855
rect 21741 13821 21775 13855
rect 10562 13753 10596 13787
rect 11805 13753 11839 13787
rect 13506 13753 13540 13787
rect 15853 13753 15887 13787
rect 6469 13685 6503 13719
rect 7297 13685 7331 13719
rect 9597 13685 9631 13719
rect 10149 13685 10183 13719
rect 11437 13685 11471 13719
rect 12633 13685 12667 13719
rect 13001 13685 13035 13719
rect 18153 13753 18187 13787
rect 18245 13753 18279 13787
rect 17233 13685 17267 13719
rect 19717 13685 19751 13719
rect 1041 13481 1075 13515
rect 6101 13481 6135 13515
rect 7067 13481 7101 13515
rect 10885 13481 10919 13515
rect 12449 13481 12483 13515
rect 13921 13481 13955 13515
rect 19073 13481 19107 13515
rect 20729 13481 20763 13515
rect 21005 13481 21039 13515
rect 2329 13413 2363 13447
rect 3525 13413 3559 13447
rect 5502 13413 5536 13447
rect 6745 13413 6779 13447
rect 8125 13413 8159 13447
rect 10051 13413 10085 13447
rect 11621 13413 11655 13447
rect 13322 13413 13356 13447
rect 15761 13413 15795 13447
rect 16037 13413 16071 13447
rect 16129 13413 16163 13447
rect 16405 13413 16439 13447
rect 16681 13413 16715 13447
rect 18245 13413 18279 13447
rect 20269 13413 20303 13447
rect 4236 13345 4270 13379
rect 5181 13345 5215 13379
rect 6377 13345 6411 13379
rect 6996 13345 7030 13379
rect 7481 13345 7515 13379
rect 15368 13345 15402 13379
rect 2237 13277 2271 13311
rect 2881 13277 2915 13311
rect 8033 13277 8067 13311
rect 9689 13277 9723 13311
rect 11529 13277 11563 13311
rect 13001 13277 13035 13311
rect 1961 13209 1995 13243
rect 8585 13209 8619 13243
rect 12081 13209 12115 13243
rect 19717 13345 19751 13379
rect 20913 13345 20947 13379
rect 21465 13345 21499 13379
rect 16589 13277 16623 13311
rect 17233 13277 17267 13311
rect 18153 13277 18187 13311
rect 18613 13277 18647 13311
rect 17601 13209 17635 13243
rect 19901 13209 19935 13243
rect 1041 13141 1075 13175
rect 1685 13141 1719 13175
rect 3157 13141 3191 13175
rect 4307 13141 4341 13175
rect 4813 13141 4847 13175
rect 8953 13141 8987 13175
rect 9321 13141 9355 13175
rect 10609 13141 10643 13175
rect 11253 13141 11287 13175
rect 12817 13141 12851 13175
rect 14565 13141 14599 13175
rect 15117 13141 15151 13175
rect 15439 13141 15473 13175
rect 16037 13141 16071 13175
rect 17877 13141 17911 13175
rect 19441 13141 19475 13175
rect 21925 13141 21959 13175
rect 22293 13141 22327 13175
rect 4123 12937 4157 12971
rect 5917 12937 5951 12971
rect 8493 12937 8527 12971
rect 10609 12937 10643 12971
rect 12265 12937 12299 12971
rect 13829 12937 13863 12971
rect 16681 12937 16715 12971
rect 19441 12937 19475 12971
rect 20913 12937 20947 12971
rect 21373 12937 21407 12971
rect 22109 12937 22143 12971
rect 3433 12869 3467 12903
rect 7113 12869 7147 12903
rect 8125 12869 8159 12903
rect 11437 12869 11471 12903
rect 14841 12869 14875 12903
rect 17417 12869 17451 12903
rect 1685 12801 1719 12835
rect 2513 12801 2547 12835
rect 4997 12801 5031 12835
rect 7205 12801 7239 12835
rect 9045 12801 9079 12835
rect 9689 12801 9723 12835
rect 15669 12801 15703 12835
rect 18797 12801 18831 12835
rect 1444 12733 1478 12767
rect 1869 12733 1903 12767
rect 3801 12733 3835 12767
rect 4052 12733 4086 12767
rect 4537 12733 4571 12767
rect 12484 12733 12518 12767
rect 12909 12733 12943 12767
rect 13921 12733 13955 12767
rect 15393 12733 15427 12767
rect 19901 12733 19935 12767
rect 20177 12733 20211 12767
rect 21189 12733 21223 12767
rect 21741 12733 21775 12767
rect 2605 12665 2639 12699
rect 3157 12665 3191 12699
rect 4905 12665 4939 12699
rect 5318 12665 5352 12699
rect 7526 12665 7560 12699
rect 9137 12665 9171 12699
rect 10885 12665 10919 12699
rect 10977 12665 11011 12699
rect 14243 12665 14277 12699
rect 16031 12665 16065 12699
rect 18153 12665 18187 12699
rect 18245 12665 18279 12699
rect 19165 12665 19199 12699
rect 2237 12597 2271 12631
rect 6193 12597 6227 12631
rect 6561 12597 6595 12631
rect 8769 12597 8803 12631
rect 10057 12597 10091 12631
rect 10517 12597 10551 12631
rect 11897 12597 11931 12631
rect 12587 12597 12621 12631
rect 13369 12597 13403 12631
rect 16865 12597 16899 12631
rect 17785 12597 17819 12631
rect 19717 12597 19751 12631
rect 949 12393 983 12427
rect 1639 12393 1673 12427
rect 2053 12393 2087 12427
rect 2651 12393 2685 12427
rect 7205 12393 7239 12427
rect 7665 12393 7699 12427
rect 11345 12393 11379 12427
rect 11713 12393 11747 12427
rect 12541 12393 12575 12427
rect 13461 12393 13495 12427
rect 14013 12393 14047 12427
rect 15393 12393 15427 12427
rect 16681 12393 16715 12427
rect 17187 12393 17221 12427
rect 19763 12393 19797 12427
rect 20177 12393 20211 12427
rect 21005 12393 21039 12427
rect 4261 12325 4295 12359
rect 6285 12325 6319 12359
rect 6377 12325 6411 12359
rect 8217 12325 8251 12359
rect 8769 12325 8803 12359
rect 14657 12325 14691 12359
rect 16405 12325 16439 12359
rect 18245 12325 18279 12359
rect 1536 12257 1570 12291
rect 2580 12257 2614 12291
rect 4813 12257 4847 12291
rect 7113 12257 7147 12291
rect 12449 12257 12483 12291
rect 12909 12257 12943 12291
rect 14264 12257 14298 12291
rect 14473 12257 14507 12291
rect 15485 12257 15519 12291
rect 15853 12257 15887 12291
rect 17116 12257 17150 12291
rect 19660 12257 19694 12291
rect 20913 12257 20947 12291
rect 21373 12257 21407 12291
rect 4169 12189 4203 12223
rect 8125 12189 8159 12223
rect 10149 12189 10183 12223
rect 5917 12121 5951 12155
rect 9413 12121 9447 12155
rect 14335 12121 14369 12155
rect 15025 12189 15059 12223
rect 18153 12189 18187 12223
rect 19073 12189 19107 12223
rect 18705 12121 18739 12155
rect 19441 12121 19475 12155
rect 2329 12053 2363 12087
rect 3065 12053 3099 12087
rect 3433 12053 3467 12087
rect 3709 12053 3743 12087
rect 5181 12053 5215 12087
rect 5549 12053 5583 12087
rect 9045 12053 9079 12087
rect 9965 12053 9999 12087
rect 11069 12053 11103 12087
rect 12081 12053 12115 12087
rect 14473 12053 14507 12087
rect 17601 12053 17635 12087
rect 17877 12053 17911 12087
rect 20453 12053 20487 12087
rect 21925 12053 21959 12087
rect 22293 12053 22327 12087
rect 6193 11849 6227 11883
rect 7757 11849 7791 11883
rect 8125 11849 8159 11883
rect 9505 11849 9539 11883
rect 14013 11849 14047 11883
rect 15071 11849 15105 11883
rect 17785 11849 17819 11883
rect 19073 11849 19107 11883
rect 19441 11849 19475 11883
rect 20913 11849 20947 11883
rect 21373 11849 21407 11883
rect 22109 11849 22143 11883
rect 5457 11781 5491 11815
rect 16865 11781 16899 11815
rect 21833 11781 21867 11815
rect 1961 11713 1995 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 8585 11713 8619 11747
rect 9873 11713 9907 11747
rect 12265 11713 12299 11747
rect 13093 11713 13127 11747
rect 15393 11713 15427 11747
rect 15945 11713 15979 11747
rect 18797 11713 18831 11747
rect 19717 11713 19751 11747
rect 3744 11645 3778 11679
rect 4169 11645 4203 11679
rect 5273 11645 5307 11679
rect 5825 11645 5859 11679
rect 10149 11645 10183 11679
rect 10885 11645 10919 11679
rect 11161 11645 11195 11679
rect 15000 11645 15034 11679
rect 17233 11645 17267 11679
rect 21189 11645 21223 11679
rect 2282 11577 2316 11611
rect 4537 11577 4571 11611
rect 4905 11577 4939 11611
rect 7158 11577 7192 11611
rect 8217 11577 8251 11611
rect 8401 11577 8435 11611
rect 8906 11577 8940 11611
rect 13455 11577 13489 11611
rect 15761 11577 15795 11611
rect 16266 11577 16300 11611
rect 18153 11577 18187 11611
rect 18245 11577 18279 11611
rect 19809 11577 19843 11611
rect 20361 11577 20395 11611
rect 1777 11509 1811 11543
rect 2881 11509 2915 11543
rect 3157 11509 3191 11543
rect 3525 11509 3559 11543
rect 3847 11509 3881 11543
rect 10701 11509 10735 11543
rect 11897 11509 11931 11543
rect 13001 11509 13035 11543
rect 14381 11509 14415 11543
rect 14841 11509 14875 11543
rect 5641 11305 5675 11339
rect 7113 11305 7147 11339
rect 7665 11305 7699 11339
rect 2558 11237 2592 11271
rect 4261 11237 4295 11271
rect 6009 11237 6043 11271
rect 3157 11169 3191 11203
rect 2237 11101 2271 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 5917 11101 5951 11135
rect 3525 11033 3559 11067
rect 4537 11033 4571 11067
rect 5273 11033 5307 11067
rect 6469 11033 6503 11067
rect 8769 11305 8803 11339
rect 9413 11305 9447 11339
rect 9873 11305 9907 11339
rect 10701 11305 10735 11339
rect 11989 11305 12023 11339
rect 14243 11305 14277 11339
rect 14933 11305 14967 11339
rect 16129 11305 16163 11339
rect 16681 11305 16715 11339
rect 17647 11305 17681 11339
rect 19717 11305 19751 11339
rect 20361 11305 20395 11339
rect 21005 11305 21039 11339
rect 11161 11237 11195 11271
rect 12633 11237 12667 11271
rect 12725 11237 12759 11271
rect 14565 11237 14599 11271
rect 18705 11237 18739 11271
rect 9689 11169 9723 11203
rect 11713 11169 11747 11203
rect 14105 11169 14139 11203
rect 15761 11169 15795 11203
rect 17509 11169 17543 11203
rect 20913 11169 20947 11203
rect 21373 11169 21407 11203
rect 7849 11101 7883 11135
rect 11069 11101 11103 11135
rect 13553 11101 13587 11135
rect 15485 11101 15519 11135
rect 18613 11101 18647 11135
rect 18889 11101 18923 11135
rect 13185 11033 13219 11067
rect 1685 10965 1719 10999
rect 1961 10965 1995 10999
rect 3893 10965 3927 10999
rect 4399 10965 4433 10999
rect 6837 10965 6871 10999
rect 7113 10965 7147 10999
rect 7297 10965 7331 10999
rect 9045 10965 9079 10999
rect 10241 10965 10275 10999
rect 12357 10965 12391 10999
rect 13921 10965 13955 10999
rect 16957 10965 16991 10999
rect 17325 10965 17359 10999
rect 18153 10965 18187 10999
rect 19993 10965 20027 10999
rect 21925 10965 21959 10999
rect 22293 10965 22327 10999
rect 1593 10761 1627 10795
rect 2421 10761 2455 10795
rect 4353 10761 4387 10795
rect 5733 10761 5767 10795
rect 9229 10761 9263 10795
rect 11345 10761 11379 10795
rect 14105 10761 14139 10795
rect 15853 10761 15887 10795
rect 17601 10761 17635 10795
rect 19073 10761 19107 10795
rect 19763 10761 19797 10795
rect 20545 10761 20579 10795
rect 20913 10761 20947 10795
rect 21741 10761 21775 10795
rect 6377 10693 6411 10727
rect 10977 10693 11011 10727
rect 21373 10693 21407 10727
rect 7573 10625 7607 10659
rect 8309 10625 8343 10659
rect 13553 10625 13587 10659
rect 14565 10625 14599 10659
rect 14841 10625 14875 10659
rect 16037 10625 16071 10659
rect 18153 10625 18187 10659
rect 19441 10625 19475 10659
rect 949 10557 983 10591
rect 1409 10557 1443 10591
rect 2513 10557 2547 10591
rect 2697 10557 2731 10591
rect 4813 10557 4847 10591
rect 8401 10557 8435 10591
rect 9413 10557 9447 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 16957 10557 16991 10591
rect 19660 10557 19694 10591
rect 20085 10557 20119 10591
rect 21189 10557 21223 10591
rect 6929 10489 6963 10523
rect 7021 10489 7055 10523
rect 1777 10421 1811 10455
rect 1961 10421 1995 10455
rect 2789 10421 2823 10455
rect 3433 10421 3467 10455
rect 3709 10421 3743 10455
rect 4721 10421 4755 10455
rect 5181 10421 5215 10455
rect 6009 10421 6043 10455
rect 1777 10217 1811 10251
rect 2605 10217 2639 10251
rect 2973 10217 3007 10251
rect 3341 10217 3375 10251
rect 3709 10217 3743 10251
rect 4169 10217 4203 10251
rect 4353 10217 4387 10251
rect 5457 10217 5491 10251
rect 7205 10217 7239 10251
rect 7751 10217 7785 10251
rect 1409 10081 1443 10115
rect 2329 9945 2363 9979
rect 2329 9673 2363 9707
rect 3571 9673 3605 9707
rect 1409 9537 1443 9571
rect 2605 9537 2639 9571
rect 6003 10149 6037 10183
rect 4664 10081 4698 10115
rect 4767 10081 4801 10115
rect 7389 10081 7423 10115
rect 5641 10013 5675 10047
rect 5181 9945 5215 9979
rect 6561 9945 6595 9979
rect 6837 9877 6871 9911
rect 8309 9877 8343 9911
rect 7665 9673 7699 9707
rect 4721 9605 4755 9639
rect 6101 9605 6135 9639
rect 7481 9605 7515 9639
rect 4813 9537 4847 9571
rect 3468 9469 3502 9503
rect 3893 9469 3927 9503
rect 4169 9469 4203 9503
rect 4592 9469 4626 9503
rect 5457 9469 5491 9503
rect 1771 9401 1805 9435
rect 4445 9401 4479 9435
rect 5181 9401 5215 9435
rect 6193 9537 6227 9571
rect 6929 9401 6963 9435
rect 7021 9401 7055 9435
rect 7849 9401 7883 9435
rect 2973 9333 3007 9367
rect 4169 9333 4203 9367
rect 5917 9333 5951 9367
rect 6101 9333 6135 9367
rect 6561 9333 6595 9367
rect 7665 9333 7699 9367
rect 12265 10489 12299 10523
rect 12541 10489 12575 10523
rect 12642 10489 12676 10523
rect 13185 10489 13219 10523
rect 14657 10489 14691 10523
rect 16358 10489 16392 10523
rect 18245 10489 18279 10523
rect 18797 10489 18831 10523
rect 8585 10421 8619 10455
rect 10425 10421 10459 10455
rect 11805 10421 11839 10455
rect 22109 10421 22143 10455
rect 9827 10217 9861 10251
rect 11253 10217 11287 10251
rect 12265 10217 12299 10251
rect 12633 10217 12667 10251
rect 13921 10217 13955 10251
rect 14565 10217 14599 10251
rect 15669 10217 15703 10251
rect 16037 10217 16071 10251
rect 16589 10217 16623 10251
rect 19717 10217 19751 10251
rect 20453 10217 20487 10251
rect 21005 10217 21039 10251
rect 8953 10149 8987 10183
rect 10333 10149 10367 10183
rect 13046 10149 13080 10183
rect 17417 10149 17451 10183
rect 18889 10149 18923 10183
rect 8677 10081 8711 10115
rect 9597 10081 9631 10115
rect 10517 10081 10551 10115
rect 10701 10081 10735 10115
rect 11529 10081 11563 10115
rect 11764 10081 11798 10115
rect 11989 10081 12023 10115
rect 12725 10081 12759 10115
rect 16164 10081 16198 10115
rect 16267 10081 16301 10115
rect 17760 10081 17794 10115
rect 20913 10081 20947 10115
rect 21465 10081 21499 10115
rect 11851 10013 11885 10047
rect 10333 9945 10367 9979
rect 9413 9877 9447 9911
rect 10149 9877 10183 9911
rect 10839 9877 10873 9911
rect 9689 9673 9723 9707
rect 10379 9673 10413 9707
rect 11391 9605 11425 9639
rect 11069 9537 11103 9571
rect 9413 9469 9447 9503
rect 10308 9469 10342 9503
rect 11320 9469 11354 9503
rect 11529 9469 11563 9503
rect 8769 9401 8803 9435
rect 8861 9401 8895 9435
rect 10793 9401 10827 9435
rect 14841 10013 14875 10047
rect 18797 10013 18831 10047
rect 20085 10013 20119 10047
rect 13645 9945 13679 9979
rect 19349 9945 19383 9979
rect 22293 9945 22327 9979
rect 16957 9877 16991 9911
rect 17969 9877 18003 9911
rect 18245 9877 18279 9911
rect 18521 9877 18555 9911
rect 21925 9877 21959 9911
rect 13093 9673 13127 9707
rect 15301 9673 15335 9707
rect 17141 9673 17175 9707
rect 17785 9673 17819 9707
rect 19763 9673 19797 9707
rect 20913 9673 20947 9707
rect 21373 9673 21407 9707
rect 15393 9605 15427 9639
rect 20637 9605 20671 9639
rect 13507 9537 13541 9571
rect 16221 9537 16255 9571
rect 18429 9537 18463 9571
rect 22109 9537 22143 9571
rect 13404 9469 13438 9503
rect 13829 9469 13863 9503
rect 14381 9469 14415 9503
rect 15393 9469 15427 9503
rect 15945 9469 15979 9503
rect 16865 9469 16899 9503
rect 19692 9469 19726 9503
rect 21189 9469 21223 9503
rect 16313 9401 16347 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 21833 9401 21867 9435
rect 8401 9333 8435 9367
rect 8585 9333 8619 9367
rect 10057 9333 10091 9367
rect 11529 9333 11563 9367
rect 11713 9333 11747 9367
rect 11989 9333 12023 9367
rect 12173 9333 12207 9367
rect 12725 9333 12759 9367
rect 14197 9333 14231 9367
rect 14749 9333 14783 9367
rect 15577 9333 15611 9367
rect 19073 9333 19107 9367
rect 19441 9333 19475 9367
rect 20177 9333 20211 9367
rect 1547 9129 1581 9163
rect 5641 9129 5675 9163
rect 1823 9061 1857 9095
rect 2145 9061 2179 9095
rect 3709 9061 3743 9095
rect 1444 8993 1478 9027
rect 1720 8993 1754 9027
rect 2697 8993 2731 9027
rect 2053 8925 2087 8959
rect 3341 8925 3375 8959
rect 857 4981 891 5015
rect 949 8857 983 8891
rect 489 4437 523 4471
rect 4997 9061 5031 9095
rect 4721 8993 4755 9027
rect 7941 9129 7975 9163
rect 8217 9129 8251 9163
rect 6653 9061 6687 9095
rect 7205 9061 7239 9095
rect 8033 8993 8067 9027
rect 6561 8925 6595 8959
rect 6285 8857 6319 8891
rect 7481 8857 7515 8891
rect 3065 8789 3099 8823
rect 4169 8789 4203 8823
rect 5917 8789 5951 8823
rect 6101 8789 6135 8823
rect 10241 9129 10275 9163
rect 10425 9129 10459 9163
rect 8585 8993 8619 9027
rect 9689 8993 9723 9027
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 11253 9129 11287 9163
rect 14473 9129 14507 9163
rect 15439 9129 15473 9163
rect 16221 9129 16255 9163
rect 19855 9129 19889 9163
rect 12909 9061 12943 9095
rect 16726 9061 16760 9095
rect 18061 9061 18095 9095
rect 18337 9061 18371 9095
rect 20545 9061 20579 9095
rect 21005 9061 21039 9095
rect 21097 9061 21131 9095
rect 10885 8993 10919 9027
rect 15368 8993 15402 9027
rect 16405 8993 16439 9027
rect 18889 8993 18923 9027
rect 19717 8993 19751 9027
rect 12173 8925 12207 8959
rect 12817 8925 12851 8959
rect 18245 8925 18279 8959
rect 20177 8925 20211 8959
rect 22293 8925 22327 8959
rect 12449 8857 12483 8891
rect 13369 8857 13403 8891
rect 17601 8857 17635 8891
rect 21557 8857 21591 8891
rect 8769 8789 8803 8823
rect 9873 8789 9907 8823
rect 10425 8789 10459 8823
rect 10609 8789 10643 8823
rect 11805 8789 11839 8823
rect 13737 8789 13771 8823
rect 14841 8789 14875 8823
rect 15761 8789 15795 8823
rect 17325 8789 17359 8823
rect 19165 8789 19199 8823
rect 19625 8789 19659 8823
rect 21925 8789 21959 8823
rect 1547 8585 1581 8619
rect 3433 8585 3467 8619
rect 3985 8585 4019 8619
rect 6101 8585 6135 8619
rect 6193 8585 6227 8619
rect 6561 8585 6595 8619
rect 8125 8585 8159 8619
rect 11713 8585 11747 8619
rect 13461 8585 13495 8619
rect 13829 8585 13863 8619
rect 15117 8585 15151 8619
rect 16405 8585 16439 8619
rect 16865 8585 16899 8619
rect 17095 8585 17129 8619
rect 19533 8585 19567 8619
rect 20913 8585 20947 8619
rect 21327 8585 21361 8619
rect 1409 8381 1443 8415
rect 1720 8381 1754 8415
rect 2237 8313 2271 8347
rect 2329 8313 2363 8347
rect 2881 8313 2915 8347
rect 3249 8313 3283 8347
rect 4997 8517 5031 8551
rect 5089 8517 5123 8551
rect 11069 8517 11103 8551
rect 16129 8517 16163 8551
rect 22017 8517 22051 8551
rect 3709 8381 3743 8415
rect 3893 8381 3927 8415
rect 1823 8245 1857 8279
rect 3433 8245 3467 8279
rect 3617 8245 3651 8279
rect 4629 8245 4663 8279
rect 5917 8449 5951 8483
rect 8677 8449 8711 8483
rect 9321 8449 9355 8483
rect 9781 8449 9815 8483
rect 10149 8449 10183 8483
rect 12541 8449 12575 8483
rect 14749 8449 14783 8483
rect 18153 8449 18187 8483
rect 19717 8449 19751 8483
rect 6837 8381 6871 8415
rect 7481 8381 7515 8415
rect 7941 8381 7975 8415
rect 5273 8313 5307 8347
rect 5365 8313 5399 8347
rect 9137 8381 9171 8415
rect 15209 8381 15243 8415
rect 17024 8381 17058 8415
rect 17417 8381 17451 8415
rect 18797 8381 18831 8415
rect 21256 8381 21290 8415
rect 21741 8381 21775 8415
rect 8401 8313 8435 8347
rect 8493 8313 8527 8347
rect 7021 8245 7055 8279
rect 7941 8245 7975 8279
rect 10511 8313 10545 8347
rect 12633 8313 12667 8347
rect 13185 8313 13219 8347
rect 15530 8313 15564 8347
rect 18245 8313 18279 8347
rect 19809 8313 19843 8347
rect 20361 8313 20395 8347
rect 11437 8245 11471 8279
rect 12173 8245 12207 8279
rect 14013 8245 14047 8279
rect 17785 8245 17819 8279
rect 19073 8245 19107 8279
rect 22477 8245 22511 8279
rect 8171 8041 8205 8075
rect 8953 8041 8987 8075
rect 10241 8041 10275 8075
rect 12449 8041 12483 8075
rect 13001 8041 13035 8075
rect 16957 8041 16991 8075
rect 2237 7973 2271 8007
rect 3065 7973 3099 8007
rect 5083 7973 5117 8007
rect 5917 7973 5951 8007
rect 6285 7973 6319 8007
rect 6561 7973 6595 8007
rect 6653 7973 6687 8007
rect 8493 7973 8527 8007
rect 1476 7905 1510 7939
rect 1736 7905 1770 7939
rect 4721 7905 4755 7939
rect 8068 7905 8102 7939
rect 1823 7837 1857 7871
rect 2145 7837 2179 7871
rect 2973 7837 3007 7871
rect 3617 7837 3651 7871
rect 2697 7769 2731 7803
rect 7113 7769 7147 7803
rect 11069 7973 11103 8007
rect 11621 7973 11655 8007
rect 13093 7973 13127 8007
rect 13553 7973 13587 8007
rect 13645 7973 13679 8007
rect 16399 7973 16433 8007
rect 17509 7973 17543 8007
rect 18106 7973 18140 8007
rect 19671 7973 19705 8007
rect 21005 7973 21039 8007
rect 21097 7973 21131 8007
rect 9689 7837 9723 7871
rect 10977 7837 11011 7871
rect 12265 7769 12299 7803
rect 16037 7905 16071 7939
rect 18705 7905 18739 7939
rect 19584 7905 19618 7939
rect 14197 7837 14231 7871
rect 17233 7837 17267 7871
rect 17509 7837 17543 7871
rect 17785 7837 17819 7871
rect 19993 7837 20027 7871
rect 21281 7837 21315 7871
rect 13277 7769 13311 7803
rect 17601 7769 17635 7803
rect 1639 7701 1673 7735
rect 4261 7701 4295 7735
rect 5641 7701 5675 7735
rect 6193 7701 6227 7735
rect 7481 7701 7515 7735
rect 7849 7701 7883 7735
rect 9137 7701 9171 7735
rect 10517 7701 10551 7735
rect 11897 7701 11931 7735
rect 13093 7701 13127 7735
rect 14565 7701 14599 7735
rect 14841 7701 14875 7735
rect 15485 7701 15519 7735
rect 15945 7701 15979 7735
rect 18981 7701 19015 7735
rect 19349 7701 19383 7735
rect 20729 7701 20763 7735
rect 21925 7701 21959 7735
rect 22293 7701 22327 7735
rect 2421 7497 2455 7531
rect 2605 7497 2639 7531
rect 5549 7497 5583 7531
rect 2053 7429 2087 7463
rect 1501 7361 1535 7395
rect 2237 7293 2271 7327
rect 1593 7225 1627 7259
rect 3157 7361 3191 7395
rect 3985 7361 4019 7395
rect 5457 7293 5491 7327
rect 2881 7225 2915 7259
rect 2973 7225 3007 7259
rect 3709 7225 3743 7259
rect 3801 7225 3835 7259
rect 4813 7225 4847 7259
rect 4905 7225 4939 7259
rect 5641 7225 5675 7259
rect 6469 7497 6503 7531
rect 7757 7497 7791 7531
rect 8125 7497 8159 7531
rect 8309 7497 8343 7531
rect 6837 7361 6871 7395
rect 9597 7497 9631 7531
rect 9781 7497 9815 7531
rect 10149 7497 10183 7531
rect 10241 7497 10275 7531
rect 11805 7497 11839 7531
rect 13645 7497 13679 7531
rect 13921 7497 13955 7531
rect 15761 7497 15795 7531
rect 16129 7497 16163 7531
rect 20913 7497 20947 7531
rect 8769 7361 8803 7395
rect 8309 7293 8343 7327
rect 9413 7293 9447 7327
rect 9597 7293 9631 7327
rect 7199 7225 7233 7259
rect 8401 7225 8435 7259
rect 8838 7225 8872 7259
rect 2605 7157 2639 7191
rect 5733 7157 5767 7191
rect 6101 7157 6135 7191
rect 6285 7157 6319 7191
rect 11529 7429 11563 7463
rect 10609 7361 10643 7395
rect 17049 7429 17083 7463
rect 18797 7429 18831 7463
rect 20361 7429 20395 7463
rect 21465 7429 21499 7463
rect 14565 7361 14599 7395
rect 15209 7361 15243 7395
rect 16497 7361 16531 7395
rect 18245 7361 18279 7395
rect 12449 7293 12483 7327
rect 13921 7293 13955 7327
rect 19533 7293 19567 7327
rect 21281 7293 21315 7327
rect 21833 7293 21867 7327
rect 10425 7225 10459 7259
rect 10971 7225 11005 7259
rect 12811 7225 12845 7259
rect 14657 7225 14691 7259
rect 16589 7225 16623 7259
rect 18337 7225 18371 7259
rect 19809 7225 19843 7259
rect 19901 7225 19935 7259
rect 10241 7157 10275 7191
rect 12265 7157 12299 7191
rect 13369 7157 13403 7191
rect 14105 7157 14139 7191
rect 17417 7157 17451 7191
rect 17785 7157 17819 7191
rect 19165 7157 19199 7191
rect 22201 7157 22235 7191
rect 2421 6953 2455 6987
rect 4077 6953 4111 6987
rect 7297 6953 7331 6987
rect 8217 6953 8251 6987
rect 11069 6953 11103 6987
rect 12173 6953 12207 6987
rect 14657 6953 14691 6987
rect 15025 6953 15059 6987
rect 16313 6953 16347 6987
rect 17877 6953 17911 6987
rect 19165 6953 19199 6987
rect 19809 6953 19843 6987
rect 1863 6885 1897 6919
rect 2697 6885 2731 6919
rect 3249 6885 3283 6919
rect 1501 6817 1535 6851
rect 3392 6817 3426 6851
rect 3668 6817 3702 6851
rect 2605 6749 2639 6783
rect 3479 6749 3513 6783
rect 4490 6885 4524 6919
rect 6009 6885 6043 6919
rect 6101 6885 6135 6919
rect 6653 6885 6687 6919
rect 6745 6885 6779 6919
rect 9873 6885 9907 6919
rect 13737 6885 13771 6919
rect 13829 6885 13863 6919
rect 15761 6885 15795 6919
rect 16818 6885 16852 6919
rect 18566 6885 18600 6919
rect 21097 6885 21131 6919
rect 4169 6749 4203 6783
rect 5733 6749 5767 6783
rect 7849 6817 7883 6851
rect 9045 6817 9079 6851
rect 9321 6817 9355 6851
rect 9413 6817 9447 6851
rect 10793 6817 10827 6851
rect 11805 6817 11839 6851
rect 13369 6817 13403 6851
rect 15368 6817 15402 6851
rect 20453 6817 20487 6851
rect 5089 6681 5123 6715
rect 6745 6681 6779 6715
rect 8769 6681 8803 6715
rect 9781 6749 9815 6783
rect 10241 6749 10275 6783
rect 14013 6749 14047 6783
rect 16497 6749 16531 6783
rect 18245 6749 18279 6783
rect 21005 6749 21039 6783
rect 21925 6749 21959 6783
rect 12725 6681 12759 6715
rect 13001 6681 13035 6715
rect 17417 6681 17451 6715
rect 21557 6681 21591 6715
rect 3755 6613 3789 6647
rect 4077 6613 4111 6647
rect 5365 6613 5399 6647
rect 6929 6613 6963 6647
rect 7757 6613 7791 6647
rect 9321 6613 9355 6647
rect 11437 6613 11471 6647
rect 15439 6613 15473 6647
rect 20085 6613 20119 6647
rect 22293 6613 22327 6647
rect 1823 6409 1857 6443
rect 3065 6409 3099 6443
rect 4951 6409 4985 6443
rect 6975 6409 7009 6443
rect 8309 6409 8343 6443
rect 12265 6409 12299 6443
rect 12633 6409 12667 6443
rect 12817 6409 12851 6443
rect 14933 6409 14967 6443
rect 16497 6409 16531 6443
rect 17785 6409 17819 6443
rect 21327 6409 21361 6443
rect 22385 6409 22419 6443
rect 1547 6341 1581 6375
rect 6423 6341 6457 6375
rect 2145 6273 2179 6307
rect 3525 6273 3559 6307
rect 5917 6273 5951 6307
rect 7389 6273 7423 6307
rect 11897 6273 11931 6307
rect 1476 6205 1510 6239
rect 1685 6205 1719 6239
rect 4880 6205 4914 6239
rect 5457 6205 5491 6239
rect 5641 6205 5675 6239
rect 6320 6205 6354 6239
rect 6904 6205 6938 6239
rect 8585 6205 8619 6239
rect 8953 6205 8987 6239
rect 14565 6341 14599 6375
rect 19073 6341 19107 6375
rect 19257 6341 19291 6375
rect 20269 6341 20303 6375
rect 20913 6341 20947 6375
rect 21649 6341 21683 6375
rect 22017 6341 22051 6375
rect 15117 6205 15151 6239
rect 16932 6205 16966 6239
rect 18797 6205 18831 6239
rect 2466 6137 2500 6171
rect 3249 6137 3283 6171
rect 3341 6137 3375 6171
rect 4077 6137 4111 6171
rect 4169 6137 4203 6171
rect 4721 6137 4755 6171
rect 7751 6137 7785 6171
rect 9229 6137 9263 6171
rect 9321 6137 9355 6171
rect 9873 6137 9907 6171
rect 10885 6137 10919 6171
rect 10977 6137 11011 6171
rect 11529 6137 11563 6171
rect 12817 6137 12851 6171
rect 13001 6137 13035 6171
rect 13093 6137 13127 6171
rect 13645 6137 13679 6171
rect 15479 6137 15513 6171
rect 17417 6137 17451 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 21224 6205 21258 6239
rect 19717 6137 19751 6171
rect 19809 6137 19843 6171
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 13921 6069 13955 6103
rect 16037 6069 16071 6103
rect 17003 6069 17037 6103
rect 19257 6069 19291 6103
rect 19441 6069 19475 6103
rect 2329 5865 2363 5899
rect 8125 5865 8159 5899
rect 9045 5865 9079 5899
rect 9229 5865 9263 5899
rect 14565 5865 14599 5899
rect 14933 5865 14967 5899
rect 16589 5865 16623 5899
rect 16865 5865 16899 5899
rect 18153 5865 18187 5899
rect 19809 5865 19843 5899
rect 21925 5865 21959 5899
rect 1771 5797 1805 5831
rect 4353 5797 4387 5831
rect 5457 5797 5491 5831
rect 6009 5797 6043 5831
rect 6285 5797 6319 5831
rect 2697 5729 2731 5763
rect 2973 5729 3007 5763
rect 3249 5729 3283 5763
rect 3755 5729 3789 5763
rect 5064 5729 5098 5763
rect 6837 5729 6871 5763
rect 7297 5729 7331 5763
rect 7573 5729 7607 5763
rect 7757 5729 7791 5763
rect 8585 5729 8619 5763
rect 1409 5661 1443 5695
rect 3157 5661 3191 5695
rect 4261 5661 4295 5695
rect 5365 5661 5399 5695
rect 6193 5661 6227 5695
rect 9229 5661 9263 5695
rect 9321 5797 9355 5831
rect 9413 5797 9447 5831
rect 9781 5797 9815 5831
rect 9873 5797 9907 5831
rect 10425 5797 10459 5831
rect 10793 5797 10827 5831
rect 11161 5797 11195 5831
rect 11799 5797 11833 5831
rect 12725 5797 12759 5831
rect 13369 5797 13403 5831
rect 15669 5797 15703 5831
rect 17233 5797 17267 5831
rect 18975 5797 19009 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 3387 5593 3421 5627
rect 4813 5593 4847 5627
rect 8723 5593 8757 5627
rect 12357 5729 12391 5763
rect 13921 5729 13955 5763
rect 16221 5729 16255 5763
rect 20177 5729 20211 5763
rect 11437 5661 11471 5695
rect 13277 5661 13311 5695
rect 15577 5661 15611 5695
rect 17141 5661 17175 5695
rect 18613 5661 18647 5695
rect 21005 5661 21039 5695
rect 13001 5593 13035 5627
rect 17693 5593 17727 5627
rect 22293 5593 22327 5627
rect 3847 5525 3881 5559
rect 5135 5525 5169 5559
rect 8401 5525 8435 5559
rect 9321 5525 9355 5559
rect 14197 5525 14231 5559
rect 18429 5525 18463 5559
rect 19533 5525 19567 5559
rect 20545 5525 20579 5559
rect 2329 5321 2363 5355
rect 11483 5321 11517 5355
rect 13461 5321 13495 5355
rect 14013 5321 14047 5355
rect 14197 5321 14231 5355
rect 16497 5321 16531 5355
rect 19993 5321 20027 5355
rect 3525 5253 3559 5287
rect 6561 5253 6595 5287
rect 9045 5253 9079 5287
rect 11805 5253 11839 5287
rect 13783 5253 13817 5287
rect 1409 5185 1443 5219
rect 4997 5185 5031 5219
rect 7849 5185 7883 5219
rect 9689 5185 9723 5219
rect 10333 5185 10367 5219
rect 13185 5185 13219 5219
rect 17785 5253 17819 5287
rect 18199 5253 18233 5287
rect 18981 5253 19015 5287
rect 20269 5253 20303 5287
rect 21327 5253 21361 5287
rect 14749 5185 14783 5219
rect 2421 5117 2455 5151
rect 3525 5117 3559 5151
rect 3985 5117 4019 5151
rect 4445 5117 4479 5151
rect 4813 5117 4847 5151
rect 7573 5117 7607 5151
rect 8769 5117 8803 5151
rect 11380 5117 11414 5151
rect 12700 5117 12734 5151
rect 13712 5117 13746 5151
rect 14013 5117 14047 5151
rect 15393 5117 15427 5151
rect 15485 5117 15519 5151
rect 15669 5117 15703 5151
rect 16037 5117 16071 5151
rect 16865 5117 16899 5151
rect 18096 5117 18130 5151
rect 18521 5117 18555 5151
rect 19073 5117 19107 5151
rect 21256 5117 21290 5151
rect 21649 5117 21683 5151
rect 5181 5049 5215 5083
rect 5273 5049 5307 5083
rect 5825 5049 5859 5083
rect 6009 5049 6043 5083
rect 6101 5049 6135 5083
rect 6929 5049 6963 5083
rect 7021 5049 7055 5083
rect 9781 5049 9815 5083
rect 14473 5049 14507 5083
rect 14841 5049 14875 5083
rect 2789 4981 2823 5015
rect 3341 4981 3375 5015
rect 8217 4981 8251 5015
rect 9413 4981 9447 5015
rect 10701 4981 10735 5015
rect 11069 4981 11103 5015
rect 12265 4981 12299 5015
rect 12771 4981 12805 5015
rect 14013 4981 14047 5015
rect 17003 5049 17037 5083
rect 18337 5049 18371 5083
rect 19394 5049 19428 5083
rect 15577 4981 15611 5015
rect 17417 4981 17451 5015
rect 20913 4981 20947 5015
rect 22017 4981 22051 5015
rect 22385 4981 22419 5015
rect 1777 4777 1811 4811
rect 2329 4777 2363 4811
rect 5549 4777 5583 4811
rect 14289 4777 14323 4811
rect 17785 4777 17819 4811
rect 21925 4777 21959 4811
rect 2742 4709 2776 4743
rect 3652 4709 3686 4743
rect 5917 4709 5951 4743
rect 6653 4709 6687 4743
rect 6745 4709 6779 4743
rect 7573 4709 7607 4743
rect 8125 4709 8159 4743
rect 8401 4709 8435 4743
rect 9873 4709 9907 4743
rect 11799 4709 11833 4743
rect 13277 4709 13311 4743
rect 13369 4709 13403 4743
rect 16542 4709 16576 4743
rect 21097 4709 21131 4743
rect 21649 4709 21683 4743
rect 2421 4641 2455 4675
rect 3433 4641 3467 4675
rect 3776 4641 3810 4675
rect 4353 4641 4387 4675
rect 4537 4641 4571 4675
rect 4905 4641 4939 4675
rect 5052 4641 5086 4675
rect 8953 4641 8987 4675
rect 11437 4641 11471 4675
rect 12357 4641 12391 4675
rect 13921 4641 13955 4675
rect 16221 4641 16255 4675
rect 17141 4641 17175 4675
rect 19763 4641 19797 4675
rect 19855 4641 19889 4675
rect 20177 4641 20211 4675
rect 20545 4641 20579 4675
rect 21741 4641 21775 4675
rect 22293 4641 22327 4675
rect 1409 4573 1443 4607
rect 4629 4573 4663 4607
rect 5273 4573 5307 4607
rect 5825 4573 5859 4607
rect 6193 4573 6227 4607
rect 7481 4573 7515 4607
rect 8309 4573 8343 4607
rect 9229 4573 9263 4607
rect 9781 4573 9815 4607
rect 11161 4573 11195 4607
rect 15577 4573 15611 4607
rect 16037 4573 16071 4607
rect 17417 4573 17451 4607
rect 17969 4573 18003 4607
rect 19165 4573 19199 4607
rect 21005 4573 21039 4607
rect 3341 4505 3375 4539
rect 7205 4505 7239 4539
rect 10333 4505 10367 4539
rect 14565 4505 14599 4539
rect 14933 4505 14967 4539
rect 18889 4505 18923 4539
rect 19533 4505 19567 4539
rect 3847 4437 3881 4471
rect 5181 4437 5215 4471
rect 10701 4437 10735 4471
rect 12725 4437 12759 4471
rect 13093 4437 13127 4471
rect 15853 4437 15887 4471
rect 16037 4437 16071 4471
rect 21741 4437 21775 4471
rect 2421 4233 2455 4267
rect 4905 4233 4939 4267
rect 6101 4233 6135 4267
rect 11483 4233 11517 4267
rect 15255 4233 15289 4267
rect 16037 4233 16071 4267
rect 17877 4233 17911 4267
rect 20913 4233 20947 4267
rect 22385 4233 22419 4267
rect 2697 4165 2731 4199
rect 4399 4165 4433 4199
rect 4721 4165 4755 4199
rect 1501 4097 1535 4131
rect 2513 4029 2547 4063
rect 2881 4029 2915 4063
rect 3249 4029 3283 4063
rect 4296 4029 4330 4063
rect 4537 4029 4571 4063
rect 8309 4165 8343 4199
rect 11805 4165 11839 4199
rect 12587 4165 12621 4199
rect 14841 4165 14875 4199
rect 19257 4165 19291 4199
rect 7757 4097 7791 4131
rect 9229 4097 9263 4131
rect 10057 4097 10091 4131
rect 10241 4097 10275 4131
rect 13369 4097 13403 4131
rect 14565 4097 14599 4131
rect 17417 4097 17451 4131
rect 18429 4097 18463 4131
rect 4997 4029 5031 4063
rect 6076 4029 6110 4063
rect 6336 4029 6370 4063
rect 6837 4029 6871 4063
rect 7297 4029 7331 4063
rect 11380 4029 11414 4063
rect 12516 4029 12550 4063
rect 12909 4029 12943 4063
rect 15152 4029 15186 4063
rect 15577 4029 15611 4063
rect 16865 4029 16899 4063
rect 19993 4097 20027 4131
rect 21224 4029 21258 4063
rect 21649 4029 21683 4063
rect 3571 3961 3605 3995
rect 4905 3961 4939 3995
rect 7849 3961 7883 3995
rect 8585 3961 8619 3995
rect 8677 3961 8711 3995
rect 9413 3961 9447 3995
rect 9505 3961 9539 3995
rect 10333 3961 10367 3995
rect 10885 3961 10919 3995
rect 13553 3961 13587 3995
rect 13645 3961 13679 3995
rect 14197 3961 14231 3995
rect 16221 3961 16255 3995
rect 16313 3961 16347 3995
rect 18153 3961 18187 3995
rect 18245 3961 18279 3995
rect 19257 3961 19291 3995
rect 19717 3961 19751 3995
rect 19809 3961 19843 3995
rect 1869 3893 1903 3927
rect 4169 3893 4203 3927
rect 5365 3893 5399 3927
rect 5917 3893 5951 3927
rect 6423 3893 6457 3927
rect 6929 3893 6963 3927
rect 11161 3893 11195 3927
rect 12265 3893 12299 3927
rect 19073 3893 19107 3927
rect 19533 3893 19567 3927
rect 21327 3893 21361 3927
rect 22017 3893 22051 3927
rect 1777 3689 1811 3723
rect 3433 3689 3467 3723
rect 4537 3689 4571 3723
rect 5089 3689 5123 3723
rect 6101 3689 6135 3723
rect 8217 3689 8251 3723
rect 10195 3689 10229 3723
rect 10793 3689 10827 3723
rect 11345 3689 11379 3723
rect 13001 3689 13035 3723
rect 14473 3689 14507 3723
rect 14749 3689 14783 3723
rect 15485 3689 15519 3723
rect 15991 3689 16025 3723
rect 17785 3689 17819 3723
rect 17877 3689 17911 3723
rect 19165 3689 19199 3723
rect 19717 3689 19751 3723
rect 20545 3689 20579 3723
rect 21925 3689 21959 3723
rect 2742 3621 2776 3655
rect 5502 3621 5536 3655
rect 6377 3621 6411 3655
rect 7659 3621 7693 3655
rect 8401 3621 8435 3655
rect 8502 3621 8536 3655
rect 9275 3621 9309 3655
rect 12311 3621 12345 3655
rect 13547 3621 13581 3655
rect 16405 3621 16439 3655
rect 16497 3621 16531 3655
rect 17186 3621 17220 3655
rect 1409 3553 1443 3587
rect 3341 3553 3375 3587
rect 3776 3553 3810 3587
rect 5181 3553 5215 3587
rect 6929 3553 6963 3587
rect 9137 3553 9171 3587
rect 9724 3553 9758 3587
rect 10092 3553 10126 3587
rect 12224 3553 12258 3587
rect 12725 3553 12759 3587
rect 14105 3553 14139 3587
rect 15920 3553 15954 3587
rect 16681 3553 16715 3587
rect 2421 3485 2455 3519
rect 6285 3485 6319 3519
rect 7021 3485 7055 3519
rect 7297 3485 7331 3519
rect 10421 3485 10455 3519
rect 13185 3485 13219 3519
rect 16497 3485 16531 3519
rect 16865 3485 16899 3519
rect 4077 3417 4111 3451
rect 8953 3417 8987 3451
rect 11989 3417 12023 3451
rect 18521 3621 18555 3655
rect 21097 3621 21131 3655
rect 18613 3553 18647 3587
rect 20269 3553 20303 3587
rect 21005 3485 21039 3519
rect 21281 3485 21315 3519
rect 18797 3417 18831 3451
rect 2329 3349 2363 3383
rect 3847 3349 3881 3383
rect 9827 3349 9861 3383
rect 11713 3349 11747 3383
rect 17877 3349 17911 3383
rect 18061 3349 18095 3383
rect 19533 3349 19567 3383
rect 22293 3349 22327 3383
rect 949 3145 983 3179
rect 4353 3145 4387 3179
rect 11943 3145 11977 3179
rect 12219 3145 12253 3179
rect 12587 3145 12621 3179
rect 17785 3145 17819 3179
rect 21741 3145 21775 3179
rect 6377 3077 6411 3111
rect 9965 3077 9999 3111
rect 13277 3077 13311 3111
rect 15669 3077 15703 3111
rect 17049 3077 17083 3111
rect 1409 3009 1443 3043
rect 3433 3009 3467 3043
rect 4445 3009 4479 3043
rect 7757 3009 7791 3043
rect 8401 3009 8435 3043
rect 8585 3009 8619 3043
rect 9229 3009 9263 3043
rect 10241 3009 10275 3043
rect 10885 3009 10919 3043
rect 11069 3009 11103 3043
rect 14565 3009 14599 3043
rect 14933 3009 14967 3043
rect 17509 3009 17543 3043
rect 18429 3009 18463 3043
rect 19441 3009 19475 3043
rect 19717 3009 19751 3043
rect 19993 3009 20027 3043
rect 2421 2941 2455 2975
rect 5457 2941 5491 2975
rect 6469 2941 6503 2975
rect 6929 2941 6963 2975
rect 7297 2941 7331 2975
rect 7573 2941 7607 2975
rect 11840 2941 11874 2975
rect 12081 2941 12115 2975
rect 12484 2941 12518 2975
rect 12909 2941 12943 2975
rect 14197 2941 14231 2975
rect 16129 2941 16163 2975
rect 16865 2941 16899 2975
rect 21189 2941 21223 2975
rect 3754 2873 3788 2907
rect 4766 2873 4800 2907
rect 5733 2873 5767 2907
rect 7849 2873 7883 2907
rect 8654 2873 8688 2907
rect 9402 2873 9436 2907
rect 9505 2873 9539 2907
rect 10333 2873 10367 2907
rect 11161 2873 11195 2907
rect 11713 2873 11747 2907
rect 13553 2873 13587 2907
rect 13645 2873 13679 2907
rect 15117 2873 15151 2907
rect 15209 2873 15243 2907
rect 18153 2873 18187 2907
rect 18245 2873 18279 2907
rect 19809 2873 19843 2907
rect 22109 2873 22143 2907
rect 1777 2805 1811 2839
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 3341 2805 3375 2839
rect 5365 2805 5399 2839
rect 6607 2805 6641 2839
rect 16773 2805 16807 2839
rect 19073 2805 19107 2839
rect 20637 2805 20671 2839
rect 21005 2805 21039 2839
rect 21373 2805 21407 2839
rect 581 2601 615 2635
rect 2329 2601 2363 2635
rect 3617 2601 3651 2635
rect 7849 2601 7883 2635
rect 14013 2601 14047 2635
rect 15025 2601 15059 2635
rect 17693 2601 17727 2635
rect 21373 2601 21407 2635
rect 22109 2601 22143 2635
rect 1771 2533 1805 2567
rect 2742 2533 2776 2567
rect 4398 2533 4432 2567
rect 5410 2533 5444 2567
rect 7250 2533 7284 2567
rect 8125 2533 8159 2567
rect 8861 2533 8895 2567
rect 8953 2533 8987 2567
rect 9505 2533 9539 2567
rect 9873 2533 9907 2567
rect 9965 2533 9999 2567
rect 10793 2533 10827 2567
rect 11345 2533 11379 2567
rect 11621 2533 11655 2567
rect 12817 2533 12851 2567
rect 16031 2533 16065 2567
rect 17969 2533 18003 2567
rect 18429 2533 18463 2567
rect 18521 2533 18555 2567
rect 19349 2533 19383 2567
rect 1409 2465 1443 2499
rect 3433 2465 3467 2499
rect 4077 2465 4111 2499
rect 6101 2465 6135 2499
rect 6494 2465 6528 2499
rect 6929 2465 6963 2499
rect 12311 2465 12345 2499
rect 13645 2465 13679 2499
rect 14264 2465 14298 2499
rect 16589 2465 16623 2499
rect 19073 2465 19107 2499
rect 19901 2465 19935 2499
rect 21189 2465 21223 2499
rect 2421 2397 2455 2431
rect 5089 2397 5123 2431
rect 8033 2397 8067 2431
rect 8677 2397 8711 2431
rect 10149 2397 10183 2431
rect 10701 2397 10735 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 12725 2397 12759 2431
rect 15669 2397 15703 2431
rect 17049 2397 17083 2431
rect 17233 2397 17267 2431
rect 19533 2397 19567 2431
rect 20453 2397 20487 2431
rect 3341 2329 3375 2363
rect 6009 2329 6043 2363
rect 6653 2329 6687 2363
rect 13277 2329 13311 2363
rect 16865 2329 16899 2363
rect 4997 2261 5031 2295
rect 6285 2261 6319 2295
rect 12403 2261 12437 2295
rect 14473 2261 14507 2295
rect 14749 2261 14783 2295
rect 17049 2261 17083 2295
rect 20821 2329 20855 2363
rect 19533 2261 19567 2295
rect 19717 2261 19751 2295
rect 20085 2261 20119 2295
rect 21741 2261 21775 2295
rect 121 85 155 119
<< metal1 >>
rect 2866 23536 2872 23588
rect 2924 23576 2930 23588
rect 8941 23579 8999 23585
rect 8941 23576 8953 23579
rect 2924 23548 8953 23576
rect 2924 23536 2930 23548
rect 8941 23545 8953 23548
rect 8987 23545 8999 23579
rect 8941 23539 8999 23545
rect 15102 23536 15108 23588
rect 15160 23576 15166 23588
rect 19334 23576 19340 23588
rect 15160 23548 19340 23576
rect 15160 23536 15166 23548
rect 19334 23536 19340 23548
rect 19392 23536 19398 23588
rect 569 23239 627 23245
rect 569 23205 581 23239
rect 615 23236 627 23239
rect 8849 23239 8907 23245
rect 8849 23236 8861 23239
rect 615 23208 8861 23236
rect 615 23205 627 23208
rect 569 23199 627 23205
rect 8849 23205 8861 23208
rect 8895 23205 8907 23239
rect 8849 23199 8907 23205
rect 3694 23128 3700 23180
rect 3752 23168 3758 23180
rect 9582 23168 9588 23180
rect 3752 23140 9588 23168
rect 3752 23128 3758 23140
rect 9582 23128 9588 23140
rect 9640 23128 9646 23180
rect 937 23103 995 23109
rect 937 23069 949 23103
rect 983 23100 995 23103
rect 7745 23103 7803 23109
rect 7745 23100 7757 23103
rect 983 23072 7757 23100
rect 983 23069 995 23072
rect 937 23063 995 23069
rect 7745 23069 7757 23072
rect 7791 23069 7803 23103
rect 7745 23063 7803 23069
rect 2222 22992 2228 23044
rect 2280 23032 2286 23044
rect 7190 23032 7196 23044
rect 2280 23004 7196 23032
rect 2280 22992 2286 23004
rect 7190 22992 7196 23004
rect 7248 22992 7254 23044
rect 7377 23035 7435 23041
rect 7377 23001 7389 23035
rect 7423 23032 7435 23035
rect 14734 23032 14740 23044
rect 7423 23004 14740 23032
rect 7423 23001 7435 23004
rect 7377 22995 7435 23001
rect 14734 22992 14740 23004
rect 14792 22992 14798 23044
rect 566 22924 572 22976
rect 624 22964 630 22976
rect 9033 22967 9091 22973
rect 9033 22964 9045 22967
rect 624 22936 9045 22964
rect 624 22924 630 22936
rect 9033 22933 9045 22936
rect 9079 22933 9091 22967
rect 9033 22927 9091 22933
rect 1118 22856 1124 22908
rect 1176 22896 1182 22908
rect 8021 22899 8079 22905
rect 8021 22896 8033 22899
rect 1176 22868 8033 22896
rect 1176 22856 1182 22868
rect 8021 22865 8033 22868
rect 8067 22865 8079 22899
rect 8021 22859 8079 22865
rect 8941 22899 8999 22905
rect 8941 22865 8953 22899
rect 8987 22896 8999 22899
rect 19150 22896 19156 22908
rect 8987 22868 19156 22896
rect 8987 22865 8999 22868
rect 8941 22859 8999 22865
rect 19150 22856 19156 22868
rect 19208 22856 19214 22908
rect 934 22788 940 22840
rect 992 22828 998 22840
rect 7558 22828 7564 22840
rect 992 22800 7564 22828
rect 992 22788 998 22800
rect 7558 22788 7564 22800
rect 7616 22788 7622 22840
rect 7650 22788 7656 22840
rect 7708 22828 7714 22840
rect 19242 22828 19248 22840
rect 7708 22800 19248 22828
rect 7708 22788 7714 22800
rect 19242 22788 19248 22800
rect 19300 22788 19306 22840
rect 2038 22720 2044 22772
rect 2096 22760 2102 22772
rect 8662 22760 8668 22772
rect 2096 22732 8668 22760
rect 2096 22720 2102 22732
rect 8662 22720 8668 22732
rect 8720 22720 8726 22772
rect 9950 22720 9956 22772
rect 10008 22760 10014 22772
rect 19334 22760 19340 22772
rect 10008 22732 19340 22760
rect 10008 22720 10014 22732
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 1854 22652 1860 22704
rect 1912 22692 1918 22704
rect 17954 22692 17960 22704
rect 1912 22664 17960 22692
rect 1912 22652 1918 22664
rect 17954 22652 17960 22664
rect 18012 22652 18018 22704
rect 1946 22584 1952 22636
rect 2004 22624 2010 22636
rect 6273 22627 6331 22633
rect 6273 22624 6285 22627
rect 2004 22596 6285 22624
rect 2004 22584 2010 22596
rect 6273 22593 6285 22596
rect 6319 22593 6331 22627
rect 6273 22587 6331 22593
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22624 8907 22627
rect 16206 22624 16212 22636
rect 8895 22596 16212 22624
rect 8895 22593 8907 22596
rect 8849 22587 8907 22593
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 1486 22516 1492 22568
rect 1544 22556 1550 22568
rect 6089 22559 6147 22565
rect 6089 22556 6101 22559
rect 1544 22528 6101 22556
rect 1544 22516 1550 22528
rect 6089 22525 6101 22528
rect 6135 22525 6147 22559
rect 6089 22519 6147 22525
rect 6181 22559 6239 22565
rect 6181 22525 6193 22559
rect 6227 22556 6239 22559
rect 13630 22556 13636 22568
rect 6227 22528 13636 22556
rect 6227 22525 6239 22528
rect 6181 22519 6239 22525
rect 13630 22516 13636 22528
rect 13688 22516 13694 22568
rect 17 22491 75 22497
rect 17 22457 29 22491
rect 63 22488 75 22491
rect 14274 22488 14280 22500
rect 63 22460 14280 22488
rect 63 22457 75 22460
rect 17 22451 75 22457
rect 14274 22448 14280 22460
rect 14332 22448 14338 22500
rect 477 22423 535 22429
rect 477 22389 489 22423
rect 523 22420 535 22423
rect 5077 22423 5135 22429
rect 5077 22420 5089 22423
rect 523 22392 5089 22420
rect 523 22389 535 22392
rect 477 22383 535 22389
rect 5077 22389 5089 22392
rect 5123 22389 5135 22423
rect 5077 22383 5135 22389
rect 6089 22423 6147 22429
rect 6089 22389 6101 22423
rect 6135 22420 6147 22423
rect 9214 22420 9220 22432
rect 6135 22392 9220 22420
rect 6135 22389 6147 22392
rect 6089 22383 6147 22389
rect 9214 22380 9220 22392
rect 9272 22380 9278 22432
rect 3694 22312 3700 22364
rect 3752 22352 3758 22364
rect 7834 22352 7840 22364
rect 3752 22324 7840 22352
rect 3752 22312 3758 22324
rect 7834 22312 7840 22324
rect 7892 22312 7898 22364
rect 8018 22312 8024 22364
rect 8076 22352 8082 22364
rect 11057 22355 11115 22361
rect 11057 22352 11069 22355
rect 8076 22324 11069 22352
rect 8076 22312 8082 22324
rect 11057 22321 11069 22324
rect 11103 22321 11115 22355
rect 11057 22315 11115 22321
rect 3234 22244 3240 22296
rect 3292 22284 3298 22296
rect 6181 22287 6239 22293
rect 6181 22284 6193 22287
rect 3292 22256 6193 22284
rect 3292 22244 3298 22256
rect 6181 22253 6193 22256
rect 6227 22253 6239 22287
rect 6181 22247 6239 22253
rect 6273 22287 6331 22293
rect 6273 22253 6285 22287
rect 6319 22284 6331 22287
rect 9766 22284 9772 22296
rect 6319 22256 9772 22284
rect 6319 22253 6331 22256
rect 6273 22247 6331 22253
rect 9766 22244 9772 22256
rect 9824 22244 9830 22296
rect 10594 22244 10600 22296
rect 10652 22284 10658 22296
rect 15654 22284 15660 22296
rect 10652 22256 15660 22284
rect 10652 22244 10658 22256
rect 15654 22244 15660 22256
rect 15712 22244 15718 22296
rect 1026 22176 1032 22228
rect 1084 22216 1090 22228
rect 9033 22219 9091 22225
rect 1084 22188 7512 22216
rect 1084 22176 1090 22188
rect 4062 22108 4068 22160
rect 4120 22148 4126 22160
rect 7377 22151 7435 22157
rect 7377 22148 7389 22151
rect 4120 22120 7389 22148
rect 4120 22108 4126 22120
rect 7377 22117 7389 22120
rect 7423 22117 7435 22151
rect 7484 22148 7512 22188
rect 9033 22185 9045 22219
rect 9079 22216 9091 22219
rect 20898 22216 20904 22228
rect 9079 22188 20904 22216
rect 9079 22185 9091 22188
rect 9033 22179 9091 22185
rect 20898 22176 20904 22188
rect 20956 22176 20962 22228
rect 10962 22148 10968 22160
rect 7484 22120 10968 22148
rect 7377 22111 7435 22117
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 11057 22151 11115 22157
rect 11057 22117 11069 22151
rect 11103 22148 11115 22151
rect 16942 22148 16948 22160
rect 11103 22120 16948 22148
rect 11103 22117 11115 22120
rect 11057 22111 11115 22117
rect 16942 22108 16948 22120
rect 17000 22108 17006 22160
rect 8021 22083 8079 22089
rect 8021 22049 8033 22083
rect 8067 22080 8079 22083
rect 19058 22080 19064 22092
rect 8067 22052 19064 22080
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 22012 7803 22015
rect 20438 22012 20444 22024
rect 7791 21984 20444 22012
rect 7791 21981 7803 21984
rect 7745 21975 7803 21981
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 3878 21904 3884 21956
rect 3936 21944 3942 21956
rect 5534 21944 5540 21956
rect 3936 21916 5540 21944
rect 3936 21904 3942 21916
rect 5534 21904 5540 21916
rect 5592 21944 5598 21956
rect 18322 21944 18328 21956
rect 5592 21916 18328 21944
rect 5592 21904 5598 21916
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 2590 21836 2596 21888
rect 2648 21876 2654 21888
rect 4706 21876 4712 21888
rect 2648 21848 4712 21876
rect 2648 21836 2654 21848
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5077 21879 5135 21885
rect 5077 21845 5089 21879
rect 5123 21876 5135 21879
rect 15470 21876 15476 21888
rect 5123 21848 15476 21876
rect 5123 21845 5135 21848
rect 5077 21839 5135 21845
rect 15470 21836 15476 21848
rect 15528 21836 15534 21888
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 845 21675 903 21681
rect 845 21641 857 21675
rect 891 21672 903 21675
rect 2133 21675 2191 21681
rect 2133 21672 2145 21675
rect 891 21644 2145 21672
rect 891 21641 903 21644
rect 845 21635 903 21641
rect 2133 21641 2145 21644
rect 2179 21672 2191 21675
rect 2222 21672 2228 21684
rect 2179 21644 2228 21672
rect 2179 21641 2191 21644
rect 2133 21635 2191 21641
rect 2222 21632 2228 21644
rect 2280 21632 2286 21684
rect 3881 21675 3939 21681
rect 3881 21641 3893 21675
rect 3927 21672 3939 21675
rect 4430 21672 4436 21684
rect 3927 21644 4436 21672
rect 3927 21641 3939 21644
rect 3881 21635 3939 21641
rect 4430 21632 4436 21644
rect 4488 21672 4494 21684
rect 5902 21672 5908 21684
rect 4488 21644 5908 21672
rect 4488 21632 4494 21644
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 6638 21632 6644 21684
rect 6696 21672 6702 21684
rect 9585 21675 9643 21681
rect 6696 21644 7649 21672
rect 6696 21632 6702 21644
rect 3418 21564 3424 21616
rect 3476 21604 3482 21616
rect 4246 21613 4252 21616
rect 4230 21607 4252 21613
rect 4230 21604 4242 21607
rect 3476 21576 4242 21604
rect 3476 21564 3482 21576
rect 4230 21573 4242 21576
rect 4304 21604 4310 21616
rect 4341 21607 4399 21613
rect 4341 21604 4353 21607
rect 4304 21576 4353 21604
rect 4230 21567 4252 21573
rect 4246 21564 4252 21567
rect 4304 21564 4310 21576
rect 4341 21573 4353 21576
rect 4387 21573 4399 21607
rect 4341 21567 4399 21573
rect 4448 21604 4476 21632
rect 4448 21576 4660 21604
rect 4448 21545 4476 21576
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21536 2007 21539
rect 2501 21539 2559 21545
rect 2501 21536 2513 21539
rect 1995 21508 2513 21536
rect 1995 21505 2007 21508
rect 1949 21499 2007 21505
rect 2501 21505 2513 21508
rect 2547 21536 2559 21539
rect 4433 21539 4491 21545
rect 2547 21508 3924 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 2133 21471 2191 21477
rect 2133 21437 2145 21471
rect 2179 21468 2191 21471
rect 2409 21471 2467 21477
rect 2409 21468 2421 21471
rect 2179 21440 2421 21468
rect 2179 21437 2191 21440
rect 2133 21431 2191 21437
rect 2409 21437 2421 21440
rect 2455 21437 2467 21471
rect 2409 21431 2467 21437
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 1210 21360 1216 21412
rect 1268 21400 1274 21412
rect 2590 21400 2596 21412
rect 1268 21372 2596 21400
rect 1268 21360 1274 21372
rect 2590 21360 2596 21372
rect 2648 21400 2654 21412
rect 2700 21400 2728 21431
rect 3142 21400 3148 21412
rect 2648 21372 2728 21400
rect 3103 21372 3148 21400
rect 2648 21360 2654 21372
rect 3142 21360 3148 21372
rect 3200 21360 3206 21412
rect 1535 21335 1593 21341
rect 1535 21301 1547 21335
rect 1581 21332 1593 21335
rect 2130 21332 2136 21344
rect 1581 21304 2136 21332
rect 1581 21301 1593 21304
rect 1535 21295 1593 21301
rect 2130 21292 2136 21304
rect 2188 21292 2194 21344
rect 3418 21332 3424 21344
rect 3379 21304 3424 21332
rect 3418 21292 3424 21304
rect 3476 21292 3482 21344
rect 3896 21332 3924 21508
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 4632 21536 4660 21576
rect 4706 21564 4712 21616
rect 4764 21604 4770 21616
rect 6365 21607 6423 21613
rect 6365 21604 6377 21607
rect 4764 21576 6377 21604
rect 4764 21564 4770 21576
rect 6365 21573 6377 21576
rect 6411 21604 6423 21607
rect 7282 21604 7288 21616
rect 6411 21576 7288 21604
rect 6411 21573 6423 21576
rect 6365 21567 6423 21573
rect 7282 21564 7288 21576
rect 7340 21564 7346 21616
rect 7621 21604 7649 21644
rect 9585 21641 9597 21675
rect 9631 21672 9643 21675
rect 10042 21672 10048 21684
rect 9631 21644 10048 21672
rect 9631 21641 9643 21644
rect 9585 21635 9643 21641
rect 10042 21632 10048 21644
rect 10100 21632 10106 21684
rect 13633 21675 13691 21681
rect 13633 21672 13645 21675
rect 10152 21644 13645 21672
rect 10152 21604 10180 21644
rect 13633 21641 13645 21644
rect 13679 21641 13691 21675
rect 13633 21635 13691 21641
rect 14461 21675 14519 21681
rect 14461 21641 14473 21675
rect 14507 21672 14519 21675
rect 15378 21672 15384 21684
rect 14507 21644 15384 21672
rect 14507 21641 14519 21644
rect 14461 21635 14519 21641
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 16485 21675 16543 21681
rect 16485 21672 16497 21675
rect 15620 21644 16497 21672
rect 15620 21632 15626 21644
rect 16485 21641 16497 21644
rect 16531 21641 16543 21675
rect 16485 21635 16543 21641
rect 16669 21675 16727 21681
rect 16669 21641 16681 21675
rect 16715 21672 16727 21675
rect 18490 21675 18548 21681
rect 18490 21672 18502 21675
rect 16715 21644 18502 21672
rect 16715 21641 16727 21644
rect 16669 21635 16727 21641
rect 18490 21641 18502 21644
rect 18536 21672 18548 21675
rect 19337 21675 19395 21681
rect 19337 21672 19349 21675
rect 18536 21644 19349 21672
rect 18536 21641 18548 21644
rect 18490 21635 18548 21641
rect 19337 21641 19349 21644
rect 19383 21641 19395 21675
rect 19337 21635 19395 21641
rect 7621 21576 10180 21604
rect 10226 21564 10232 21616
rect 10284 21604 10290 21616
rect 11563 21607 11621 21613
rect 11563 21604 11575 21607
rect 10284 21576 11575 21604
rect 10284 21564 10290 21576
rect 11563 21573 11575 21576
rect 11609 21573 11621 21607
rect 11563 21567 11621 21573
rect 12526 21564 12532 21616
rect 12584 21604 12590 21616
rect 12894 21604 12900 21616
rect 12584 21576 12900 21604
rect 12584 21564 12590 21576
rect 12894 21564 12900 21576
rect 12952 21564 12958 21616
rect 13265 21607 13323 21613
rect 13265 21573 13277 21607
rect 13311 21604 13323 21607
rect 16117 21607 16175 21613
rect 16117 21604 16129 21607
rect 13311 21576 16129 21604
rect 13311 21573 13323 21576
rect 13265 21567 13323 21573
rect 16117 21573 16129 21576
rect 16163 21604 16175 21607
rect 18046 21604 18052 21616
rect 16163 21576 18052 21604
rect 16163 21573 16175 21576
rect 16117 21567 16175 21573
rect 18046 21564 18052 21576
rect 18104 21564 18110 21616
rect 18138 21564 18144 21616
rect 18196 21604 18202 21616
rect 18598 21604 18604 21616
rect 18196 21576 18368 21604
rect 18559 21576 18604 21604
rect 18196 21564 18202 21576
rect 4798 21536 4804 21548
rect 4632 21508 4804 21536
rect 4433 21499 4491 21505
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 6733 21539 6791 21545
rect 6733 21536 6745 21539
rect 5552 21508 6745 21536
rect 3970 21428 3976 21480
rect 4028 21468 4034 21480
rect 4065 21471 4123 21477
rect 4065 21468 4077 21471
rect 4028 21440 4077 21468
rect 4028 21428 4034 21440
rect 4065 21437 4077 21440
rect 4111 21437 4123 21471
rect 5552 21468 5580 21508
rect 6733 21505 6745 21508
rect 6779 21536 6791 21539
rect 7006 21536 7012 21548
rect 6779 21508 7012 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 18340 21536 18368 21576
rect 18598 21564 18604 21576
rect 18656 21564 18662 21616
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 9640 21508 18276 21536
rect 18340 21508 18705 21536
rect 9640 21496 9646 21508
rect 5664 21471 5722 21477
rect 5664 21468 5676 21471
rect 4065 21431 4123 21437
rect 4595 21440 5580 21468
rect 4595 21332 4623 21440
rect 5644 21437 5676 21468
rect 5710 21437 5722 21471
rect 5644 21431 5722 21437
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 7282 21468 7288 21480
rect 7239 21440 7288 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 5644 21400 5672 21431
rect 5460 21372 5672 21400
rect 5460 21344 5488 21372
rect 6840 21344 6868 21431
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 7653 21471 7711 21477
rect 7653 21437 7665 21471
rect 7699 21468 7711 21471
rect 7834 21468 7840 21480
rect 7699 21440 7840 21468
rect 7699 21437 7711 21440
rect 7653 21431 7711 21437
rect 7834 21428 7840 21440
rect 7892 21428 7898 21480
rect 8570 21428 8576 21480
rect 8628 21468 8634 21480
rect 8700 21471 8758 21477
rect 8700 21468 8712 21471
rect 8628 21440 8712 21468
rect 8628 21428 8634 21440
rect 8700 21437 8712 21440
rect 8746 21468 8758 21471
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8746 21440 9137 21468
rect 8746 21437 8758 21440
rect 8700 21431 8758 21437
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 10042 21468 10048 21480
rect 10003 21440 10048 21468
rect 9125 21431 9183 21437
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 10321 21471 10379 21477
rect 10321 21437 10333 21471
rect 10367 21437 10379 21471
rect 10321 21431 10379 21437
rect 7098 21360 7104 21412
rect 7156 21400 7162 21412
rect 8297 21403 8355 21409
rect 8297 21400 8309 21403
rect 7156 21372 8309 21400
rect 7156 21360 7162 21372
rect 8297 21369 8309 21372
rect 8343 21369 8355 21403
rect 8297 21363 8355 21369
rect 8803 21403 8861 21409
rect 8803 21369 8815 21403
rect 8849 21400 8861 21403
rect 9306 21400 9312 21412
rect 8849 21372 9312 21400
rect 8849 21369 8861 21372
rect 8803 21363 8861 21369
rect 9306 21360 9312 21372
rect 9364 21360 9370 21412
rect 9398 21360 9404 21412
rect 9456 21400 9462 21412
rect 10336 21400 10364 21431
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 11460 21471 11518 21477
rect 11460 21468 11472 21471
rect 10468 21440 11472 21468
rect 10468 21428 10474 21440
rect 11460 21437 11472 21440
rect 11506 21468 11518 21471
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 11506 21440 11897 21468
rect 11506 21437 11518 21440
rect 11460 21431 11518 21437
rect 11885 21437 11897 21440
rect 11931 21468 11943 21471
rect 12158 21468 12164 21480
rect 11931 21440 12164 21468
rect 11931 21437 11943 21440
rect 11885 21431 11943 21437
rect 12158 21428 12164 21440
rect 12216 21428 12222 21480
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21468 14335 21471
rect 17072 21471 17130 21477
rect 17072 21468 17084 21471
rect 14323 21440 14964 21468
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 9456 21372 9771 21400
rect 10336 21372 10916 21400
rect 9456 21360 9462 21372
rect 4706 21332 4712 21344
rect 3896 21304 4623 21332
rect 4667 21304 4712 21332
rect 4706 21292 4712 21304
rect 4764 21292 4770 21344
rect 5074 21332 5080 21344
rect 5035 21304 5080 21332
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 5442 21332 5448 21344
rect 5403 21304 5448 21332
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 5767 21335 5825 21341
rect 5767 21301 5779 21335
rect 5813 21332 5825 21335
rect 5994 21332 6000 21344
rect 5813 21304 6000 21332
rect 5813 21301 5825 21304
rect 5767 21295 5825 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 6822 21332 6828 21344
rect 6735 21304 6828 21332
rect 6822 21292 6828 21304
rect 6880 21332 6886 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 6880 21304 8033 21332
rect 6880 21292 6886 21304
rect 8021 21301 8033 21304
rect 8067 21332 8079 21335
rect 8110 21332 8116 21344
rect 8067 21304 8116 21332
rect 8067 21301 8079 21304
rect 8021 21295 8079 21301
rect 8110 21292 8116 21304
rect 8168 21292 8174 21344
rect 9743 21332 9771 21372
rect 10888 21341 10916 21372
rect 11238 21360 11244 21412
rect 11296 21400 11302 21412
rect 12345 21403 12403 21409
rect 12345 21400 12357 21403
rect 11296 21372 12357 21400
rect 11296 21360 11302 21372
rect 12345 21369 12357 21372
rect 12391 21400 12403 21403
rect 12526 21400 12532 21412
rect 12391 21372 12532 21400
rect 12391 21369 12403 21372
rect 12345 21363 12403 21369
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 12710 21360 12716 21412
rect 12768 21400 12774 21412
rect 12805 21403 12863 21409
rect 12805 21400 12817 21403
rect 12768 21372 12817 21400
rect 12768 21360 12774 21372
rect 12805 21369 12817 21372
rect 12851 21400 12863 21403
rect 12894 21400 12900 21412
rect 12851 21372 12900 21400
rect 12851 21369 12863 21372
rect 12805 21363 12863 21369
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 9861 21335 9919 21341
rect 9861 21332 9873 21335
rect 9743 21304 9873 21332
rect 9861 21301 9873 21304
rect 9907 21301 9919 21335
rect 9861 21295 9919 21301
rect 10873 21335 10931 21341
rect 10873 21301 10885 21335
rect 10919 21332 10931 21335
rect 11054 21332 11060 21344
rect 10919 21304 11060 21332
rect 10919 21301 10931 21304
rect 10873 21295 10931 21301
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 11330 21292 11336 21344
rect 11388 21332 11394 21344
rect 14936 21341 14964 21440
rect 16868 21440 17084 21468
rect 15010 21360 15016 21412
rect 15068 21400 15074 21412
rect 15197 21403 15255 21409
rect 15197 21400 15209 21403
rect 15068 21372 15209 21400
rect 15068 21360 15074 21372
rect 15197 21369 15209 21372
rect 15243 21369 15255 21403
rect 15562 21400 15568 21412
rect 15523 21372 15568 21400
rect 15197 21363 15255 21369
rect 15562 21360 15568 21372
rect 15620 21360 15626 21412
rect 15657 21403 15715 21409
rect 15657 21369 15669 21403
rect 15703 21400 15715 21403
rect 15746 21400 15752 21412
rect 15703 21372 15752 21400
rect 15703 21369 15715 21372
rect 15657 21363 15715 21369
rect 15746 21360 15752 21372
rect 15804 21360 15810 21412
rect 14921 21335 14979 21341
rect 11388 21304 11433 21332
rect 11388 21292 11394 21304
rect 14921 21301 14933 21335
rect 14967 21332 14979 21335
rect 15102 21332 15108 21344
rect 14967 21304 15108 21332
rect 14967 21301 14979 21304
rect 14921 21295 14979 21301
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 16080 21304 16681 21332
rect 16080 21292 16086 21304
rect 16669 21301 16681 21304
rect 16715 21301 16727 21335
rect 16669 21295 16727 21301
rect 16758 21292 16764 21344
rect 16816 21332 16822 21344
rect 16868 21341 16896 21440
rect 17072 21437 17084 21440
rect 17118 21437 17130 21471
rect 17770 21468 17776 21480
rect 17683 21440 17776 21468
rect 17072 21431 17130 21437
rect 17770 21428 17776 21440
rect 17828 21468 17834 21480
rect 18138 21468 18144 21480
rect 17828 21440 18144 21468
rect 17828 21428 17834 21440
rect 18138 21428 18144 21440
rect 18196 21428 18202 21480
rect 18248 21468 18276 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18782 21496 18788 21548
rect 18840 21536 18846 21548
rect 21315 21539 21373 21545
rect 21315 21536 21327 21539
rect 18840 21508 21327 21536
rect 18840 21496 18846 21508
rect 21315 21505 21327 21508
rect 21361 21505 21373 21539
rect 21315 21499 21373 21505
rect 19924 21471 19982 21477
rect 19924 21468 19936 21471
rect 18248 21440 19936 21468
rect 19924 21437 19936 21440
rect 19970 21468 19982 21471
rect 20349 21471 20407 21477
rect 20349 21468 20361 21471
rect 19970 21440 20361 21468
rect 19970 21437 19982 21440
rect 19924 21431 19982 21437
rect 20349 21437 20361 21440
rect 20395 21437 20407 21471
rect 20349 21431 20407 21437
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 21212 21471 21270 21477
rect 21212 21468 21224 21471
rect 20772 21440 21224 21468
rect 20772 21428 20778 21440
rect 21212 21437 21224 21440
rect 21258 21468 21270 21471
rect 21637 21471 21695 21477
rect 21637 21468 21649 21471
rect 21258 21440 21649 21468
rect 21258 21437 21270 21440
rect 21212 21431 21270 21437
rect 21637 21437 21649 21440
rect 21683 21437 21695 21471
rect 21637 21431 21695 21437
rect 16942 21360 16948 21412
rect 17000 21400 17006 21412
rect 17175 21403 17233 21409
rect 17175 21400 17187 21403
rect 17000 21372 17187 21400
rect 17000 21360 17006 21372
rect 17175 21369 17187 21372
rect 17221 21369 17233 21403
rect 18322 21400 18328 21412
rect 18283 21372 18328 21400
rect 17175 21363 17233 21369
rect 18322 21360 18328 21372
rect 18380 21400 18386 21412
rect 19705 21403 19763 21409
rect 19705 21400 19717 21403
rect 18380 21372 19717 21400
rect 18380 21360 18386 21372
rect 19705 21369 19717 21372
rect 19751 21369 19763 21403
rect 19705 21363 19763 21369
rect 16853 21335 16911 21341
rect 16853 21332 16865 21335
rect 16816 21304 16865 21332
rect 16816 21292 16822 21304
rect 16853 21301 16865 21304
rect 16899 21301 16911 21335
rect 16853 21295 16911 21301
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 18141 21335 18199 21341
rect 18141 21332 18153 21335
rect 17552 21304 18153 21332
rect 17552 21292 17558 21304
rect 18141 21301 18153 21304
rect 18187 21332 18199 21335
rect 18598 21332 18604 21344
rect 18187 21304 18604 21332
rect 18187 21301 18199 21304
rect 18141 21295 18199 21301
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 18690 21292 18696 21344
rect 18748 21332 18754 21344
rect 18969 21335 19027 21341
rect 18969 21332 18981 21335
rect 18748 21304 18981 21332
rect 18748 21292 18754 21304
rect 18969 21301 18981 21304
rect 19015 21301 19027 21335
rect 18969 21295 19027 21301
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 20027 21335 20085 21341
rect 20027 21332 20039 21335
rect 19484 21304 20039 21332
rect 19484 21292 19490 21304
rect 20027 21301 20039 21304
rect 20073 21301 20085 21335
rect 20027 21295 20085 21301
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 1394 21088 1400 21140
rect 1452 21128 1458 21140
rect 2869 21131 2927 21137
rect 2869 21128 2881 21131
rect 1452 21100 2881 21128
rect 1452 21088 1458 21100
rect 2869 21097 2881 21100
rect 2915 21097 2927 21131
rect 2869 21091 2927 21097
rect 4246 21088 4252 21140
rect 4304 21128 4310 21140
rect 5074 21128 5080 21140
rect 4304 21100 5080 21128
rect 4304 21088 4310 21100
rect 2590 21060 2596 21072
rect 2551 21032 2596 21060
rect 2590 21020 2596 21032
rect 2648 21020 2654 21072
rect 3142 21020 3148 21072
rect 3200 21060 3206 21072
rect 4338 21060 4344 21072
rect 3200 21032 4344 21060
rect 3200 21020 3206 21032
rect 4338 21020 4344 21032
rect 4396 21020 4402 21072
rect 4525 21063 4583 21069
rect 4525 21029 4537 21063
rect 4571 21060 4583 21063
rect 4614 21060 4620 21072
rect 4571 21032 4620 21060
rect 4571 21029 4583 21032
rect 4525 21023 4583 21029
rect 4614 21020 4620 21032
rect 4672 21020 4678 21072
rect 1762 20992 1768 21004
rect 1723 20964 1768 20992
rect 1762 20952 1768 20964
rect 1820 20952 1826 21004
rect 2041 20995 2099 21001
rect 2041 20961 2053 20995
rect 2087 20992 2099 20995
rect 2774 20992 2780 21004
rect 2087 20964 2780 20992
rect 2087 20961 2099 20964
rect 2041 20955 2099 20961
rect 2774 20952 2780 20964
rect 2832 20952 2838 21004
rect 3329 20995 3387 21001
rect 3329 20961 3341 20995
rect 3375 20992 3387 20995
rect 3418 20992 3424 21004
rect 3375 20964 3424 20992
rect 3375 20961 3387 20964
rect 3329 20955 3387 20961
rect 3418 20952 3424 20964
rect 3476 20992 3482 21004
rect 3476 20964 4108 20992
rect 3476 20952 3482 20964
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20924 2283 20927
rect 3510 20924 3516 20936
rect 2271 20896 3516 20924
rect 2271 20893 2283 20896
rect 2225 20887 2283 20893
rect 3510 20884 3516 20896
rect 3568 20884 3574 20936
rect 2406 20816 2412 20868
rect 2464 20856 2470 20868
rect 3789 20859 3847 20865
rect 3789 20856 3801 20859
rect 2464 20828 3801 20856
rect 2464 20816 2470 20828
rect 3789 20825 3801 20828
rect 3835 20856 3847 20859
rect 3970 20856 3976 20868
rect 3835 20828 3976 20856
rect 3835 20825 3847 20828
rect 3789 20819 3847 20825
rect 3970 20816 3976 20828
rect 4028 20816 4034 20868
rect 4080 20856 4108 20964
rect 4430 20924 4436 20936
rect 4391 20896 4436 20924
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 4724 20924 4752 21100
rect 5074 21088 5080 21100
rect 5132 21088 5138 21140
rect 5902 21128 5908 21140
rect 5863 21100 5908 21128
rect 5902 21088 5908 21100
rect 5960 21088 5966 21140
rect 7101 21131 7159 21137
rect 7101 21097 7113 21131
rect 7147 21128 7159 21131
rect 7834 21128 7840 21140
rect 7147 21100 7840 21128
rect 7147 21097 7159 21100
rect 7101 21091 7159 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 8754 21088 8760 21140
rect 8812 21128 8818 21140
rect 12253 21131 12311 21137
rect 12253 21128 12265 21131
rect 8812 21100 12265 21128
rect 8812 21088 8818 21100
rect 12253 21097 12265 21100
rect 12299 21097 12311 21131
rect 13998 21128 14004 21140
rect 13959 21100 14004 21128
rect 12253 21091 12311 21097
rect 5629 21063 5687 21069
rect 5629 21029 5641 21063
rect 5675 21060 5687 21063
rect 5810 21060 5816 21072
rect 5675 21032 5816 21060
rect 5675 21029 5687 21032
rect 5629 21023 5687 21029
rect 5810 21020 5816 21032
rect 5868 21020 5874 21072
rect 7190 21020 7196 21072
rect 7248 21060 7254 21072
rect 9582 21060 9588 21072
rect 7248 21032 9588 21060
rect 7248 21020 7254 21032
rect 9582 21020 9588 21032
rect 9640 21060 9646 21072
rect 11882 21060 11888 21072
rect 9640 21032 11888 21060
rect 9640 21020 9646 21032
rect 5261 20995 5319 21001
rect 5261 20961 5273 20995
rect 5307 20992 5319 20995
rect 6178 20992 6184 21004
rect 5307 20964 6184 20992
rect 5307 20961 5319 20964
rect 5261 20955 5319 20961
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6362 20992 6368 21004
rect 6323 20964 6368 20992
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 6549 20995 6607 21001
rect 6549 20961 6561 20995
rect 6595 20992 6607 20995
rect 7466 20992 7472 21004
rect 6595 20964 7472 20992
rect 6595 20961 6607 20964
rect 6549 20955 6607 20961
rect 4893 20927 4951 20933
rect 4893 20924 4905 20927
rect 4724 20896 4905 20924
rect 4893 20893 4905 20896
rect 4939 20924 4951 20927
rect 5718 20924 5724 20936
rect 4939 20896 5724 20924
rect 4939 20893 4951 20896
rect 4893 20887 4951 20893
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 5902 20884 5908 20936
rect 5960 20924 5966 20936
rect 6564 20924 6592 20955
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 7926 20992 7932 21004
rect 7887 20964 7932 20992
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 8205 20995 8263 21001
rect 8205 20961 8217 20995
rect 8251 20992 8263 20995
rect 8573 20995 8631 21001
rect 8251 20964 8524 20992
rect 8251 20961 8263 20964
rect 8205 20955 8263 20961
rect 6730 20924 6736 20936
rect 5960 20896 6592 20924
rect 6691 20896 6736 20924
rect 5960 20884 5966 20896
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 7558 20884 7564 20936
rect 7616 20924 7622 20936
rect 8220 20924 8248 20955
rect 7616 20896 8248 20924
rect 8297 20927 8355 20933
rect 7616 20884 7622 20896
rect 8297 20893 8309 20927
rect 8343 20893 8355 20927
rect 8496 20924 8524 20964
rect 8573 20961 8585 20995
rect 8619 20992 8631 20995
rect 9214 20992 9220 21004
rect 8619 20964 9220 20992
rect 8619 20961 8631 20964
rect 8573 20955 8631 20961
rect 9214 20952 9220 20964
rect 9272 20952 9278 21004
rect 9692 21001 9720 21032
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20961 9735 20995
rect 9950 20992 9956 21004
rect 9911 20964 9956 20992
rect 9677 20955 9735 20961
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 11256 21001 11284 21032
rect 11882 21020 11888 21032
rect 11940 21020 11946 21072
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 11480 20964 11529 20992
rect 11480 20952 11486 20964
rect 11517 20961 11529 20964
rect 11563 20961 11575 20995
rect 11517 20955 11575 20961
rect 10137 20927 10195 20933
rect 10137 20924 10149 20927
rect 8496 20896 10149 20924
rect 8297 20887 8355 20893
rect 4338 20856 4344 20868
rect 4080 20828 4344 20856
rect 4338 20816 4344 20828
rect 4396 20816 4402 20868
rect 4706 20816 4712 20868
rect 4764 20856 4770 20868
rect 5350 20856 5356 20868
rect 4764 20828 5356 20856
rect 4764 20816 4770 20828
rect 5350 20816 5356 20828
rect 5408 20816 5414 20868
rect 5626 20816 5632 20868
rect 5684 20856 5690 20868
rect 7469 20859 7527 20865
rect 7469 20856 7481 20859
rect 5684 20828 7481 20856
rect 5684 20816 5690 20828
rect 7469 20825 7481 20828
rect 7515 20825 7527 20859
rect 7469 20819 7527 20825
rect 7650 20816 7656 20868
rect 7708 20856 7714 20868
rect 8312 20856 8340 20887
rect 9692 20868 9720 20896
rect 10137 20893 10149 20896
rect 10183 20893 10195 20927
rect 11330 20924 11336 20936
rect 10137 20887 10195 20893
rect 10244 20896 11336 20924
rect 7708 20828 8340 20856
rect 7708 20816 7714 20828
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 9033 20859 9091 20865
rect 9033 20856 9045 20859
rect 8536 20828 9045 20856
rect 8536 20816 8542 20828
rect 9033 20825 9045 20828
rect 9079 20825 9091 20859
rect 9033 20819 9091 20825
rect 9674 20816 9680 20868
rect 9732 20816 9738 20868
rect 9769 20859 9827 20865
rect 9769 20825 9781 20859
rect 9815 20856 9827 20859
rect 10244 20856 10272 20896
rect 11330 20884 11336 20896
rect 11388 20924 11394 20936
rect 11974 20924 11980 20936
rect 11388 20896 11606 20924
rect 11935 20896 11980 20924
rect 11388 20884 11394 20896
rect 9815 20828 10272 20856
rect 11578 20856 11606 20896
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 12268 20924 12296 21091
rect 13998 21088 14004 21100
rect 14056 21128 14062 21140
rect 14550 21128 14556 21140
rect 14056 21100 14556 21128
rect 14056 21088 14062 21100
rect 14550 21088 14556 21100
rect 14608 21088 14614 21140
rect 15010 21128 15016 21140
rect 14971 21100 15016 21128
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 15562 21128 15568 21140
rect 15344 21100 15568 21128
rect 15344 21088 15350 21100
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 15028 21060 15056 21088
rect 15381 21063 15439 21069
rect 15381 21060 15393 21063
rect 15028 21032 15393 21060
rect 15381 21029 15393 21032
rect 15427 21029 15439 21063
rect 15381 21023 15439 21029
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 15528 21032 15573 21060
rect 15528 21020 15534 21032
rect 16758 21020 16764 21072
rect 16816 21060 16822 21072
rect 17037 21063 17095 21069
rect 17037 21060 17049 21063
rect 16816 21032 17049 21060
rect 16816 21020 16822 21032
rect 17037 21029 17049 21032
rect 17083 21029 17095 21063
rect 17037 21023 17095 21029
rect 18046 21020 18052 21072
rect 18104 21060 18110 21072
rect 18506 21060 18512 21072
rect 18104 21032 18512 21060
rect 18104 21020 18110 21032
rect 18506 21020 18512 21032
rect 18564 21020 18570 21072
rect 18601 21063 18659 21069
rect 18601 21029 18613 21063
rect 18647 21060 18659 21063
rect 18966 21060 18972 21072
rect 18647 21032 18972 21060
rect 18647 21029 18659 21032
rect 18601 21023 18659 21029
rect 18966 21020 18972 21032
rect 19024 21020 19030 21072
rect 20806 21020 20812 21072
rect 20864 21060 20870 21072
rect 20993 21063 21051 21069
rect 20993 21060 21005 21063
rect 20864 21032 21005 21060
rect 20864 21020 20870 21032
rect 20993 21029 21005 21032
rect 21039 21029 21051 21063
rect 20993 21023 21051 21029
rect 21085 21063 21143 21069
rect 21085 21029 21097 21063
rect 21131 21060 21143 21063
rect 21358 21060 21364 21072
rect 21131 21032 21364 21060
rect 21131 21029 21143 21032
rect 21085 21023 21143 21029
rect 21358 21020 21364 21032
rect 21416 21020 21422 21072
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12860 20964 12909 20992
rect 12860 20952 12866 20964
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 12986 20952 12992 21004
rect 13044 20992 13050 21004
rect 13541 20995 13599 21001
rect 13541 20992 13553 20995
rect 13044 20964 13553 20992
rect 13044 20952 13050 20964
rect 13541 20961 13553 20964
rect 13587 20992 13599 20995
rect 14826 20992 14832 21004
rect 13587 20964 14832 20992
rect 13587 20961 13599 20964
rect 13541 20955 13599 20961
rect 14826 20952 14832 20964
rect 14884 20952 14890 21004
rect 12268 20896 13814 20924
rect 12986 20856 12992 20868
rect 11578 20828 12992 20856
rect 9815 20825 9827 20828
rect 9769 20819 9827 20825
rect 4522 20748 4528 20800
rect 4580 20788 4586 20800
rect 4663 20791 4721 20797
rect 4663 20788 4675 20791
rect 4580 20760 4675 20788
rect 4580 20748 4586 20760
rect 4663 20757 4675 20760
rect 4709 20757 4721 20791
rect 4663 20751 4721 20757
rect 4801 20791 4859 20797
rect 4801 20757 4813 20791
rect 4847 20788 4859 20791
rect 5442 20788 5448 20800
rect 4847 20760 5448 20788
rect 4847 20757 4859 20760
rect 4801 20751 4859 20757
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 7190 20748 7196 20800
rect 7248 20788 7254 20800
rect 8665 20791 8723 20797
rect 8665 20788 8677 20791
rect 7248 20760 8677 20788
rect 7248 20748 7254 20760
rect 8665 20757 8677 20760
rect 8711 20757 8723 20791
rect 8665 20751 8723 20757
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 9401 20791 9459 20797
rect 9401 20788 9413 20791
rect 8996 20760 9413 20788
rect 8996 20748 9002 20760
rect 9401 20757 9413 20760
rect 9447 20788 9459 20791
rect 9784 20788 9812 20819
rect 12986 20816 12992 20828
rect 13044 20816 13050 20868
rect 13786 20856 13814 20896
rect 14918 20884 14924 20936
rect 14976 20924 14982 20936
rect 15746 20924 15752 20936
rect 14976 20896 15752 20924
rect 14976 20884 14982 20896
rect 15746 20884 15752 20896
rect 15804 20884 15810 20936
rect 16666 20884 16672 20936
rect 16724 20924 16730 20936
rect 16945 20927 17003 20933
rect 16945 20924 16957 20927
rect 16724 20896 16957 20924
rect 16724 20884 16730 20896
rect 16945 20893 16957 20896
rect 16991 20893 17003 20927
rect 16945 20887 17003 20893
rect 17589 20927 17647 20933
rect 17589 20893 17601 20927
rect 17635 20924 17647 20927
rect 19153 20927 19211 20933
rect 19153 20924 19165 20927
rect 17635 20896 19165 20924
rect 17635 20893 17647 20896
rect 17589 20887 17647 20893
rect 19153 20893 19165 20896
rect 19199 20924 19211 20927
rect 21266 20924 21272 20936
rect 19199 20896 21272 20924
rect 19199 20893 19211 20896
rect 19153 20887 19211 20893
rect 15933 20859 15991 20865
rect 15933 20856 15945 20859
rect 13786 20828 15945 20856
rect 15933 20825 15945 20828
rect 15979 20856 15991 20859
rect 17604 20856 17632 20887
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 21542 20856 21548 20868
rect 15979 20828 17632 20856
rect 21503 20828 21548 20856
rect 15979 20825 15991 20828
rect 15933 20819 15991 20825
rect 21542 20816 21548 20828
rect 21600 20816 21606 20868
rect 10686 20788 10692 20800
rect 9447 20760 9812 20788
rect 10647 20760 10692 20788
rect 9447 20757 9459 20760
rect 9401 20751 9459 20757
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 11149 20791 11207 20797
rect 11149 20757 11161 20791
rect 11195 20788 11207 20791
rect 11422 20788 11428 20800
rect 11195 20760 11428 20788
rect 11195 20757 11207 20760
rect 11149 20751 11207 20757
rect 11422 20748 11428 20760
rect 11480 20748 11486 20800
rect 12618 20788 12624 20800
rect 12579 20760 12624 20788
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 16114 20788 16120 20800
rect 14792 20760 16120 20788
rect 14792 20748 14798 20760
rect 16114 20748 16120 20760
rect 16172 20788 16178 20800
rect 17678 20788 17684 20800
rect 16172 20760 17684 20788
rect 16172 20748 16178 20760
rect 17678 20748 17684 20760
rect 17736 20788 17742 20800
rect 18690 20788 18696 20800
rect 17736 20760 18696 20788
rect 17736 20748 17742 20760
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3418 20584 3424 20596
rect 3099 20556 3424 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 4249 20587 4307 20593
rect 4249 20553 4261 20587
rect 4295 20584 4307 20587
rect 4614 20584 4620 20596
rect 4295 20556 4620 20584
rect 4295 20553 4307 20556
rect 4249 20547 4307 20553
rect 4614 20544 4620 20556
rect 4672 20584 4678 20596
rect 5442 20584 5448 20596
rect 4672 20556 5448 20584
rect 4672 20544 4678 20556
rect 5442 20544 5448 20556
rect 5500 20544 5506 20596
rect 5718 20584 5724 20596
rect 5679 20556 5724 20584
rect 5718 20544 5724 20556
rect 5776 20584 5782 20596
rect 6089 20587 6147 20593
rect 6089 20584 6101 20587
rect 5776 20556 6101 20584
rect 5776 20544 5782 20556
rect 6089 20553 6101 20556
rect 6135 20553 6147 20587
rect 6089 20547 6147 20553
rect 7282 20544 7288 20596
rect 7340 20584 7346 20596
rect 9217 20587 9275 20593
rect 9217 20584 9229 20587
rect 7340 20556 9229 20584
rect 7340 20544 7346 20556
rect 9217 20553 9229 20556
rect 9263 20584 9275 20587
rect 9950 20584 9956 20596
rect 9263 20556 9956 20584
rect 9263 20553 9275 20556
rect 9217 20547 9275 20553
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 11425 20587 11483 20593
rect 11425 20553 11437 20587
rect 11471 20584 11483 20587
rect 13722 20584 13728 20596
rect 11471 20556 13728 20584
rect 11471 20553 11483 20556
rect 11425 20547 11483 20553
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 18564 20556 19441 20584
rect 18564 20544 18570 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 20806 20584 20812 20596
rect 20767 20556 20812 20584
rect 19429 20547 19487 20553
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 21450 20584 21456 20596
rect 21411 20556 21456 20584
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 3326 20516 3332 20528
rect 3160 20488 3332 20516
rect 3160 20457 3188 20488
rect 3326 20476 3332 20488
rect 3384 20516 3390 20528
rect 3384 20488 3648 20516
rect 3384 20476 3390 20488
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20448 2743 20451
rect 3145 20451 3203 20457
rect 3145 20448 3157 20451
rect 2731 20420 3157 20448
rect 2731 20417 2743 20420
rect 2685 20411 2743 20417
rect 3145 20417 3157 20420
rect 3191 20417 3203 20451
rect 3620 20448 3648 20488
rect 4154 20476 4160 20528
rect 4212 20516 4218 20528
rect 4479 20519 4537 20525
rect 4479 20516 4491 20519
rect 4212 20488 4491 20516
rect 4212 20476 4218 20488
rect 4479 20485 4491 20488
rect 4525 20485 4537 20519
rect 4479 20479 4537 20485
rect 5902 20476 5908 20528
rect 5960 20516 5966 20528
rect 6822 20516 6828 20528
rect 5960 20488 6828 20516
rect 5960 20476 5966 20488
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 8481 20519 8539 20525
rect 8481 20516 8493 20519
rect 8352 20488 8493 20516
rect 8352 20476 8358 20488
rect 8481 20485 8493 20488
rect 8527 20485 8539 20519
rect 9582 20516 9588 20528
rect 8481 20479 8539 20485
rect 8588 20488 8892 20516
rect 9543 20488 9588 20516
rect 3881 20451 3939 20457
rect 3881 20448 3893 20451
rect 3620 20420 3893 20448
rect 3145 20411 3203 20417
rect 3881 20417 3893 20420
rect 3927 20448 3939 20451
rect 4614 20448 4620 20460
rect 3927 20420 4620 20448
rect 3927 20417 3939 20420
rect 3881 20411 3939 20417
rect 4614 20408 4620 20420
rect 4672 20448 4678 20460
rect 4709 20451 4767 20457
rect 4709 20448 4721 20451
rect 4672 20420 4721 20448
rect 4672 20408 4678 20420
rect 4709 20417 4721 20420
rect 4755 20417 4767 20451
rect 4709 20411 4767 20417
rect 4890 20408 4896 20460
rect 4948 20448 4954 20460
rect 8588 20448 8616 20488
rect 4948 20420 8616 20448
rect 8864 20448 8892 20488
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 9674 20476 9680 20528
rect 9732 20516 9738 20528
rect 10689 20519 10747 20525
rect 10689 20516 10701 20519
rect 9732 20488 10701 20516
rect 9732 20476 9738 20488
rect 9743 20448 9771 20488
rect 10689 20485 10701 20488
rect 10735 20485 10747 20519
rect 10689 20479 10747 20485
rect 11054 20476 11060 20528
rect 11112 20516 11118 20528
rect 12342 20516 12348 20528
rect 11112 20488 12348 20516
rect 11112 20476 11118 20488
rect 12342 20476 12348 20488
rect 12400 20476 12406 20528
rect 16850 20516 16856 20528
rect 14384 20488 16856 20516
rect 13909 20451 13967 20457
rect 8864 20420 13768 20448
rect 4948 20408 4954 20420
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 2924 20383 2982 20389
rect 1443 20352 2084 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 106 20204 112 20256
rect 164 20244 170 20256
rect 2056 20253 2084 20352
rect 2924 20349 2936 20383
rect 2970 20380 2982 20383
rect 3418 20380 3424 20392
rect 2970 20352 3424 20380
rect 2970 20349 2982 20352
rect 2924 20343 2982 20349
rect 3418 20340 3424 20352
rect 3476 20340 3482 20392
rect 3602 20340 3608 20392
rect 3660 20380 3666 20392
rect 6822 20380 6828 20392
rect 3660 20352 6828 20380
rect 3660 20340 3666 20352
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20349 7251 20383
rect 7193 20343 7251 20349
rect 7469 20383 7527 20389
rect 7469 20349 7481 20383
rect 7515 20380 7527 20383
rect 7834 20380 7840 20392
rect 7515 20352 7840 20380
rect 7515 20349 7527 20352
rect 7469 20343 7527 20349
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20312 2835 20315
rect 4154 20312 4160 20324
rect 2823 20284 4160 20312
rect 2823 20281 2835 20284
rect 2777 20275 2835 20281
rect 4154 20272 4160 20284
rect 4212 20312 4218 20324
rect 4341 20315 4399 20321
rect 4341 20312 4353 20315
rect 4212 20284 4353 20312
rect 4212 20272 4218 20284
rect 4341 20281 4353 20284
rect 4387 20312 4399 20315
rect 4982 20312 4988 20324
rect 4387 20284 4988 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 4982 20272 4988 20284
rect 5040 20272 5046 20324
rect 5077 20315 5135 20321
rect 5077 20281 5089 20315
rect 5123 20312 5135 20315
rect 5718 20312 5724 20324
rect 5123 20284 5724 20312
rect 5123 20281 5135 20284
rect 5077 20275 5135 20281
rect 5718 20272 5724 20284
rect 5776 20272 5782 20324
rect 6362 20272 6368 20324
rect 6420 20312 6426 20324
rect 6549 20315 6607 20321
rect 6549 20312 6561 20315
rect 6420 20284 6561 20312
rect 6420 20272 6426 20284
rect 6549 20281 6561 20284
rect 6595 20312 6607 20315
rect 7208 20312 7236 20343
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 8700 20383 8758 20389
rect 8700 20380 8712 20383
rect 8352 20352 8712 20380
rect 8352 20340 8358 20352
rect 8700 20349 8712 20352
rect 8746 20349 8758 20383
rect 8700 20343 8758 20349
rect 9030 20340 9036 20392
rect 9088 20380 9094 20392
rect 9677 20383 9735 20389
rect 9088 20352 9674 20380
rect 9088 20340 9094 20352
rect 7282 20312 7288 20324
rect 6595 20284 7288 20312
rect 6595 20281 6607 20284
rect 6549 20275 6607 20281
rect 7282 20272 7288 20284
rect 7340 20312 7346 20324
rect 7926 20312 7932 20324
rect 7340 20284 7932 20312
rect 7340 20272 7346 20284
rect 7926 20272 7932 20284
rect 7984 20312 7990 20324
rect 8021 20315 8079 20321
rect 8021 20312 8033 20315
rect 7984 20284 8033 20312
rect 7984 20272 7990 20284
rect 8021 20281 8033 20284
rect 8067 20312 8079 20315
rect 8803 20315 8861 20321
rect 8067 20284 8616 20312
rect 8067 20281 8079 20284
rect 8021 20275 8079 20281
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 164 20216 1593 20244
rect 164 20204 170 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 1581 20207 1639 20213
rect 2041 20247 2099 20253
rect 2041 20213 2053 20247
rect 2087 20244 2099 20247
rect 2682 20244 2688 20256
rect 2087 20216 2688 20244
rect 2087 20213 2099 20216
rect 2041 20207 2099 20213
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 3421 20247 3479 20253
rect 3421 20213 3433 20247
rect 3467 20244 3479 20247
rect 3694 20244 3700 20256
rect 3467 20216 3700 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 3694 20204 3700 20216
rect 3752 20204 3758 20256
rect 3878 20204 3884 20256
rect 3936 20244 3942 20256
rect 4890 20244 4896 20256
rect 3936 20216 4896 20244
rect 3936 20204 3942 20216
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7009 20247 7067 20253
rect 7009 20244 7021 20247
rect 6972 20216 7021 20244
rect 6972 20204 6978 20216
rect 7009 20213 7021 20216
rect 7055 20213 7067 20247
rect 8588 20244 8616 20284
rect 8803 20281 8815 20315
rect 8849 20312 8861 20315
rect 9646 20312 9674 20352
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 9743 20380 9771 20420
rect 9723 20352 9771 20380
rect 10229 20383 10287 20389
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 10229 20349 10241 20383
rect 10275 20349 10287 20383
rect 10229 20343 10287 20349
rect 9766 20312 9772 20324
rect 8849 20284 9772 20312
rect 8849 20281 8861 20284
rect 8803 20275 8861 20281
rect 9766 20272 9772 20284
rect 9824 20312 9830 20324
rect 10244 20312 10272 20343
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 11241 20383 11299 20389
rect 11241 20380 11253 20383
rect 10836 20352 11253 20380
rect 10836 20340 10842 20352
rect 11241 20349 11253 20352
rect 11287 20349 11299 20383
rect 11882 20380 11888 20392
rect 11843 20352 11888 20380
rect 11241 20343 11299 20349
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12434 20380 12440 20392
rect 12299 20352 12440 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 12710 20340 12716 20392
rect 12768 20380 12774 20392
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12768 20352 12909 20380
rect 12768 20340 12774 20352
rect 12897 20349 12909 20352
rect 12943 20349 12955 20383
rect 13740 20380 13768 20420
rect 13909 20417 13921 20451
rect 13955 20448 13967 20451
rect 13998 20448 14004 20460
rect 13955 20420 14004 20448
rect 13955 20417 13967 20420
rect 13909 20411 13967 20417
rect 13998 20408 14004 20420
rect 14056 20448 14062 20460
rect 14384 20448 14412 20488
rect 16850 20476 16856 20488
rect 16908 20476 16914 20528
rect 16942 20476 16948 20528
rect 17000 20516 17006 20528
rect 20070 20516 20076 20528
rect 17000 20488 20076 20516
rect 17000 20476 17006 20488
rect 20070 20476 20076 20488
rect 20128 20476 20134 20528
rect 20165 20519 20223 20525
rect 20165 20485 20177 20519
rect 20211 20516 20223 20519
rect 22646 20516 22652 20528
rect 20211 20488 22652 20516
rect 20211 20485 20223 20488
rect 20165 20479 20223 20485
rect 18874 20448 18880 20460
rect 14056 20420 14412 20448
rect 14056 20408 14062 20420
rect 14277 20383 14335 20389
rect 13740 20352 13952 20380
rect 12897 20343 12955 20349
rect 10410 20312 10416 20324
rect 9824 20284 10272 20312
rect 10371 20284 10416 20312
rect 9824 20272 9830 20284
rect 10042 20244 10048 20256
rect 8588 20216 10048 20244
rect 7009 20207 7067 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 10244 20244 10272 20284
rect 10410 20272 10416 20284
rect 10468 20272 10474 20324
rect 11698 20272 11704 20324
rect 11756 20312 11762 20324
rect 13924 20312 13952 20352
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 14384 20380 14412 20420
rect 15856 20420 18880 20448
rect 14550 20380 14556 20392
rect 14323 20352 14412 20380
rect 14511 20352 14556 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 14792 20352 15025 20380
rect 14792 20340 14798 20352
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15856 20389 15884 20420
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 15252 20352 15485 20380
rect 15252 20340 15258 20352
rect 15473 20349 15485 20352
rect 15519 20380 15531 20383
rect 15841 20383 15899 20389
rect 15841 20380 15853 20383
rect 15519 20352 15853 20380
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 15841 20349 15853 20352
rect 15887 20349 15899 20383
rect 16114 20380 16120 20392
rect 16075 20352 16120 20380
rect 15841 20343 15899 20349
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20349 18383 20383
rect 18325 20343 18383 20349
rect 15378 20312 15384 20324
rect 11756 20284 12480 20312
rect 13924 20284 15384 20312
rect 11756 20272 11762 20284
rect 11146 20244 11152 20256
rect 10244 20216 11152 20244
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 12452 20244 12480 20284
rect 15378 20272 15384 20284
rect 15436 20272 15442 20324
rect 16758 20272 16764 20324
rect 16816 20312 16822 20324
rect 16853 20315 16911 20321
rect 16853 20312 16865 20315
rect 16816 20284 16865 20312
rect 16816 20272 16822 20284
rect 16853 20281 16865 20284
rect 16899 20281 16911 20315
rect 16853 20275 16911 20281
rect 17865 20315 17923 20321
rect 17865 20281 17877 20315
rect 17911 20312 17923 20315
rect 18340 20312 18368 20343
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18472 20352 18521 20380
rect 18472 20340 18478 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 19680 20383 19738 20389
rect 19680 20349 19692 20383
rect 19726 20380 19738 20383
rect 20180 20380 20208 20479
rect 22646 20476 22652 20488
rect 22704 20476 22710 20528
rect 19726 20352 20208 20380
rect 20968 20383 21026 20389
rect 19726 20349 19738 20352
rect 19680 20343 19738 20349
rect 20968 20349 20980 20383
rect 21014 20380 21026 20383
rect 21450 20380 21456 20392
rect 21014 20352 21456 20380
rect 21014 20349 21026 20352
rect 20968 20343 21026 20349
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 19518 20312 19524 20324
rect 17911 20284 19524 20312
rect 17911 20281 17923 20284
rect 17865 20275 17923 20281
rect 19518 20272 19524 20284
rect 19576 20272 19582 20324
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 21358 20312 21364 20324
rect 20588 20284 21364 20312
rect 20588 20272 20594 20284
rect 21358 20272 21364 20284
rect 21416 20312 21422 20324
rect 21729 20315 21787 20321
rect 21729 20312 21741 20315
rect 21416 20284 21741 20312
rect 21416 20272 21422 20284
rect 21729 20281 21741 20284
rect 21775 20281 21787 20315
rect 21729 20275 21787 20281
rect 12529 20247 12587 20253
rect 12529 20244 12541 20247
rect 12452 20216 12541 20244
rect 12529 20213 12541 20216
rect 12575 20213 12587 20247
rect 12529 20207 12587 20213
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 13449 20247 13507 20253
rect 13449 20244 13461 20247
rect 12860 20216 13461 20244
rect 12860 20204 12866 20216
rect 13449 20213 13461 20216
rect 13495 20244 13507 20247
rect 13538 20244 13544 20256
rect 13495 20216 13544 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 14093 20247 14151 20253
rect 14093 20213 14105 20247
rect 14139 20244 14151 20247
rect 14182 20244 14188 20256
rect 14139 20216 14188 20244
rect 14139 20213 14151 20216
rect 14093 20207 14151 20213
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 15654 20244 15660 20256
rect 15615 20216 15660 20244
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 16666 20204 16672 20256
rect 16724 20244 16730 20256
rect 17221 20247 17279 20253
rect 17221 20244 17233 20247
rect 16724 20216 17233 20244
rect 16724 20204 16730 20216
rect 17221 20213 17233 20216
rect 17267 20213 17279 20247
rect 18138 20244 18144 20256
rect 18099 20216 18144 20244
rect 17221 20207 17279 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 19024 20216 19073 20244
rect 19024 20204 19030 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19751 20247 19809 20253
rect 19751 20244 19763 20247
rect 19668 20216 19763 20244
rect 19668 20204 19674 20216
rect 19751 20213 19763 20216
rect 19797 20213 19809 20247
rect 19751 20207 19809 20213
rect 19886 20204 19892 20256
rect 19944 20244 19950 20256
rect 21039 20247 21097 20253
rect 21039 20244 21051 20247
rect 19944 20216 21051 20244
rect 19944 20204 19950 20216
rect 21039 20213 21051 20216
rect 21085 20213 21097 20247
rect 21039 20207 21097 20213
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 1535 20043 1593 20049
rect 1535 20009 1547 20043
rect 1581 20040 1593 20043
rect 1670 20040 1676 20052
rect 1581 20012 1676 20040
rect 1581 20009 1593 20012
rect 1535 20003 1593 20009
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 1762 20000 1768 20052
rect 1820 20040 1826 20052
rect 1857 20043 1915 20049
rect 1857 20040 1869 20043
rect 1820 20012 1869 20040
rect 1820 20000 1826 20012
rect 1857 20009 1869 20012
rect 1903 20040 1915 20043
rect 3786 20040 3792 20052
rect 1903 20012 3792 20040
rect 1903 20009 1915 20012
rect 1857 20003 1915 20009
rect 3786 20000 3792 20012
rect 3844 20040 3850 20052
rect 3844 20012 4844 20040
rect 3844 20000 3850 20012
rect 3694 19972 3700 19984
rect 2424 19944 3700 19972
rect 1464 19907 1522 19913
rect 1464 19873 1476 19907
rect 1510 19904 1522 19907
rect 2314 19904 2320 19916
rect 1510 19876 2320 19904
rect 1510 19873 1522 19876
rect 1464 19867 1522 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2424 19913 2452 19944
rect 3694 19932 3700 19944
rect 3752 19932 3758 19984
rect 3881 19975 3939 19981
rect 3881 19941 3893 19975
rect 3927 19972 3939 19975
rect 3970 19972 3976 19984
rect 3927 19944 3976 19972
rect 3927 19941 3939 19944
rect 3881 19935 3939 19941
rect 3970 19932 3976 19944
rect 4028 19932 4034 19984
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 4212 19944 4292 19972
rect 4212 19932 4218 19944
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 2590 19864 2596 19916
rect 2648 19904 2654 19916
rect 2685 19907 2743 19913
rect 2685 19904 2697 19907
rect 2648 19876 2697 19904
rect 2648 19864 2654 19876
rect 2685 19873 2697 19876
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 3050 19836 3056 19848
rect 1820 19808 3056 19836
rect 1820 19796 1826 19808
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3970 19836 3976 19848
rect 3191 19808 3976 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3970 19796 3976 19808
rect 4028 19836 4034 19848
rect 4264 19845 4292 19944
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 4028 19808 4261 19836
rect 4028 19796 4034 19808
rect 4249 19805 4261 19808
rect 4295 19836 4307 19839
rect 4448 19836 4476 19867
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 4663 19907 4721 19913
rect 4663 19904 4675 19907
rect 4580 19876 4675 19904
rect 4580 19864 4586 19876
rect 4663 19873 4675 19876
rect 4709 19873 4721 19907
rect 4816 19904 4844 20012
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5445 20043 5503 20049
rect 5445 20040 5457 20043
rect 5040 20012 5457 20040
rect 5040 20000 5046 20012
rect 5445 20009 5457 20012
rect 5491 20040 5503 20043
rect 5534 20040 5540 20052
rect 5491 20012 5540 20040
rect 5491 20009 5503 20012
rect 5445 20003 5503 20009
rect 5534 20000 5540 20012
rect 5592 20040 5598 20052
rect 5902 20040 5908 20052
rect 5592 20012 5810 20040
rect 5863 20012 5908 20040
rect 5592 20000 5598 20012
rect 5782 19984 5810 20012
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 6086 20040 6092 20052
rect 6047 20012 6092 20040
rect 6086 20000 6092 20012
rect 6144 20000 6150 20052
rect 6454 20000 6460 20052
rect 6512 20000 6518 20052
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 15378 20040 15384 20052
rect 6880 20012 13814 20040
rect 15339 20012 15384 20040
rect 6880 20000 6886 20012
rect 5782 19944 5816 19984
rect 5810 19932 5816 19944
rect 5868 19932 5874 19984
rect 6472 19972 6500 20000
rect 6012 19944 6500 19972
rect 7101 19975 7159 19981
rect 6012 19913 6040 19944
rect 7101 19941 7113 19975
rect 7147 19972 7159 19975
rect 7282 19972 7288 19984
rect 7147 19944 7288 19972
rect 7147 19941 7159 19944
rect 7101 19935 7159 19941
rect 7282 19932 7288 19944
rect 7340 19932 7346 19984
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 7653 19975 7711 19981
rect 7653 19972 7665 19975
rect 7616 19944 7665 19972
rect 7616 19932 7622 19944
rect 7653 19941 7665 19944
rect 7699 19941 7711 19975
rect 7653 19935 7711 19941
rect 7742 19932 7748 19984
rect 7800 19972 7806 19984
rect 10413 19975 10471 19981
rect 10413 19972 10425 19975
rect 7800 19944 10425 19972
rect 7800 19932 7806 19944
rect 10413 19941 10425 19944
rect 10459 19941 10471 19975
rect 10413 19935 10471 19941
rect 11146 19932 11152 19984
rect 11204 19972 11210 19984
rect 12066 19972 12072 19984
rect 11204 19944 12072 19972
rect 11204 19932 11210 19944
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 4816 19876 6009 19904
rect 4663 19867 4721 19873
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 5997 19867 6055 19873
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 6457 19907 6515 19913
rect 6457 19904 6469 19907
rect 6420 19876 6469 19904
rect 6420 19864 6426 19876
rect 6457 19873 6469 19876
rect 6503 19873 6515 19907
rect 8294 19904 8300 19916
rect 8255 19876 8300 19904
rect 6457 19867 6515 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 8481 19907 8539 19913
rect 8481 19904 8493 19907
rect 8444 19876 8493 19904
rect 8444 19864 8450 19876
rect 8481 19873 8493 19876
rect 8527 19873 8539 19907
rect 8481 19867 8539 19873
rect 8938 19864 8944 19916
rect 8996 19904 9002 19916
rect 8996 19876 9041 19904
rect 8996 19864 9002 19876
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9640 19876 9689 19904
rect 9640 19864 9646 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9916 19876 10149 19904
rect 9916 19864 9922 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11716 19913 11744 19944
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 12250 19932 12256 19984
rect 12308 19972 12314 19984
rect 13786 19972 13814 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16945 20043 17003 20049
rect 16945 20040 16957 20043
rect 16172 20012 16957 20040
rect 16172 20000 16178 20012
rect 16945 20009 16957 20012
rect 16991 20009 17003 20043
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 16945 20003 17003 20009
rect 17052 20012 18521 20040
rect 15654 19972 15660 19984
rect 12308 19944 13124 19972
rect 13786 19944 15660 19972
rect 12308 19932 12314 19944
rect 11241 19907 11299 19913
rect 11241 19904 11253 19907
rect 11112 19876 11253 19904
rect 11112 19864 11118 19876
rect 11241 19873 11253 19876
rect 11287 19873 11299 19907
rect 11241 19867 11299 19873
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19873 11759 19907
rect 12802 19904 12808 19916
rect 11701 19867 11759 19873
rect 11808 19876 12808 19904
rect 4798 19836 4804 19848
rect 4295 19808 4476 19836
rect 4759 19808 4804 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19836 5227 19839
rect 7650 19836 7656 19848
rect 5215 19808 7656 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 7650 19796 7656 19808
rect 7708 19796 7714 19848
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 11808 19836 11836 19876
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 13096 19913 13124 19944
rect 15654 19932 15660 19944
rect 15712 19932 15718 19984
rect 16574 19932 16580 19984
rect 16632 19972 16638 19984
rect 17052 19972 17080 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21634 20040 21640 20052
rect 21131 20012 21640 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 16632 19944 17080 19972
rect 17420 19944 18920 19972
rect 16632 19932 16638 19944
rect 17420 19916 17448 19944
rect 13081 19907 13139 19913
rect 12952 19876 12997 19904
rect 12952 19864 12958 19876
rect 13081 19873 13093 19907
rect 13127 19904 13139 19907
rect 13354 19904 13360 19916
rect 13127 19876 13360 19904
rect 13127 19873 13139 19876
rect 13081 19867 13139 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 15010 19904 15016 19916
rect 13786 19876 15016 19904
rect 11974 19836 11980 19848
rect 8168 19808 11836 19836
rect 11935 19808 11980 19836
rect 8168 19796 8174 19808
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 12400 19808 13277 19836
rect 12400 19796 12406 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 13786 19836 13814 19876
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 15562 19904 15568 19916
rect 15523 19876 15568 19904
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15672 19876 15761 19904
rect 13504 19808 13814 19836
rect 13504 19796 13510 19808
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 14056 19808 14381 19836
rect 14056 19796 14062 19808
rect 14369 19805 14381 19808
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19836 15163 19839
rect 15470 19836 15476 19848
rect 15151 19808 15476 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 2498 19768 2504 19780
rect 2459 19740 2504 19768
rect 2498 19728 2504 19740
rect 2556 19728 2562 19780
rect 3602 19728 3608 19780
rect 3660 19768 3666 19780
rect 9490 19768 9496 19780
rect 3660 19740 9496 19768
rect 3660 19728 3666 19740
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 10042 19728 10048 19780
rect 10100 19768 10106 19780
rect 10100 19740 12572 19768
rect 10100 19728 10106 19740
rect 1210 19660 1216 19712
rect 1268 19700 1274 19712
rect 2222 19700 2228 19712
rect 1268 19672 2228 19700
rect 1268 19660 1274 19672
rect 2222 19660 2228 19672
rect 2280 19660 2286 19712
rect 2314 19660 2320 19712
rect 2372 19700 2378 19712
rect 2866 19700 2872 19712
rect 2372 19672 2872 19700
rect 2372 19660 2378 19672
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19700 3482 19712
rect 4246 19700 4252 19712
rect 3476 19672 4252 19700
rect 3476 19660 3482 19672
rect 4246 19660 4252 19672
rect 4304 19700 4310 19712
rect 4614 19709 4620 19712
rect 4571 19703 4620 19709
rect 4571 19700 4583 19703
rect 4304 19672 4583 19700
rect 4304 19660 4310 19672
rect 4571 19669 4583 19672
rect 4617 19669 4620 19703
rect 4571 19663 4620 19669
rect 4614 19660 4620 19663
rect 4672 19660 4678 19712
rect 5718 19660 5724 19712
rect 5776 19700 5782 19712
rect 6362 19700 6368 19712
rect 5776 19672 6368 19700
rect 5776 19660 5782 19672
rect 6362 19660 6368 19672
rect 6420 19700 6426 19712
rect 7282 19700 7288 19712
rect 6420 19672 7288 19700
rect 6420 19660 6426 19672
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 8754 19660 8760 19712
rect 8812 19700 8818 19712
rect 9033 19703 9091 19709
rect 9033 19700 9045 19703
rect 8812 19672 9045 19700
rect 8812 19660 8818 19672
rect 9033 19669 9045 19672
rect 9079 19669 9091 19703
rect 9033 19663 9091 19669
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19700 9459 19703
rect 9950 19700 9956 19712
rect 9447 19672 9956 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10778 19700 10784 19712
rect 10739 19672 10784 19700
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 11149 19703 11207 19709
rect 11149 19669 11161 19703
rect 11195 19700 11207 19703
rect 11422 19700 11428 19712
rect 11195 19672 11428 19700
rect 11195 19669 11207 19672
rect 11149 19663 11207 19669
rect 11422 19660 11428 19672
rect 11480 19700 11486 19712
rect 12250 19700 12256 19712
rect 11480 19672 12256 19700
rect 11480 19660 11486 19672
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12544 19709 12572 19740
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 14182 19768 14188 19780
rect 13688 19740 14188 19768
rect 13688 19728 13694 19740
rect 14182 19728 14188 19740
rect 14240 19728 14246 19780
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 15672 19768 15700 19876
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 16850 19904 16856 19916
rect 16811 19876 16856 19904
rect 15749 19867 15807 19873
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 17402 19904 17408 19916
rect 17363 19876 17408 19904
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 18598 19904 18604 19916
rect 18559 19876 18604 19904
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 18892 19913 18920 19944
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19904 18935 19907
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 18923 19876 19625 19904
rect 18923 19873 18935 19876
rect 18877 19867 18935 19873
rect 19613 19873 19625 19876
rect 19659 19904 19671 19907
rect 19978 19904 19984 19916
rect 19659 19876 19984 19904
rect 19659 19873 19671 19876
rect 19613 19867 19671 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 15838 19768 15844 19780
rect 14608 19740 15844 19768
rect 14608 19728 14614 19740
rect 15838 19728 15844 19740
rect 15896 19768 15902 19780
rect 18049 19771 18107 19777
rect 18049 19768 18061 19771
rect 15896 19740 18061 19768
rect 15896 19728 15902 19740
rect 18049 19737 18061 19740
rect 18095 19768 18107 19771
rect 18322 19768 18328 19780
rect 18095 19740 18328 19768
rect 18095 19737 18107 19740
rect 18049 19731 18107 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 12710 19700 12716 19712
rect 12575 19672 12716 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 14090 19700 14096 19712
rect 14003 19672 14096 19700
rect 14090 19660 14096 19672
rect 14148 19700 14154 19712
rect 16022 19700 16028 19712
rect 14148 19672 16028 19700
rect 14148 19660 14154 19672
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 21358 19700 21364 19712
rect 16724 19672 21364 19700
rect 16724 19660 16730 19672
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 2280 19468 2912 19496
rect 2280 19456 2286 19468
rect 2130 19388 2136 19440
rect 2188 19428 2194 19440
rect 2501 19431 2559 19437
rect 2188 19400 2452 19428
rect 2188 19388 2194 19400
rect 2424 19360 2452 19400
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2590 19428 2596 19440
rect 2547 19400 2596 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 2774 19428 2780 19440
rect 2735 19400 2780 19428
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 2884 19360 2912 19468
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 3878 19496 3884 19508
rect 3108 19468 3884 19496
rect 3108 19456 3114 19468
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 4798 19456 4804 19508
rect 4856 19496 4862 19508
rect 4985 19499 5043 19505
rect 4985 19496 4997 19499
rect 4856 19468 4997 19496
rect 4856 19456 4862 19468
rect 4985 19465 4997 19468
rect 5031 19496 5043 19499
rect 5031 19468 5304 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 5276 19440 5304 19468
rect 5442 19456 5448 19508
rect 5500 19496 5506 19508
rect 6362 19496 6368 19508
rect 5500 19468 6368 19496
rect 5500 19456 5506 19468
rect 6362 19456 6368 19468
rect 6420 19496 6426 19508
rect 6420 19468 7144 19496
rect 6420 19456 6426 19468
rect 4706 19428 4712 19440
rect 4264 19400 4712 19428
rect 4264 19360 4292 19400
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 5258 19388 5264 19440
rect 5316 19428 5322 19440
rect 5997 19431 6055 19437
rect 5997 19428 6009 19431
rect 5316 19400 6009 19428
rect 5316 19388 5322 19400
rect 5997 19397 6009 19400
rect 6043 19397 6055 19431
rect 5997 19391 6055 19397
rect 6273 19431 6331 19437
rect 6273 19397 6285 19431
rect 6319 19428 6331 19431
rect 6454 19428 6460 19440
rect 6319 19400 6460 19428
rect 6319 19397 6331 19400
rect 6273 19391 6331 19397
rect 6454 19388 6460 19400
rect 6512 19388 6518 19440
rect 7006 19428 7012 19440
rect 6967 19400 7012 19428
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 7116 19428 7144 19468
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 9217 19499 9275 19505
rect 9217 19496 9229 19499
rect 7524 19468 9229 19496
rect 7524 19456 7530 19468
rect 9217 19465 9229 19468
rect 9263 19496 9275 19499
rect 9309 19499 9367 19505
rect 9309 19496 9321 19499
rect 9263 19468 9321 19496
rect 9263 19465 9275 19468
rect 9217 19459 9275 19465
rect 9309 19465 9321 19468
rect 9355 19465 9367 19499
rect 9309 19459 9367 19465
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 10597 19499 10655 19505
rect 10597 19496 10609 19499
rect 9640 19468 10609 19496
rect 9640 19456 9646 19468
rect 10597 19465 10609 19468
rect 10643 19496 10655 19499
rect 11146 19496 11152 19508
rect 10643 19468 11152 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 11146 19456 11152 19468
rect 11204 19456 11210 19508
rect 11241 19499 11299 19505
rect 11241 19465 11253 19499
rect 11287 19496 11299 19499
rect 11606 19496 11612 19508
rect 11287 19468 11612 19496
rect 11287 19465 11299 19468
rect 11241 19459 11299 19465
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 13538 19496 13544 19508
rect 13499 19468 13544 19496
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 13633 19499 13691 19505
rect 13633 19465 13645 19499
rect 13679 19496 13691 19499
rect 13906 19496 13912 19508
rect 13679 19468 13912 19496
rect 13679 19465 13691 19468
rect 13633 19459 13691 19465
rect 13906 19456 13912 19468
rect 13964 19456 13970 19508
rect 14090 19456 14096 19508
rect 14148 19505 14154 19508
rect 14148 19499 14197 19505
rect 14148 19465 14151 19499
rect 14185 19465 14197 19499
rect 14148 19459 14197 19465
rect 14148 19456 14154 19459
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 16666 19496 16672 19508
rect 15436 19468 16672 19496
rect 15436 19456 15442 19468
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 16850 19496 16856 19508
rect 16811 19468 16856 19496
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 21315 19499 21373 19505
rect 21315 19496 21327 19499
rect 20680 19468 21327 19496
rect 20680 19456 20686 19468
rect 21315 19465 21327 19468
rect 21361 19465 21373 19499
rect 21315 19459 21373 19465
rect 7116 19400 8524 19428
rect 2424 19346 2820 19360
rect 2424 19332 2780 19346
rect 1210 19252 1216 19304
rect 1268 19292 1274 19304
rect 1397 19295 1455 19301
rect 1397 19292 1409 19295
rect 1268 19264 1409 19292
rect 1268 19252 1274 19264
rect 1397 19261 1409 19264
rect 1443 19261 1455 19295
rect 1397 19255 1455 19261
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19292 2007 19295
rect 2130 19292 2136 19304
rect 1995 19264 2136 19292
rect 1995 19261 2007 19264
rect 1949 19255 2007 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 2774 19294 2780 19332
rect 2832 19294 2838 19346
rect 2884 19332 4292 19360
rect 2996 19295 3054 19301
rect 2996 19261 3008 19295
rect 3042 19261 3054 19295
rect 3970 19292 3976 19304
rect 3931 19264 3976 19292
rect 2996 19255 3054 19261
rect 661 19227 719 19233
rect 661 19193 673 19227
rect 707 19224 719 19227
rect 3011 19224 3039 19255
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4264 19292 4292 19332
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 5353 19363 5411 19369
rect 5353 19360 5365 19363
rect 4672 19332 5365 19360
rect 4672 19320 4678 19332
rect 5353 19329 5365 19332
rect 5399 19360 5411 19363
rect 5810 19360 5816 19372
rect 5399 19332 5816 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 6178 19320 6184 19372
rect 6236 19360 6242 19372
rect 8496 19360 8524 19400
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 14277 19431 14335 19437
rect 14277 19428 14289 19431
rect 8628 19400 14044 19428
rect 8628 19388 8634 19400
rect 9030 19360 9036 19372
rect 6236 19332 8432 19360
rect 8496 19332 9036 19360
rect 6236 19320 6242 19332
rect 4430 19292 4436 19304
rect 4212 19264 4292 19292
rect 4391 19264 4436 19292
rect 4212 19252 4218 19264
rect 4430 19252 4436 19264
rect 4488 19252 4494 19304
rect 4522 19252 4528 19304
rect 4580 19292 4586 19304
rect 5537 19295 5595 19301
rect 5537 19292 5549 19295
rect 4580 19264 5549 19292
rect 4580 19252 4586 19264
rect 5537 19261 5549 19264
rect 5583 19292 5595 19295
rect 6089 19295 6147 19301
rect 6089 19292 6101 19295
rect 5583 19264 6101 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 6089 19261 6101 19264
rect 6135 19261 6147 19295
rect 6089 19255 6147 19261
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6696 19264 6837 19292
rect 6696 19252 6702 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7190 19292 7196 19304
rect 6972 19264 7196 19292
rect 6972 19252 6978 19264
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19292 7711 19295
rect 7926 19292 7932 19304
rect 7699 19264 7932 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8404 19301 8432 19332
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 11238 19360 11244 19372
rect 9508 19332 11244 19360
rect 9508 19301 9536 19332
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 13633 19363 13691 19369
rect 12124 19332 12940 19360
rect 12124 19320 12130 19332
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8367 19264 8401 19292
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 9217 19295 9275 19301
rect 8389 19255 8447 19261
rect 8496 19264 8978 19292
rect 3421 19227 3479 19233
rect 3421 19224 3433 19227
rect 707 19196 3433 19224
rect 707 19193 719 19196
rect 661 19187 719 19193
rect 3421 19193 3433 19196
rect 3467 19193 3479 19227
rect 3421 19187 3479 19193
rect 3694 19184 3700 19236
rect 3752 19224 3758 19236
rect 5902 19224 5908 19236
rect 3752 19196 5908 19224
rect 3752 19184 3758 19196
rect 5902 19184 5908 19196
rect 5960 19184 5966 19236
rect 5997 19227 6055 19233
rect 5997 19193 6009 19227
rect 6043 19224 6055 19227
rect 8404 19224 8432 19255
rect 8496 19224 8524 19264
rect 6043 19196 8524 19224
rect 8950 19224 8978 19264
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 9493 19295 9551 19301
rect 9493 19292 9505 19295
rect 9263 19264 9505 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 9493 19261 9505 19264
rect 9539 19261 9551 19295
rect 10042 19292 10048 19304
rect 10003 19264 10048 19292
rect 9493 19255 9551 19261
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 11057 19295 11115 19301
rect 11057 19261 11069 19295
rect 11103 19292 11115 19295
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11103 19264 11529 19292
rect 11103 19261 11115 19264
rect 11057 19255 11115 19261
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 11624 19264 12388 19292
rect 8950 19196 9674 19224
rect 6043 19193 6055 19196
rect 5997 19187 6055 19193
rect 753 19159 811 19165
rect 753 19125 765 19159
rect 799 19156 811 19159
rect 1489 19159 1547 19165
rect 1489 19156 1501 19159
rect 799 19128 1501 19156
rect 799 19125 811 19128
rect 753 19119 811 19125
rect 1489 19125 1501 19128
rect 1535 19125 1547 19159
rect 1489 19119 1547 19125
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 3099 19159 3157 19165
rect 3099 19156 3111 19159
rect 2924 19128 3111 19156
rect 2924 19116 2930 19128
rect 3099 19125 3111 19128
rect 3145 19125 3157 19159
rect 3878 19156 3884 19168
rect 3839 19128 3884 19156
rect 3099 19119 3157 19125
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4246 19156 4252 19168
rect 4207 19128 4252 19156
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 5718 19156 5724 19168
rect 5679 19128 5724 19156
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6319 19128 6561 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6549 19125 6561 19128
rect 6595 19156 6607 19159
rect 6638 19156 6644 19168
rect 6595 19128 6644 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 7377 19159 7435 19165
rect 7377 19156 7389 19159
rect 7248 19128 7389 19156
rect 7248 19116 7254 19128
rect 7377 19125 7389 19128
rect 7423 19156 7435 19159
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 7423 19128 7665 19156
rect 7423 19125 7435 19128
rect 7377 19119 7435 19125
rect 7653 19125 7665 19128
rect 7699 19156 7711 19159
rect 7745 19159 7803 19165
rect 7745 19156 7757 19159
rect 7699 19128 7757 19156
rect 7699 19125 7711 19128
rect 7653 19119 7711 19125
rect 7745 19125 7757 19128
rect 7791 19125 7803 19159
rect 8018 19156 8024 19168
rect 7979 19128 8024 19156
rect 7745 19119 7803 19125
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 8404 19156 8432 19196
rect 8757 19159 8815 19165
rect 8757 19156 8769 19159
rect 8352 19128 8769 19156
rect 8352 19116 8358 19128
rect 8757 19125 8769 19128
rect 8803 19125 8815 19159
rect 9646 19156 9674 19196
rect 10134 19184 10140 19236
rect 10192 19224 10198 19236
rect 10229 19227 10287 19233
rect 10229 19224 10241 19227
rect 10192 19196 10241 19224
rect 10192 19184 10198 19196
rect 10229 19193 10241 19196
rect 10275 19193 10287 19227
rect 11624 19224 11652 19264
rect 10229 19187 10287 19193
rect 10796 19196 11652 19224
rect 12360 19224 12388 19264
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 12912 19301 12940 19332
rect 13633 19329 13645 19363
rect 13679 19360 13691 19363
rect 13814 19360 13820 19372
rect 13679 19332 13820 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 13814 19320 13820 19332
rect 13872 19320 13878 19372
rect 14016 19334 14044 19400
rect 13924 19306 14044 19334
rect 14108 19400 14289 19428
rect 12897 19295 12955 19301
rect 12492 19264 12537 19292
rect 12492 19252 12498 19264
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 13078 19292 13084 19304
rect 12943 19264 13084 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 13725 19295 13783 19301
rect 13725 19261 13737 19295
rect 13771 19292 13783 19295
rect 13924 19292 13952 19306
rect 13771 19264 13952 19292
rect 14108 19292 14136 19400
rect 14277 19397 14289 19400
rect 14323 19397 14335 19431
rect 17770 19428 17776 19440
rect 14277 19391 14335 19397
rect 14384 19400 17776 19428
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14384 19369 14412 19400
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 18506 19388 18512 19440
rect 18564 19428 18570 19440
rect 18693 19431 18751 19437
rect 18693 19428 18705 19431
rect 18564 19400 18705 19428
rect 18564 19388 18570 19400
rect 18693 19397 18705 19400
rect 18739 19397 18751 19431
rect 18693 19391 18751 19397
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 14240 19332 14381 19360
rect 14240 19320 14246 19332
rect 14369 19329 14381 19332
rect 14415 19329 14427 19363
rect 14369 19323 14427 19329
rect 15488 19332 16436 19360
rect 15488 19292 15516 19332
rect 14108 19264 15516 19292
rect 15565 19295 15623 19301
rect 13771 19261 13783 19264
rect 13725 19255 13783 19261
rect 13170 19224 13176 19236
rect 12360 19196 13176 19224
rect 10796 19156 10824 19196
rect 13170 19184 13176 19196
rect 13228 19184 13234 19236
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 14000 19227 14058 19233
rect 14000 19224 14012 19227
rect 13964 19196 14012 19224
rect 13964 19184 13970 19196
rect 14000 19193 14012 19196
rect 14046 19193 14058 19227
rect 14000 19187 14058 19193
rect 9646 19128 10824 19156
rect 10965 19159 11023 19165
rect 8757 19119 8815 19125
rect 10965 19125 10977 19159
rect 11011 19156 11023 19159
rect 11054 19156 11060 19168
rect 11011 19128 11060 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 11517 19159 11575 19165
rect 11517 19125 11529 19159
rect 11563 19156 11575 19159
rect 11701 19159 11759 19165
rect 11701 19156 11713 19159
rect 11563 19128 11713 19156
rect 11563 19125 11575 19128
rect 11517 19119 11575 19125
rect 11701 19125 11713 19128
rect 11747 19156 11759 19159
rect 11882 19156 11888 19168
rect 11747 19128 11888 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 12529 19159 12587 19165
rect 12529 19156 12541 19159
rect 12308 19128 12541 19156
rect 12308 19116 12314 19128
rect 12529 19125 12541 19128
rect 12575 19125 12587 19159
rect 12529 19119 12587 19125
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13320 19128 13829 19156
rect 13320 19116 13326 19128
rect 13817 19125 13829 19128
rect 13863 19156 13875 19159
rect 14108 19156 14136 19264
rect 15565 19261 15577 19295
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 14458 19184 14464 19236
rect 14516 19224 14522 19236
rect 15381 19227 15439 19233
rect 15381 19224 15393 19227
rect 14516 19196 15393 19224
rect 14516 19184 14522 19196
rect 15381 19193 15393 19196
rect 15427 19224 15439 19227
rect 15580 19224 15608 19255
rect 15838 19252 15844 19304
rect 15896 19292 15902 19304
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 15896 19264 16037 19292
rect 15896 19252 15902 19264
rect 16025 19261 16037 19264
rect 16071 19261 16083 19295
rect 16408 19292 16436 19332
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 20165 19363 20223 19369
rect 20165 19360 20177 19363
rect 16540 19332 20177 19360
rect 16540 19320 16546 19332
rect 20165 19329 20177 19332
rect 20211 19329 20223 19363
rect 20165 19323 20223 19329
rect 17494 19292 17500 19304
rect 16408 19264 17500 19292
rect 16025 19255 16083 19261
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19536 19264 19625 19292
rect 15427 19196 15608 19224
rect 15427 19193 15439 19196
rect 15381 19187 15439 19193
rect 15746 19184 15752 19236
rect 15804 19224 15810 19236
rect 18138 19224 18144 19236
rect 15804 19196 18144 19224
rect 15804 19184 15810 19196
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 18288 19196 18333 19224
rect 18288 19184 18294 19196
rect 19536 19168 19564 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 19978 19252 19984 19304
rect 20036 19292 20042 19304
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 20036 19264 20085 19292
rect 20036 19252 20042 19264
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 20438 19252 20444 19304
rect 20496 19292 20502 19304
rect 21212 19295 21270 19301
rect 21212 19292 21224 19295
rect 20496 19264 21224 19292
rect 20496 19252 20502 19264
rect 21212 19261 21224 19264
rect 21258 19292 21270 19295
rect 21637 19295 21695 19301
rect 21637 19292 21649 19295
rect 21258 19264 21649 19292
rect 21258 19261 21270 19264
rect 21212 19255 21270 19261
rect 21637 19261 21649 19264
rect 21683 19292 21695 19295
rect 23566 19292 23572 19304
rect 21683 19264 23572 19292
rect 21683 19261 21695 19264
rect 21637 19255 21695 19261
rect 23566 19252 23572 19264
rect 23624 19252 23630 19304
rect 13863 19128 14136 19156
rect 13863 19125 13875 19128
rect 13817 19119 13875 19125
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 14829 19159 14887 19165
rect 14829 19156 14841 19159
rect 14792 19128 14841 19156
rect 14792 19116 14798 19128
rect 14829 19125 14841 19128
rect 14875 19125 14887 19159
rect 14829 19119 14887 19125
rect 15105 19159 15163 19165
rect 15105 19125 15117 19159
rect 15151 19156 15163 19159
rect 15470 19156 15476 19168
rect 15151 19128 15476 19156
rect 15151 19125 15163 19128
rect 15105 19119 15163 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15654 19156 15660 19168
rect 15615 19128 15660 19156
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17402 19156 17408 19168
rect 17359 19128 17408 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17402 19116 17408 19128
rect 17460 19156 17466 19168
rect 17773 19159 17831 19165
rect 17773 19156 17785 19159
rect 17460 19128 17785 19156
rect 17460 19116 17466 19128
rect 17773 19125 17785 19128
rect 17819 19125 17831 19159
rect 17773 19119 17831 19125
rect 18598 19116 18604 19168
rect 18656 19156 18662 19168
rect 19061 19159 19119 19165
rect 19061 19156 19073 19159
rect 18656 19128 19073 19156
rect 18656 19116 18662 19128
rect 19061 19125 19073 19128
rect 19107 19125 19119 19159
rect 19518 19156 19524 19168
rect 19479 19128 19524 19156
rect 19061 19119 19119 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20806 19156 20812 19168
rect 20404 19128 20812 19156
rect 20404 19116 20410 19128
rect 20806 19116 20812 19128
rect 20864 19156 20870 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20864 19128 20913 19156
rect 20864 19116 20870 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 14 18912 20 18964
rect 72 18952 78 18964
rect 5718 18952 5724 18964
rect 72 18924 5724 18952
rect 72 18912 78 18924
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 6733 18955 6791 18961
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 7282 18952 7288 18964
rect 6779 18924 7288 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 7282 18912 7288 18924
rect 7340 18952 7346 18964
rect 8297 18955 8355 18961
rect 7340 18924 7788 18952
rect 7340 18912 7346 18924
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 3602 18884 3608 18896
rect 2188 18856 3608 18884
rect 2188 18844 2194 18856
rect 3602 18844 3608 18856
rect 3660 18844 3666 18896
rect 4338 18884 4344 18896
rect 4264 18856 4344 18884
rect 2041 18819 2099 18825
rect 2041 18785 2053 18819
rect 2087 18816 2099 18819
rect 2222 18816 2228 18828
rect 2087 18788 2228 18816
rect 2087 18785 2099 18788
rect 2041 18779 2099 18785
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 2038 18640 2044 18692
rect 2096 18680 2102 18692
rect 2332 18680 2360 18779
rect 3234 18776 3240 18828
rect 3292 18816 3298 18828
rect 3329 18819 3387 18825
rect 3329 18816 3341 18819
rect 3292 18788 3341 18816
rect 3292 18776 3298 18788
rect 3329 18785 3341 18788
rect 3375 18816 3387 18819
rect 3878 18816 3884 18828
rect 3375 18788 3884 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 3878 18776 3884 18788
rect 3936 18776 3942 18828
rect 4264 18825 4292 18856
rect 4338 18844 4344 18856
rect 4396 18844 4402 18896
rect 5902 18884 5908 18896
rect 5815 18856 5908 18884
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18785 4307 18819
rect 4430 18816 4436 18828
rect 4389 18788 4436 18816
rect 4249 18779 4307 18785
rect 4430 18776 4436 18788
rect 4488 18825 4494 18828
rect 5828 18825 5856 18856
rect 5902 18844 5908 18856
rect 5960 18884 5966 18896
rect 7558 18884 7564 18896
rect 5960 18856 7564 18884
rect 5960 18844 5966 18856
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 4488 18819 4537 18825
rect 4488 18785 4491 18819
rect 4525 18785 4537 18819
rect 4488 18779 4537 18785
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18785 5871 18819
rect 6178 18816 6184 18828
rect 6139 18788 6184 18816
rect 5813 18779 5871 18785
rect 4488 18776 4522 18779
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 7190 18776 7196 18828
rect 7248 18816 7254 18828
rect 7469 18819 7527 18825
rect 7469 18816 7481 18819
rect 7248 18788 7481 18816
rect 7248 18776 7254 18788
rect 7469 18785 7481 18788
rect 7515 18785 7527 18819
rect 7650 18816 7656 18828
rect 7611 18788 7656 18816
rect 7469 18779 7527 18785
rect 2498 18748 2504 18760
rect 2459 18720 2504 18748
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 4494 18748 4522 18776
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 3844 18720 4629 18748
rect 3844 18708 3850 18720
rect 2869 18683 2927 18689
rect 2869 18680 2881 18683
rect 2096 18652 2881 18680
rect 2096 18640 2102 18652
rect 2869 18649 2881 18652
rect 2915 18680 2927 18683
rect 3878 18680 3884 18692
rect 2915 18652 3884 18680
rect 2915 18649 2927 18652
rect 2869 18643 2927 18649
rect 3878 18640 3884 18652
rect 3936 18680 3942 18692
rect 4494 18680 4522 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 5350 18708 5356 18760
rect 5408 18748 5414 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 5408 18720 5457 18748
rect 5408 18708 5414 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18748 6423 18751
rect 6454 18748 6460 18760
rect 6411 18720 6460 18748
rect 6411 18717 6423 18720
rect 6365 18711 6423 18717
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 7484 18748 7512 18779
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 7760 18816 7788 18924
rect 8297 18921 8309 18955
rect 8343 18952 8355 18955
rect 8386 18952 8392 18964
rect 8343 18924 8392 18952
rect 8343 18921 8355 18924
rect 8297 18915 8355 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 9907 18955 9965 18961
rect 8628 18924 9628 18952
rect 8628 18912 8634 18924
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 9600 18884 9628 18924
rect 9907 18921 9919 18955
rect 9953 18952 9965 18955
rect 12618 18952 12624 18964
rect 9953 18924 12624 18952
rect 9953 18921 9965 18924
rect 9907 18915 9965 18921
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 13170 18912 13176 18964
rect 13228 18952 13234 18964
rect 14001 18955 14059 18961
rect 14001 18952 14013 18955
rect 13228 18924 14013 18952
rect 13228 18912 13234 18924
rect 14001 18921 14013 18924
rect 14047 18952 14059 18955
rect 14182 18952 14188 18964
rect 14047 18924 14188 18952
rect 14047 18921 14059 18924
rect 14001 18915 14059 18921
rect 14182 18912 14188 18924
rect 14240 18912 14246 18964
rect 15105 18955 15163 18961
rect 15105 18921 15117 18955
rect 15151 18952 15163 18955
rect 15838 18952 15844 18964
rect 15151 18924 15844 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15838 18912 15844 18924
rect 15896 18952 15902 18964
rect 16301 18955 16359 18961
rect 16301 18952 16313 18955
rect 15896 18924 16313 18952
rect 15896 18912 15902 18924
rect 16301 18921 16313 18924
rect 16347 18921 16359 18955
rect 16301 18915 16359 18921
rect 16776 18924 18092 18952
rect 10229 18887 10287 18893
rect 10229 18884 10241 18887
rect 7892 18856 10241 18884
rect 7892 18844 7898 18856
rect 9600 18825 9628 18856
rect 10229 18853 10241 18856
rect 10275 18884 10287 18887
rect 10318 18884 10324 18896
rect 10275 18856 10324 18884
rect 10275 18853 10287 18856
rect 10229 18847 10287 18853
rect 10318 18844 10324 18856
rect 10376 18844 10382 18896
rect 12066 18884 12072 18896
rect 12027 18856 12072 18884
rect 12066 18844 12072 18856
rect 12124 18884 12130 18896
rect 12437 18887 12495 18893
rect 12437 18884 12449 18887
rect 12124 18856 12449 18884
rect 12124 18844 12130 18856
rect 12437 18853 12449 18856
rect 12483 18853 12495 18887
rect 12437 18847 12495 18853
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 7760 18788 9413 18816
rect 9401 18785 9413 18788
rect 9447 18785 9459 18819
rect 9401 18779 9459 18785
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18785 9643 18819
rect 9585 18779 9643 18785
rect 7558 18748 7564 18760
rect 7484 18720 7564 18748
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7926 18748 7932 18760
rect 7887 18720 7932 18748
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8628 18720 8953 18748
rect 8628 18708 8634 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 9416 18748 9444 18779
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 9804 18819 9862 18825
rect 9804 18816 9816 18819
rect 9732 18788 9816 18816
rect 9732 18776 9738 18788
rect 9804 18785 9816 18788
rect 9850 18785 9862 18819
rect 11054 18816 11060 18828
rect 11015 18788 11060 18816
rect 9804 18779 9862 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 11517 18819 11575 18825
rect 11517 18816 11529 18819
rect 11480 18788 11529 18816
rect 11480 18776 11486 18788
rect 11517 18785 11529 18788
rect 11563 18785 11575 18819
rect 12452 18816 12480 18847
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 12860 18856 13216 18884
rect 12860 18844 12866 18856
rect 12618 18816 12624 18828
rect 12452 18788 12624 18816
rect 11517 18779 11575 18785
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 12897 18819 12955 18825
rect 12897 18785 12909 18819
rect 12943 18785 12955 18819
rect 13078 18816 13084 18828
rect 13039 18788 13084 18816
rect 12897 18779 12955 18785
rect 9950 18748 9956 18760
rect 9416 18720 9956 18748
rect 8941 18711 8999 18717
rect 9950 18708 9956 18720
rect 10008 18748 10014 18760
rect 11793 18751 11851 18757
rect 10008 18720 11468 18748
rect 10008 18708 10014 18720
rect 6178 18680 6184 18692
rect 3936 18652 6184 18680
rect 3936 18640 3942 18652
rect 6178 18640 6184 18652
rect 6236 18640 6242 18692
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 10597 18683 10655 18689
rect 10597 18680 10609 18683
rect 6604 18652 10609 18680
rect 6604 18640 6610 18652
rect 10597 18649 10609 18652
rect 10643 18649 10655 18683
rect 11146 18680 11152 18692
rect 10597 18643 10655 18649
rect 11047 18652 11152 18680
rect 1670 18612 1676 18624
rect 1631 18584 1676 18612
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 5077 18615 5135 18621
rect 5077 18612 5089 18615
rect 4856 18584 5089 18612
rect 4856 18572 4862 18584
rect 5077 18581 5089 18584
rect 5123 18612 5135 18615
rect 5534 18612 5540 18624
rect 5123 18584 5540 18612
rect 5123 18581 5135 18584
rect 5077 18575 5135 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 7006 18612 7012 18624
rect 6967 18584 7012 18612
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 8573 18615 8631 18621
rect 8573 18612 8585 18615
rect 8444 18584 8585 18612
rect 8444 18572 8450 18584
rect 8573 18581 8585 18584
rect 8619 18581 8631 18615
rect 8573 18575 8631 18581
rect 8938 18572 8944 18624
rect 8996 18612 9002 18624
rect 11047 18612 11075 18652
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 11440 18680 11468 18720
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 12526 18748 12532 18760
rect 11839 18720 12532 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 12066 18680 12072 18692
rect 11440 18652 12072 18680
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 12912 18680 12940 18779
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 13188 18816 13216 18856
rect 13906 18844 13912 18896
rect 13964 18884 13970 18896
rect 14918 18884 14924 18896
rect 13964 18856 14924 18884
rect 13964 18844 13970 18856
rect 14918 18844 14924 18856
rect 14976 18884 14982 18896
rect 16022 18884 16028 18896
rect 14976 18856 15884 18884
rect 15983 18856 16028 18884
rect 14976 18844 14982 18856
rect 14252 18819 14310 18825
rect 13188 18788 13814 18816
rect 13262 18748 13268 18760
rect 13223 18720 13268 18748
rect 13262 18708 13268 18720
rect 13320 18708 13326 18760
rect 13786 18748 13814 18788
rect 14252 18785 14264 18819
rect 14298 18816 14310 18819
rect 15010 18816 15016 18828
rect 14298 18788 15016 18816
rect 14298 18785 14310 18788
rect 14252 18779 14310 18785
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15381 18819 15439 18825
rect 15381 18816 15393 18819
rect 15252 18788 15393 18816
rect 15252 18776 15258 18788
rect 15381 18785 15393 18788
rect 15427 18785 15439 18819
rect 15856 18816 15884 18856
rect 16022 18844 16028 18856
rect 16080 18844 16086 18896
rect 16776 18816 16804 18924
rect 17402 18884 17408 18896
rect 17328 18856 17408 18884
rect 16942 18816 16948 18828
rect 15856 18788 16804 18816
rect 16903 18788 16948 18816
rect 15381 18779 15439 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17218 18776 17224 18828
rect 17276 18816 17282 18828
rect 17328 18825 17356 18856
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 18064 18884 18092 18924
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18877 18955 18935 18961
rect 18877 18952 18889 18955
rect 18196 18924 18889 18952
rect 18196 18912 18202 18924
rect 18877 18921 18889 18924
rect 18923 18921 18935 18955
rect 18877 18915 18935 18921
rect 20806 18884 20812 18896
rect 18064 18856 20812 18884
rect 20806 18844 20812 18856
rect 20864 18884 20870 18896
rect 21085 18887 21143 18893
rect 21085 18884 21097 18887
rect 20864 18856 21097 18884
rect 20864 18844 20870 18856
rect 21085 18853 21097 18856
rect 21131 18853 21143 18887
rect 21085 18847 21143 18853
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 17276 18788 17325 18816
rect 17276 18776 17282 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18816 18199 18819
rect 18230 18816 18236 18828
rect 18187 18788 18236 18816
rect 18187 18785 18199 18788
rect 18141 18779 18199 18785
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 13786 18720 14657 18748
rect 14645 18717 14657 18720
rect 14691 18748 14703 18751
rect 16390 18748 16396 18760
rect 14691 18720 16396 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 17402 18748 17408 18760
rect 17363 18720 17408 18748
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 13814 18680 13820 18692
rect 12912 18652 13820 18680
rect 13814 18640 13820 18652
rect 13872 18640 13878 18692
rect 14182 18640 14188 18692
rect 14240 18680 14246 18692
rect 18156 18680 18184 18779
rect 18230 18776 18236 18788
rect 18288 18776 18294 18828
rect 18325 18819 18383 18825
rect 18325 18785 18337 18819
rect 18371 18816 18383 18819
rect 18414 18816 18420 18828
rect 18371 18788 18420 18816
rect 18371 18785 18383 18788
rect 18325 18779 18383 18785
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 19426 18816 19432 18828
rect 19387 18788 19432 18816
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 18555 18751 18613 18757
rect 18555 18717 18567 18751
rect 18601 18748 18613 18751
rect 19610 18748 19616 18760
rect 18601 18720 19616 18748
rect 18601 18717 18613 18720
rect 18555 18711 18613 18717
rect 19610 18708 19616 18720
rect 19668 18708 19674 18760
rect 20622 18708 20628 18760
rect 20680 18748 20686 18760
rect 20993 18751 21051 18757
rect 20993 18748 21005 18751
rect 20680 18720 21005 18748
rect 20680 18708 20686 18720
rect 20993 18717 21005 18720
rect 21039 18717 21051 18751
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 20993 18711 21051 18717
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 14240 18652 18184 18680
rect 14240 18640 14246 18652
rect 8996 18584 11075 18612
rect 8996 18572 9002 18584
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 12860 18584 13645 18612
rect 12860 18572 12866 18584
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 13909 18615 13967 18621
rect 13909 18581 13921 18615
rect 13955 18612 13967 18615
rect 14090 18612 14096 18624
rect 13955 18584 14096 18612
rect 13955 18581 13967 18584
rect 13909 18575 13967 18581
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14323 18615 14381 18621
rect 14323 18581 14335 18615
rect 14369 18612 14381 18615
rect 14550 18612 14556 18624
rect 14369 18584 14556 18612
rect 14369 18581 14381 18584
rect 14323 18575 14381 18581
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 19567 18615 19625 18621
rect 19567 18612 19579 18615
rect 16080 18584 19579 18612
rect 16080 18572 16086 18584
rect 19567 18581 19579 18584
rect 19613 18581 19625 18615
rect 19567 18575 19625 18581
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 3418 18417 3424 18420
rect 2777 18411 2835 18417
rect 2777 18377 2789 18411
rect 2823 18408 2835 18411
rect 3402 18411 3424 18417
rect 3402 18408 3414 18411
rect 2823 18380 3414 18408
rect 2823 18377 2835 18380
rect 2777 18371 2835 18377
rect 3402 18377 3414 18380
rect 3476 18408 3482 18420
rect 3602 18408 3608 18420
rect 3476 18380 3608 18408
rect 3402 18371 3424 18377
rect 3418 18368 3424 18371
rect 3476 18368 3482 18380
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 3878 18408 3884 18420
rect 3839 18380 3884 18408
rect 3878 18368 3884 18380
rect 3936 18368 3942 18420
rect 3970 18368 3976 18420
rect 4028 18368 4034 18420
rect 4338 18408 4344 18420
rect 4299 18380 4344 18408
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 5629 18411 5687 18417
rect 5629 18408 5641 18411
rect 4908 18380 5641 18408
rect 109 18343 167 18349
rect 109 18309 121 18343
rect 155 18340 167 18343
rect 3234 18340 3240 18352
rect 155 18312 3240 18340
rect 155 18309 167 18312
rect 109 18303 167 18309
rect 3234 18300 3240 18312
rect 3292 18340 3298 18352
rect 3513 18343 3571 18349
rect 3513 18340 3525 18343
rect 3292 18312 3525 18340
rect 3292 18300 3298 18312
rect 3513 18309 3525 18312
rect 3559 18309 3571 18343
rect 3988 18340 4016 18368
rect 4908 18352 4936 18380
rect 5629 18377 5641 18380
rect 5675 18377 5687 18411
rect 5902 18408 5908 18420
rect 5863 18380 5908 18408
rect 5629 18371 5687 18377
rect 5902 18368 5908 18380
rect 5960 18368 5966 18420
rect 6178 18408 6184 18420
rect 6139 18380 6184 18408
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 9490 18408 9496 18420
rect 7616 18380 9496 18408
rect 7616 18368 7622 18380
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 9585 18411 9643 18417
rect 9585 18377 9597 18411
rect 9631 18408 9643 18411
rect 9674 18408 9680 18420
rect 9631 18380 9680 18408
rect 9631 18377 9643 18380
rect 9585 18371 9643 18377
rect 9674 18368 9680 18380
rect 9732 18408 9738 18420
rect 9769 18411 9827 18417
rect 9769 18408 9781 18411
rect 9732 18380 9781 18408
rect 9732 18368 9738 18380
rect 9769 18377 9781 18380
rect 9815 18377 9827 18411
rect 9769 18371 9827 18377
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 11054 18408 11060 18420
rect 10008 18380 11060 18408
rect 10008 18368 10014 18380
rect 11054 18368 11060 18380
rect 11112 18368 11118 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 12253 18411 12311 18417
rect 12253 18408 12265 18411
rect 11204 18380 12265 18408
rect 11204 18368 11210 18380
rect 12253 18377 12265 18380
rect 12299 18408 12311 18411
rect 12342 18408 12348 18420
rect 12299 18380 12348 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 12342 18368 12348 18380
rect 12400 18408 12406 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 12400 18380 14841 18408
rect 12400 18368 12406 18380
rect 4890 18340 4896 18352
rect 3988 18312 4896 18340
rect 3513 18303 3571 18309
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 5920 18340 5948 18368
rect 10226 18340 10232 18352
rect 5184 18312 5948 18340
rect 6012 18312 10232 18340
rect 3145 18275 3203 18281
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3326 18272 3332 18284
rect 3191 18244 3332 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 3326 18232 3332 18244
rect 3384 18272 3390 18284
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 3384 18244 3617 18272
rect 3384 18232 3390 18244
rect 3605 18241 3617 18244
rect 3651 18272 3663 18275
rect 3970 18272 3976 18284
rect 3651 18244 3976 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 3970 18232 3976 18244
rect 4028 18232 4034 18284
rect 1670 18204 1676 18216
rect 1583 18176 1676 18204
rect 1670 18164 1676 18176
rect 1728 18164 1734 18216
rect 1949 18207 2007 18213
rect 1949 18173 1961 18207
rect 1995 18204 2007 18207
rect 2038 18204 2044 18216
rect 1995 18176 2044 18204
rect 1995 18173 2007 18176
rect 1949 18167 2007 18173
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 3418 18164 3424 18216
rect 3476 18204 3482 18216
rect 4246 18204 4252 18216
rect 3476 18176 4252 18204
rect 3476 18164 3482 18176
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18204 4767 18207
rect 5077 18207 5135 18213
rect 5077 18204 5089 18207
rect 4755 18176 5089 18204
rect 4755 18173 4767 18176
rect 4709 18167 4767 18173
rect 5077 18173 5089 18176
rect 5123 18204 5135 18207
rect 5184 18204 5212 18312
rect 5350 18272 5356 18284
rect 5311 18244 5356 18272
rect 5350 18232 5356 18244
rect 5408 18232 5414 18284
rect 5442 18232 5448 18284
rect 5500 18272 5506 18284
rect 6012 18272 6040 18312
rect 10226 18300 10232 18312
rect 10284 18300 10290 18352
rect 7374 18272 7380 18284
rect 5500 18244 6040 18272
rect 6380 18244 7380 18272
rect 5500 18232 5506 18244
rect 5123 18176 5212 18204
rect 5123 18173 5135 18176
rect 5077 18167 5135 18173
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5629 18207 5687 18213
rect 5316 18176 5361 18204
rect 5316 18164 5322 18176
rect 5629 18173 5641 18207
rect 5675 18204 5687 18207
rect 6380 18204 6408 18244
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 11422 18272 11428 18284
rect 7616 18244 7741 18272
rect 7616 18232 7622 18244
rect 5675 18176 6408 18204
rect 6457 18207 6515 18213
rect 5675 18173 5687 18176
rect 5629 18167 5687 18173
rect 6457 18173 6469 18207
rect 6503 18204 6515 18207
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6503 18176 6837 18204
rect 6503 18173 6515 18176
rect 6457 18167 6515 18173
rect 6825 18173 6837 18176
rect 6871 18204 6883 18207
rect 7190 18204 7196 18216
rect 6871 18176 7196 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 934 18028 940 18080
rect 992 18068 998 18080
rect 1489 18071 1547 18077
rect 1489 18068 1501 18071
rect 992 18040 1501 18068
rect 992 18028 998 18040
rect 1489 18037 1501 18040
rect 1535 18037 1547 18071
rect 1688 18068 1716 18164
rect 2774 18096 2780 18148
rect 2832 18136 2838 18148
rect 3234 18136 3240 18148
rect 2832 18108 3240 18136
rect 2832 18096 2838 18108
rect 3234 18096 3240 18108
rect 3292 18096 3298 18148
rect 3694 18096 3700 18148
rect 3752 18096 3758 18148
rect 5276 18136 5304 18164
rect 7006 18136 7012 18148
rect 5276 18108 7012 18136
rect 7006 18096 7012 18108
rect 7064 18136 7070 18148
rect 7300 18136 7328 18167
rect 7558 18136 7564 18148
rect 7064 18108 7328 18136
rect 7519 18108 7564 18136
rect 7064 18096 7070 18108
rect 7558 18096 7564 18108
rect 7616 18096 7622 18148
rect 3712 18068 3740 18096
rect 1688 18040 3740 18068
rect 1489 18031 1547 18037
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 6457 18071 6515 18077
rect 6457 18068 6469 18071
rect 4396 18040 6469 18068
rect 4396 18028 4402 18040
rect 6457 18037 6469 18040
rect 6503 18068 6515 18071
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 6503 18040 6561 18068
rect 6503 18037 6515 18040
rect 6457 18031 6515 18037
rect 6549 18037 6561 18040
rect 6595 18037 6607 18071
rect 7713 18068 7741 18244
rect 8956 18244 11428 18272
rect 7834 18164 7840 18216
rect 7892 18204 7898 18216
rect 8956 18213 8984 18244
rect 11422 18232 11428 18244
rect 11480 18272 11486 18284
rect 11609 18275 11667 18281
rect 11609 18272 11621 18275
rect 11480 18244 11621 18272
rect 11480 18232 11486 18244
rect 11609 18241 11621 18244
rect 11655 18241 11667 18275
rect 11609 18235 11667 18241
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 7892 18176 8401 18204
rect 7892 18164 7898 18176
rect 7834 18068 7840 18080
rect 7713 18040 7840 18068
rect 6549 18031 6607 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 8220 18077 8248 18176
rect 8389 18173 8401 18176
rect 8435 18173 8447 18207
rect 8389 18167 8447 18173
rect 8941 18207 8999 18213
rect 8941 18173 8953 18207
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 8294 18096 8300 18148
rect 8352 18136 8358 18148
rect 8956 18136 8984 18167
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9950 18204 9956 18216
rect 9088 18176 9956 18204
rect 9088 18164 9094 18176
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 10318 18204 10324 18216
rect 10279 18176 10324 18204
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 12636 18213 12664 18380
rect 14829 18377 14841 18380
rect 14875 18377 14887 18411
rect 14829 18371 14887 18377
rect 15194 18368 15200 18420
rect 15252 18408 15258 18420
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 15252 18380 15393 18408
rect 15252 18368 15258 18380
rect 15381 18377 15393 18380
rect 15427 18377 15439 18411
rect 15381 18371 15439 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 16942 18408 16948 18420
rect 15528 18380 16948 18408
rect 15528 18368 15534 18380
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 19242 18368 19248 18420
rect 19300 18408 19306 18420
rect 19702 18408 19708 18420
rect 19300 18380 19708 18408
rect 19300 18368 19306 18380
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 21315 18411 21373 18417
rect 21315 18408 21327 18411
rect 20128 18380 21327 18408
rect 20128 18368 20134 18380
rect 21315 18377 21327 18380
rect 21361 18377 21373 18411
rect 21315 18371 21373 18377
rect 14090 18300 14096 18352
rect 14148 18340 14154 18352
rect 16850 18340 16856 18352
rect 14148 18312 16856 18340
rect 14148 18300 14154 18312
rect 16850 18300 16856 18312
rect 16908 18300 16914 18352
rect 18506 18300 18512 18352
rect 18564 18340 18570 18352
rect 18564 18312 20024 18340
rect 18564 18300 18570 18312
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 19705 18275 19763 18281
rect 19705 18272 19717 18275
rect 14608 18244 19717 18272
rect 14608 18232 14614 18244
rect 19705 18241 19717 18244
rect 19751 18272 19763 18275
rect 19794 18272 19800 18284
rect 19751 18244 19800 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 19794 18232 19800 18244
rect 19852 18232 19858 18284
rect 19996 18281 20024 18312
rect 20254 18300 20260 18352
rect 20312 18340 20318 18352
rect 20312 18312 20392 18340
rect 20312 18300 20318 18312
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18173 12679 18207
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12621 18167 12679 18173
rect 8352 18108 8984 18136
rect 9125 18139 9183 18145
rect 8352 18096 8358 18108
rect 9125 18105 9137 18139
rect 9171 18105 9183 18139
rect 9125 18099 9183 18105
rect 9493 18139 9551 18145
rect 9493 18105 9505 18139
rect 9539 18136 9551 18139
rect 10042 18136 10048 18148
rect 9539 18108 10048 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 8205 18071 8263 18077
rect 8205 18037 8217 18071
rect 8251 18068 8263 18071
rect 8846 18068 8852 18080
rect 8251 18040 8852 18068
rect 8251 18037 8263 18040
rect 8205 18031 8263 18037
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9140 18068 9168 18099
rect 10042 18096 10048 18108
rect 10100 18136 10106 18148
rect 10594 18136 10600 18148
rect 10100 18108 10600 18136
rect 10100 18096 10106 18108
rect 10594 18096 10600 18108
rect 10652 18136 10658 18148
rect 10704 18136 10732 18167
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18173 14335 18207
rect 14458 18204 14464 18216
rect 14419 18176 14464 18204
rect 14277 18167 14335 18173
rect 10652 18108 10732 18136
rect 10652 18096 10658 18108
rect 12710 18096 12716 18148
rect 12768 18136 12774 18148
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 12768 18108 13921 18136
rect 12768 18096 12774 18108
rect 13909 18105 13921 18108
rect 13955 18136 13967 18139
rect 14292 18136 14320 18167
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18204 14887 18207
rect 15841 18207 15899 18213
rect 14875 18176 15792 18204
rect 14875 18173 14887 18176
rect 14829 18167 14887 18173
rect 14734 18136 14740 18148
rect 13955 18108 14740 18136
rect 13955 18105 13967 18108
rect 13909 18099 13967 18105
rect 14734 18096 14740 18108
rect 14792 18136 14798 18148
rect 15764 18136 15792 18176
rect 15841 18173 15853 18207
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18204 16175 18207
rect 16298 18204 16304 18216
rect 16163 18176 16304 18204
rect 16163 18173 16175 18176
rect 16117 18167 16175 18173
rect 15856 18136 15884 18167
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 16393 18207 16451 18213
rect 16393 18173 16405 18207
rect 16439 18204 16451 18207
rect 17865 18207 17923 18213
rect 17865 18204 17877 18207
rect 16439 18176 17877 18204
rect 16439 18173 16451 18176
rect 16393 18167 16451 18173
rect 17865 18173 17877 18176
rect 17911 18204 17923 18207
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17911 18176 18061 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 18049 18173 18061 18176
rect 18095 18204 18107 18207
rect 18138 18204 18144 18216
rect 18095 18176 18144 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 18322 18164 18328 18216
rect 18380 18204 18386 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18380 18176 18521 18204
rect 18380 18164 18386 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 20364 18204 20392 18312
rect 20806 18300 20812 18352
rect 20864 18340 20870 18352
rect 20901 18343 20959 18349
rect 20901 18340 20913 18343
rect 20864 18312 20913 18340
rect 20864 18300 20870 18312
rect 20901 18309 20913 18312
rect 20947 18309 20959 18343
rect 20901 18303 20959 18309
rect 21212 18207 21270 18213
rect 21212 18204 21224 18207
rect 20364 18176 21224 18204
rect 18509 18167 18567 18173
rect 21212 18173 21224 18176
rect 21258 18204 21270 18207
rect 21637 18207 21695 18213
rect 21637 18204 21649 18207
rect 21258 18176 21649 18204
rect 21258 18173 21270 18176
rect 21212 18167 21270 18173
rect 21637 18173 21649 18176
rect 21683 18204 21695 18207
rect 22186 18204 22192 18216
rect 21683 18176 22192 18204
rect 21683 18173 21695 18176
rect 21637 18167 21695 18173
rect 22186 18164 22192 18176
rect 22244 18164 22250 18216
rect 14792 18108 16712 18136
rect 14792 18096 14798 18108
rect 9582 18068 9588 18080
rect 9140 18040 9588 18068
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10226 18028 10232 18080
rect 10284 18068 10290 18080
rect 10321 18071 10379 18077
rect 10321 18068 10333 18071
rect 10284 18040 10333 18068
rect 10284 18028 10290 18040
rect 10321 18037 10333 18040
rect 10367 18037 10379 18071
rect 10321 18031 10379 18037
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 11112 18040 11345 18068
rect 11112 18028 11118 18040
rect 11333 18037 11345 18040
rect 11379 18068 11391 18071
rect 11790 18068 11796 18080
rect 11379 18040 11796 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 12529 18071 12587 18077
rect 12529 18068 12541 18071
rect 12400 18040 12541 18068
rect 12400 18028 12406 18040
rect 12529 18037 12541 18040
rect 12575 18037 12587 18071
rect 12529 18031 12587 18037
rect 13541 18071 13599 18077
rect 13541 18037 13553 18071
rect 13587 18068 13599 18071
rect 13814 18068 13820 18080
rect 13587 18040 13820 18068
rect 13587 18037 13599 18040
rect 13541 18031 13599 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14090 18068 14096 18080
rect 14051 18040 14096 18068
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 15010 18068 15016 18080
rect 14971 18040 15016 18068
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15194 18028 15200 18080
rect 15252 18068 15258 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 15252 18040 15669 18068
rect 15252 18028 15258 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 15764 18068 15792 18108
rect 16684 18080 16712 18108
rect 16758 18096 16764 18148
rect 16816 18136 16822 18148
rect 17218 18136 17224 18148
rect 16816 18108 17224 18136
rect 16816 18096 16822 18108
rect 17218 18096 17224 18108
rect 17276 18136 17282 18148
rect 17313 18139 17371 18145
rect 17313 18136 17325 18139
rect 17276 18108 17325 18136
rect 17276 18096 17282 18108
rect 17313 18105 17325 18108
rect 17359 18105 17371 18139
rect 17313 18099 17371 18105
rect 19797 18139 19855 18145
rect 19797 18105 19809 18139
rect 19843 18136 19855 18139
rect 20530 18136 20536 18148
rect 19843 18108 20536 18136
rect 19843 18105 19855 18108
rect 19797 18099 19855 18105
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 15764 18040 16405 18068
rect 15657 18031 15715 18037
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 16666 18068 16672 18080
rect 16627 18040 16672 18068
rect 16393 18031 16451 18037
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18141 18071 18199 18077
rect 18141 18068 18153 18071
rect 17920 18040 18153 18068
rect 17920 18028 17926 18040
rect 18141 18037 18153 18040
rect 18187 18037 18199 18071
rect 18141 18031 18199 18037
rect 18414 18028 18420 18080
rect 18472 18068 18478 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 18472 18040 19073 18068
rect 18472 18028 18478 18040
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19061 18031 19119 18037
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 19300 18040 19441 18068
rect 19300 18028 19306 18040
rect 19429 18037 19441 18040
rect 19475 18068 19487 18071
rect 19812 18068 19840 18099
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 20622 18096 20628 18148
rect 20680 18136 20686 18148
rect 22005 18139 22063 18145
rect 22005 18136 22017 18139
rect 20680 18108 22017 18136
rect 20680 18096 20686 18108
rect 22005 18105 22017 18108
rect 22051 18105 22063 18139
rect 22005 18099 22063 18105
rect 19475 18040 19840 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 937 17867 995 17873
rect 937 17833 949 17867
rect 983 17864 995 17867
rect 1670 17864 1676 17876
rect 983 17836 1676 17864
rect 983 17833 995 17836
rect 937 17827 995 17833
rect 1479 17737 1507 17836
rect 1670 17824 1676 17836
rect 1728 17864 1734 17876
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1728 17836 1869 17864
rect 1728 17824 1734 17836
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 3878 17864 3884 17876
rect 3839 17836 3884 17864
rect 1857 17827 1915 17833
rect 3878 17824 3884 17836
rect 3936 17864 3942 17876
rect 3936 17836 4292 17864
rect 3936 17824 3942 17836
rect 3142 17756 3148 17808
rect 3200 17796 3206 17808
rect 3326 17796 3332 17808
rect 3200 17768 3332 17796
rect 3200 17756 3206 17768
rect 3326 17756 3332 17768
rect 3384 17756 3390 17808
rect 1464 17731 1522 17737
rect 1464 17697 1476 17731
rect 1510 17697 1522 17731
rect 2682 17728 2688 17740
rect 2643 17700 2688 17728
rect 1464 17691 1522 17697
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 2866 17688 2872 17740
rect 2924 17728 2930 17740
rect 2961 17731 3019 17737
rect 2961 17728 2973 17731
rect 2924 17700 2973 17728
rect 2924 17688 2930 17700
rect 2961 17697 2973 17700
rect 3007 17728 3019 17731
rect 3896 17728 3924 17824
rect 4264 17805 4292 17836
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 6273 17867 6331 17873
rect 6273 17864 6285 17867
rect 4764 17836 6285 17864
rect 4764 17824 4770 17836
rect 6273 17833 6285 17836
rect 6319 17833 6331 17867
rect 6638 17864 6644 17876
rect 6599 17836 6644 17864
rect 6273 17827 6331 17833
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 6822 17824 6828 17876
rect 6880 17864 6886 17876
rect 7466 17864 7472 17876
rect 6880 17836 7472 17864
rect 6880 17824 6886 17836
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 8389 17867 8447 17873
rect 8389 17864 8401 17867
rect 8352 17836 8401 17864
rect 8352 17824 8358 17836
rect 8389 17833 8401 17836
rect 8435 17833 8447 17867
rect 8389 17827 8447 17833
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 8904 17836 10149 17864
rect 8904 17824 8910 17836
rect 10137 17833 10149 17836
rect 10183 17833 10195 17867
rect 11422 17864 11428 17876
rect 11383 17836 11428 17864
rect 10137 17827 10195 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 11514 17824 11520 17876
rect 11572 17864 11578 17876
rect 11701 17867 11759 17873
rect 11701 17864 11713 17867
rect 11572 17836 11713 17864
rect 11572 17824 11578 17836
rect 11701 17833 11713 17836
rect 11747 17833 11759 17867
rect 11701 17827 11759 17833
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 15381 17867 15439 17873
rect 15381 17864 15393 17867
rect 12492 17836 15393 17864
rect 12492 17824 12498 17836
rect 15381 17833 15393 17836
rect 15427 17833 15439 17867
rect 15381 17827 15439 17833
rect 15562 17824 15568 17876
rect 15620 17864 15626 17876
rect 16298 17864 16304 17876
rect 15620 17836 16304 17864
rect 15620 17824 15626 17836
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 18046 17864 18052 17876
rect 17644 17836 18052 17864
rect 17644 17824 17650 17836
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18141 17867 18199 17873
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 18322 17864 18328 17876
rect 18187 17836 18328 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 18506 17864 18512 17876
rect 18467 17836 18512 17864
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 19794 17864 19800 17876
rect 19755 17836 19800 17864
rect 19794 17824 19800 17836
rect 19852 17824 19858 17876
rect 19978 17824 19984 17876
rect 20036 17864 20042 17876
rect 20993 17867 21051 17873
rect 20993 17864 21005 17867
rect 20036 17836 21005 17864
rect 20036 17824 20042 17836
rect 20993 17833 21005 17836
rect 21039 17833 21051 17867
rect 20993 17827 21051 17833
rect 4249 17799 4307 17805
rect 4249 17765 4261 17799
rect 4295 17765 4307 17799
rect 4249 17759 4307 17765
rect 4614 17756 4620 17808
rect 4672 17796 4678 17808
rect 9033 17799 9091 17805
rect 9033 17796 9045 17799
rect 4672 17768 9045 17796
rect 4672 17756 4678 17768
rect 9033 17765 9045 17768
rect 9079 17765 9091 17799
rect 9033 17759 9091 17765
rect 10318 17756 10324 17808
rect 10376 17796 10382 17808
rect 10870 17796 10876 17808
rect 10376 17768 10876 17796
rect 10376 17756 10382 17768
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 11440 17796 11468 17824
rect 12710 17796 12716 17808
rect 11440 17768 12716 17796
rect 3007 17700 3924 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 4890 17688 4896 17740
rect 4948 17728 4954 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 4948 17700 4997 17728
rect 4948 17688 4954 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 4985 17691 5043 17697
rect 5258 17688 5264 17740
rect 5316 17728 5322 17740
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 5316 17700 5457 17728
rect 5316 17688 5322 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 6822 17728 6828 17740
rect 6783 17700 6828 17728
rect 5445 17691 5503 17697
rect 3142 17660 3148 17672
rect 3103 17632 3148 17660
rect 3142 17620 3148 17632
rect 3200 17620 3206 17672
rect 3694 17620 3700 17672
rect 3752 17660 3758 17672
rect 5166 17660 5172 17672
rect 3752 17632 5172 17660
rect 3752 17620 3758 17632
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 2222 17552 2228 17604
rect 2280 17592 2286 17604
rect 2317 17595 2375 17601
rect 2317 17592 2329 17595
rect 2280 17564 2329 17592
rect 2280 17552 2286 17564
rect 2317 17561 2329 17564
rect 2363 17592 2375 17595
rect 4246 17592 4252 17604
rect 2363 17564 4252 17592
rect 2363 17561 2375 17564
rect 2317 17555 2375 17561
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 293 17527 351 17533
rect 293 17493 305 17527
rect 339 17524 351 17527
rect 1486 17524 1492 17536
rect 339 17496 1492 17524
rect 339 17493 351 17496
rect 293 17487 351 17493
rect 1486 17484 1492 17496
rect 1544 17533 1550 17536
rect 1544 17527 1593 17533
rect 1544 17493 1547 17527
rect 1581 17493 1593 17527
rect 1544 17487 1593 17493
rect 1544 17484 1550 17487
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3513 17527 3571 17533
rect 3513 17524 3525 17527
rect 3292 17496 3525 17524
rect 3292 17484 3298 17496
rect 3513 17493 3525 17496
rect 3559 17524 3571 17527
rect 4062 17524 4068 17536
rect 3559 17496 4068 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4430 17484 4436 17536
rect 4488 17524 4494 17536
rect 4893 17527 4951 17533
rect 4893 17524 4905 17527
rect 4488 17496 4905 17524
rect 4488 17484 4494 17496
rect 4893 17493 4905 17496
rect 4939 17524 4951 17527
rect 5460 17524 5488 17691
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6972 17700 7021 17728
rect 6972 17688 6978 17700
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 8608 17731 8666 17737
rect 8608 17728 8620 17731
rect 7009 17691 7067 17697
rect 8036 17700 8620 17728
rect 5626 17660 5632 17672
rect 5587 17632 5632 17660
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 6328 17632 7941 17660
rect 6328 17620 6334 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 5810 17552 5816 17604
rect 5868 17592 5874 17604
rect 6365 17595 6423 17601
rect 6365 17592 6377 17595
rect 5868 17564 6377 17592
rect 5868 17552 5874 17564
rect 6365 17561 6377 17564
rect 6411 17561 6423 17595
rect 8036 17592 8064 17700
rect 8608 17697 8620 17700
rect 8654 17728 8666 17731
rect 9214 17728 9220 17740
rect 8654 17700 9220 17728
rect 8654 17697 8666 17700
rect 8608 17691 8666 17697
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9732 17700 10057 17728
rect 9732 17688 9738 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10594 17728 10600 17740
rect 10555 17700 10600 17728
rect 10045 17691 10103 17697
rect 10594 17688 10600 17700
rect 10652 17688 10658 17740
rect 11606 17728 11612 17740
rect 11567 17700 11612 17728
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 12084 17737 12112 17768
rect 12710 17756 12716 17768
rect 12768 17796 12774 17808
rect 12894 17796 12900 17808
rect 12768 17768 12900 17796
rect 12768 17756 12774 17768
rect 12894 17756 12900 17768
rect 12952 17796 12958 17808
rect 12989 17799 13047 17805
rect 12989 17796 13001 17799
rect 12952 17768 13001 17796
rect 12952 17756 12958 17768
rect 12989 17765 13001 17768
rect 13035 17796 13047 17799
rect 13035 17768 13676 17796
rect 13035 17765 13047 17768
rect 12989 17759 13047 17765
rect 12069 17731 12127 17737
rect 12069 17697 12081 17731
rect 12115 17697 12127 17731
rect 12618 17728 12624 17740
rect 12579 17700 12624 17728
rect 12069 17691 12127 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 13170 17728 13176 17740
rect 13131 17700 13176 17728
rect 13170 17688 13176 17700
rect 13228 17728 13234 17740
rect 13538 17728 13544 17740
rect 13228 17700 13544 17728
rect 13228 17688 13234 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13648 17737 13676 17768
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 16853 17799 16911 17805
rect 16853 17796 16865 17799
rect 14976 17768 16865 17796
rect 14976 17756 14982 17768
rect 16853 17765 16865 17768
rect 16899 17765 16911 17799
rect 18340 17796 18368 17824
rect 18340 17768 18920 17796
rect 16853 17759 16911 17765
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17697 13691 17731
rect 13633 17691 13691 17697
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13872 17700 14289 17728
rect 13872 17688 13878 17700
rect 14277 17697 14289 17700
rect 14323 17728 14335 17731
rect 14458 17728 14464 17740
rect 14323 17700 14464 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 14458 17688 14464 17700
rect 14516 17728 14522 17740
rect 14642 17728 14648 17740
rect 14516 17700 14648 17728
rect 14516 17688 14522 17700
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 15470 17728 15476 17740
rect 15431 17700 15476 17728
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15841 17731 15899 17737
rect 15841 17697 15853 17731
rect 15887 17697 15899 17731
rect 17494 17728 17500 17740
rect 17455 17700 17500 17728
rect 15841 17691 15899 17697
rect 12802 17660 12808 17672
rect 6365 17555 6423 17561
rect 7202 17564 8064 17592
rect 8220 17632 12808 17660
rect 5718 17524 5724 17536
rect 4939 17496 5724 17524
rect 4939 17493 4951 17496
rect 4893 17487 4951 17493
rect 5718 17484 5724 17496
rect 5776 17524 5782 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5776 17496 6009 17524
rect 5776 17484 5782 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 6273 17527 6331 17533
rect 6273 17493 6285 17527
rect 6319 17524 6331 17527
rect 7202 17524 7230 17564
rect 7650 17524 7656 17536
rect 6319 17496 7230 17524
rect 7563 17496 7656 17524
rect 6319 17493 6331 17496
rect 6273 17487 6331 17493
rect 7650 17484 7656 17496
rect 7708 17524 7714 17536
rect 8220 17524 8248 17632
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 15102 17660 15108 17672
rect 14139 17632 15108 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 15102 17620 15108 17632
rect 15160 17660 15166 17672
rect 15856 17660 15884 17691
rect 17494 17688 17500 17700
rect 17552 17688 17558 17740
rect 18233 17731 18291 17737
rect 18233 17697 18245 17731
rect 18279 17728 18291 17731
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 18279 17700 18429 17728
rect 18279 17697 18291 17700
rect 18233 17691 18291 17697
rect 18417 17697 18429 17700
rect 18463 17728 18475 17731
rect 18598 17728 18604 17740
rect 18463 17700 18604 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 18598 17688 18604 17700
rect 18656 17688 18662 17740
rect 18892 17737 18920 17768
rect 19058 17756 19064 17808
rect 19116 17796 19122 17808
rect 20070 17796 20076 17808
rect 19116 17768 20076 17796
rect 19116 17756 19122 17768
rect 20070 17756 20076 17768
rect 20128 17756 20134 17808
rect 18877 17731 18935 17737
rect 18877 17697 18889 17731
rect 18923 17697 18935 17731
rect 18877 17691 18935 17697
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20864 17700 20913 17728
rect 20864 17688 20870 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 21450 17728 21456 17740
rect 21411 17700 21456 17728
rect 20901 17691 20959 17697
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 15160 17632 18368 17660
rect 15160 17620 15166 17632
rect 9861 17595 9919 17601
rect 9861 17561 9873 17595
rect 9907 17592 9919 17595
rect 10042 17592 10048 17604
rect 9907 17564 10048 17592
rect 9907 17561 9919 17564
rect 9861 17555 9919 17561
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 10870 17552 10876 17604
rect 10928 17592 10934 17604
rect 14921 17595 14979 17601
rect 14921 17592 14933 17595
rect 10928 17564 14933 17592
rect 10928 17552 10934 17564
rect 14921 17561 14933 17564
rect 14967 17561 14979 17595
rect 14921 17555 14979 17561
rect 15838 17552 15844 17604
rect 15896 17592 15902 17604
rect 18233 17595 18291 17601
rect 18233 17592 18245 17595
rect 15896 17564 18245 17592
rect 15896 17552 15902 17564
rect 18233 17561 18245 17564
rect 18279 17561 18291 17595
rect 18340 17592 18368 17632
rect 21450 17592 21456 17604
rect 18340 17564 21456 17592
rect 18233 17555 18291 17561
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 7708 17496 8248 17524
rect 8711 17527 8769 17533
rect 7708 17484 7714 17496
rect 8711 17493 8723 17527
rect 8757 17524 8769 17527
rect 8846 17524 8852 17536
rect 8757 17496 8852 17524
rect 8757 17493 8769 17496
rect 8711 17487 8769 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 9401 17527 9459 17533
rect 9401 17524 9413 17527
rect 9364 17496 9413 17524
rect 9364 17484 9370 17496
rect 9401 17493 9413 17496
rect 9447 17493 9459 17527
rect 9401 17487 9459 17493
rect 9950 17484 9956 17536
rect 10008 17524 10014 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10008 17496 11069 17524
rect 10008 17484 10014 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 12676 17496 14105 17524
rect 12676 17484 12682 17496
rect 14093 17493 14105 17496
rect 14139 17493 14151 17527
rect 14550 17524 14556 17536
rect 14511 17496 14556 17524
rect 14093 17487 14151 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 16758 17524 16764 17536
rect 16719 17496 16764 17524
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 19426 17524 19432 17536
rect 18656 17496 19432 17524
rect 18656 17484 18662 17496
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 14 17416 20 17468
rect 72 17456 78 17468
rect 72 17428 117 17456
rect 1104 17434 22816 17456
rect 72 17416 78 17428
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 17 17323 75 17329
rect 17 17289 29 17323
rect 63 17320 75 17323
rect 2222 17320 2228 17332
rect 63 17292 2228 17320
rect 63 17289 75 17292
rect 17 17283 75 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2682 17320 2688 17332
rect 2547 17292 2688 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 2866 17320 2872 17332
rect 2827 17292 2872 17320
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 3329 17323 3387 17329
rect 3329 17289 3341 17323
rect 3375 17320 3387 17323
rect 4338 17320 4344 17332
rect 3375 17292 4344 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 6178 17320 6184 17332
rect 4479 17292 6184 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 6178 17280 6184 17292
rect 6236 17280 6242 17332
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 8110 17320 8116 17332
rect 6512 17292 8116 17320
rect 6512 17280 6518 17292
rect 8110 17280 8116 17292
rect 8168 17280 8174 17332
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 8352 17292 8978 17320
rect 8352 17280 8358 17292
rect 2038 17212 2044 17264
rect 2096 17252 2102 17264
rect 4706 17252 4712 17264
rect 2096 17224 4712 17252
rect 2096 17212 2102 17224
rect 4706 17212 4712 17224
rect 4764 17252 4770 17264
rect 6641 17255 6699 17261
rect 6641 17252 6653 17255
rect 4764 17224 6653 17252
rect 4764 17212 4770 17224
rect 6641 17221 6653 17224
rect 6687 17252 6699 17255
rect 6822 17252 6828 17264
rect 6687 17224 6828 17252
rect 6687 17221 6699 17224
rect 6641 17215 6699 17221
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 7466 17252 7472 17264
rect 7427 17224 7472 17252
rect 7466 17212 7472 17224
rect 7524 17252 7530 17264
rect 8950 17252 8978 17292
rect 9214 17280 9220 17332
rect 9272 17320 9278 17332
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 9272 17292 9413 17320
rect 9272 17280 9278 17292
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 9732 17292 9965 17320
rect 9732 17280 9738 17292
rect 9953 17289 9965 17292
rect 9999 17320 10011 17323
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9999 17292 10057 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10045 17289 10057 17292
rect 10091 17289 10103 17323
rect 13538 17320 13544 17332
rect 13499 17292 13544 17320
rect 10045 17283 10103 17289
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17320 13783 17323
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13771 17292 13829 17320
rect 13771 17289 13783 17292
rect 13725 17283 13783 17289
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 16761 17323 16819 17329
rect 16761 17320 16773 17323
rect 13817 17283 13875 17289
rect 14660 17292 16773 17320
rect 10597 17255 10655 17261
rect 10597 17252 10609 17255
rect 7524 17224 8800 17252
rect 8950 17224 10609 17252
rect 7524 17212 7530 17224
rect 2056 17184 2084 17212
rect 1688 17156 2084 17184
rect 3513 17187 3571 17193
rect 1688 17125 1716 17156
rect 3513 17153 3525 17187
rect 3559 17184 3571 17187
rect 4154 17184 4160 17196
rect 3559 17156 4160 17184
rect 3559 17153 3571 17156
rect 3513 17147 3571 17153
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 2406 17116 2412 17128
rect 1995 17088 2412 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2406 17076 2412 17088
rect 2464 17116 2470 17128
rect 2866 17116 2872 17128
rect 2464 17088 2872 17116
rect 2464 17076 2470 17088
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3896 17125 3924 17156
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4246 17144 4252 17196
rect 4304 17184 4310 17196
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 4304 17156 5089 17184
rect 4304 17144 4310 17156
rect 5077 17153 5089 17156
rect 5123 17184 5135 17187
rect 6178 17184 6184 17196
rect 5123 17156 6184 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17085 3939 17119
rect 3881 17079 3939 17085
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 4028 17088 4077 17116
rect 4028 17076 4034 17088
rect 4065 17085 4077 17088
rect 4111 17116 4123 17119
rect 4430 17116 4436 17128
rect 4111 17088 4436 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 5460 17125 5488 17156
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7006 17184 7012 17196
rect 6963 17156 7012 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 8478 17184 8484 17196
rect 7432 17156 8484 17184
rect 7432 17144 7438 17156
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 8772 17193 8800 17224
rect 10597 17221 10609 17224
rect 10643 17252 10655 17255
rect 11606 17252 11612 17264
rect 10643 17224 11612 17252
rect 10643 17221 10655 17224
rect 10597 17215 10655 17221
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 9674 17184 9680 17196
rect 8803 17156 9680 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 9674 17144 9680 17156
rect 9732 17184 9738 17196
rect 10870 17184 10876 17196
rect 9732 17156 10876 17184
rect 9732 17144 9738 17156
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17085 5503 17119
rect 5445 17079 5503 17085
rect 5718 17076 5724 17128
rect 5776 17116 5782 17128
rect 5776 17088 5821 17116
rect 5776 17076 5782 17088
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 10980 17125 11008 17224
rect 11606 17212 11612 17224
rect 11664 17252 11670 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11664 17224 11805 17252
rect 11664 17212 11670 17224
rect 11793 17221 11805 17224
rect 11839 17252 11851 17255
rect 12618 17252 12624 17264
rect 11839 17224 12624 17252
rect 11839 17221 11851 17224
rect 11793 17215 11851 17221
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 13354 17212 13360 17264
rect 13412 17252 13418 17264
rect 14660 17252 14688 17292
rect 16761 17289 16773 17292
rect 16807 17289 16819 17323
rect 16761 17283 16819 17289
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 17494 17320 17500 17332
rect 16991 17292 17500 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 18690 17280 18696 17332
rect 18748 17320 18754 17332
rect 19058 17320 19064 17332
rect 18748 17292 19064 17320
rect 18748 17280 18754 17292
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 19429 17323 19487 17329
rect 19429 17320 19441 17323
rect 19392 17292 19441 17320
rect 19392 17280 19398 17292
rect 19429 17289 19441 17292
rect 19475 17289 19487 17323
rect 21358 17320 21364 17332
rect 21319 17292 21364 17320
rect 19429 17283 19487 17289
rect 13412 17224 14688 17252
rect 13412 17212 13418 17224
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 13633 17187 13691 17193
rect 11296 17156 13353 17184
rect 11296 17144 11302 17156
rect 10965 17119 11023 17125
rect 7892 17088 8242 17116
rect 7892 17076 7898 17088
rect 201 17051 259 17057
rect 201 17017 213 17051
rect 247 17048 259 17051
rect 3329 17051 3387 17057
rect 3329 17048 3341 17051
rect 247 17020 3341 17048
rect 247 17017 259 17020
rect 201 17011 259 17017
rect 3329 17017 3341 17020
rect 3375 17017 3387 17051
rect 4338 17048 4344 17060
rect 4299 17020 4344 17048
rect 3329 17011 3387 17017
rect 4338 17008 4344 17020
rect 4396 17008 4402 17060
rect 4709 17051 4767 17057
rect 4709 17017 4721 17051
rect 4755 17048 4767 17051
rect 4890 17048 4896 17060
rect 4755 17020 4896 17048
rect 4755 17017 4767 17020
rect 4709 17011 4767 17017
rect 4890 17008 4896 17020
rect 4948 17008 4954 17060
rect 5258 17008 5264 17060
rect 5316 17048 5322 17060
rect 5902 17048 5908 17060
rect 5316 17020 5666 17048
rect 5863 17020 5908 17048
rect 5316 17008 5322 17020
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 4430 16980 4436 16992
rect 4391 16952 4436 16980
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 5442 16980 5448 16992
rect 5224 16952 5448 16980
rect 5224 16940 5230 16952
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 5638 16980 5666 17020
rect 5902 17008 5908 17020
rect 5960 17008 5966 17060
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 8214 17048 8242 17088
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17085 11391 17119
rect 11333 17079 11391 17085
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17116 11575 17119
rect 11790 17116 11796 17128
rect 11563 17088 11796 17116
rect 11563 17085 11575 17088
rect 11517 17079 11575 17085
rect 8478 17048 8484 17060
rect 7064 17020 7109 17048
rect 8214 17020 8484 17048
rect 7064 17008 7070 17020
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 8573 17051 8631 17057
rect 8573 17017 8585 17051
rect 8619 17017 8631 17051
rect 11348 17048 11376 17079
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12176 17088 12449 17116
rect 11606 17048 11612 17060
rect 11348 17020 11612 17048
rect 8573 17011 8631 17017
rect 6181 16983 6239 16989
rect 6181 16980 6193 16983
rect 5638 16952 6193 16980
rect 6181 16949 6193 16952
rect 6227 16980 6239 16983
rect 6822 16980 6828 16992
rect 6227 16952 6828 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7190 16940 7196 16992
rect 7248 16980 7254 16992
rect 7837 16983 7895 16989
rect 7837 16980 7849 16983
rect 7248 16952 7849 16980
rect 7248 16940 7254 16952
rect 7837 16949 7849 16952
rect 7883 16949 7895 16983
rect 8294 16980 8300 16992
rect 8255 16952 8300 16980
rect 7837 16943 7895 16949
rect 8294 16940 8300 16952
rect 8352 16980 8358 16992
rect 8588 16980 8616 17011
rect 11606 17008 11612 17020
rect 11664 17008 11670 17060
rect 8352 16952 8616 16980
rect 9953 16983 10011 16989
rect 8352 16940 8358 16952
rect 9953 16949 9965 16983
rect 9999 16980 10011 16983
rect 11054 16980 11060 16992
rect 9999 16952 11060 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 11054 16940 11060 16952
rect 11112 16980 11118 16992
rect 12176 16989 12204 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12768 17088 12909 17116
rect 12768 17076 12774 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 13325 17116 13353 17156
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 13679 17156 15485 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 15473 17153 15485 17156
rect 15519 17184 15531 17187
rect 15838 17184 15844 17196
rect 15519 17156 15844 17184
rect 15519 17153 15531 17156
rect 15473 17147 15531 17153
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13325 17088 13737 17116
rect 12897 17079 12955 17085
rect 13725 17085 13737 17088
rect 13771 17116 13783 17119
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13771 17088 14013 17116
rect 13771 17085 13783 17088
rect 13725 17079 13783 17085
rect 14001 17085 14013 17088
rect 14047 17085 14059 17119
rect 14458 17116 14464 17128
rect 14419 17088 14464 17116
rect 14001 17079 14059 17085
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 15580 17125 15608 17156
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 15930 17144 15936 17196
rect 15988 17184 15994 17196
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 15988 17156 18061 17184
rect 15988 17144 15994 17156
rect 18049 17153 18061 17156
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17085 15623 17119
rect 16022 17116 16028 17128
rect 15983 17088 16028 17116
rect 15565 17079 15623 17085
rect 16022 17076 16028 17088
rect 16080 17116 16086 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 16080 17088 17233 17116
rect 16080 17076 16086 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17828 17088 18153 17116
rect 17828 17076 17834 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 19444 17116 19472 17283
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 21450 17280 21456 17332
rect 21508 17320 21514 17332
rect 21729 17323 21787 17329
rect 21729 17320 21741 17323
rect 21508 17292 21741 17320
rect 21508 17280 21514 17292
rect 21729 17289 21741 17292
rect 21775 17289 21787 17323
rect 21729 17283 21787 17289
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19444 17088 19717 17116
rect 18141 17079 18199 17085
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 20254 17076 20260 17128
rect 20312 17116 20318 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20312 17088 21189 17116
rect 20312 17076 20318 17088
rect 21177 17085 21189 17088
rect 21223 17116 21235 17119
rect 22097 17119 22155 17125
rect 22097 17116 22109 17119
rect 21223 17088 22109 17116
rect 21223 17085 21235 17088
rect 21177 17079 21235 17085
rect 22097 17085 22109 17088
rect 22143 17085 22155 17119
rect 22097 17079 22155 17085
rect 13170 17048 13176 17060
rect 13131 17020 13176 17048
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 15105 17051 15163 17057
rect 15105 17048 15117 17051
rect 13596 17020 15117 17048
rect 13596 17008 13602 17020
rect 15105 17017 15117 17020
rect 15151 17048 15163 17051
rect 15470 17048 15476 17060
rect 15151 17020 15476 17048
rect 15151 17017 15163 17020
rect 15105 17011 15163 17017
rect 15470 17008 15476 17020
rect 15528 17048 15534 17060
rect 15930 17048 15936 17060
rect 15528 17020 15936 17048
rect 15528 17008 15534 17020
rect 15930 17008 15936 17020
rect 15988 17008 15994 17060
rect 16298 17048 16304 17060
rect 16259 17020 16304 17048
rect 16298 17008 16304 17020
rect 16356 17008 16362 17060
rect 16761 17051 16819 17057
rect 16761 17017 16773 17051
rect 16807 17048 16819 17051
rect 18690 17048 18696 17060
rect 16807 17020 18696 17048
rect 16807 17017 16819 17020
rect 16761 17011 16819 17017
rect 18690 17008 18696 17020
rect 18748 17048 18754 17060
rect 19613 17051 19671 17057
rect 19613 17048 19625 17051
rect 18748 17020 19625 17048
rect 18748 17008 18754 17020
rect 19613 17017 19625 17020
rect 19659 17017 19671 17051
rect 19613 17011 19671 17017
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11112 16952 12173 16980
rect 11112 16940 11118 16952
rect 12161 16949 12173 16952
rect 12207 16980 12219 16983
rect 13633 16983 13691 16989
rect 13633 16980 13645 16983
rect 12207 16952 13645 16980
rect 12207 16949 12219 16952
rect 12161 16943 12219 16949
rect 13633 16949 13645 16952
rect 13679 16949 13691 16983
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 13633 16943 13691 16949
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15378 16980 15384 16992
rect 15068 16952 15384 16980
rect 15068 16940 15074 16952
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 20806 16980 20812 16992
rect 19576 16952 20812 16980
rect 19576 16940 19582 16952
rect 20806 16940 20812 16952
rect 20864 16980 20870 16992
rect 20901 16983 20959 16989
rect 20901 16980 20913 16983
rect 20864 16952 20913 16980
rect 20864 16940 20870 16952
rect 20901 16949 20913 16952
rect 20947 16949 20959 16983
rect 20901 16943 20959 16949
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 658 16776 664 16788
rect 619 16748 664 16776
rect 658 16736 664 16748
rect 716 16736 722 16788
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2406 16776 2412 16788
rect 2367 16748 2412 16776
rect 2406 16736 2412 16748
rect 2464 16776 2470 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 2464 16748 2697 16776
rect 2464 16736 2470 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 2685 16739 2743 16745
rect 3697 16779 3755 16785
rect 3697 16745 3709 16779
rect 3743 16776 3755 16779
rect 3970 16776 3976 16788
rect 3743 16748 3976 16776
rect 3743 16745 3755 16748
rect 3697 16739 3755 16745
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 4126 16748 9413 16776
rect 937 16711 995 16717
rect 937 16677 949 16711
rect 983 16708 995 16711
rect 4126 16708 4154 16748
rect 9401 16745 9413 16748
rect 9447 16745 9459 16779
rect 10318 16776 10324 16788
rect 9401 16739 9459 16745
rect 9743 16748 10324 16776
rect 983 16680 4154 16708
rect 5623 16711 5681 16717
rect 983 16677 995 16680
rect 937 16671 995 16677
rect 5623 16677 5635 16711
rect 5669 16708 5681 16711
rect 6086 16708 6092 16720
rect 5669 16680 6092 16708
rect 5669 16677 5681 16680
rect 5623 16671 5681 16677
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 7282 16708 7288 16720
rect 6972 16680 7288 16708
rect 6972 16668 6978 16680
rect 7282 16668 7288 16680
rect 7340 16708 7346 16720
rect 7469 16711 7527 16717
rect 7469 16708 7481 16711
rect 7340 16680 7481 16708
rect 7340 16668 7346 16680
rect 7469 16677 7481 16680
rect 7515 16677 7527 16711
rect 7469 16671 7527 16677
rect 7834 16668 7840 16720
rect 7892 16708 7898 16720
rect 8110 16708 8116 16720
rect 7892 16680 8116 16708
rect 7892 16668 7898 16680
rect 8110 16668 8116 16680
rect 8168 16708 8174 16720
rect 8205 16711 8263 16717
rect 8205 16708 8217 16711
rect 8168 16680 8217 16708
rect 8168 16668 8174 16680
rect 8205 16677 8217 16680
rect 8251 16677 8263 16711
rect 8205 16671 8263 16677
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 8757 16711 8815 16717
rect 8757 16708 8769 16711
rect 8628 16680 8769 16708
rect 8628 16668 8634 16680
rect 8757 16677 8769 16680
rect 8803 16677 8815 16711
rect 8757 16671 8815 16677
rect 8938 16668 8944 16720
rect 8996 16708 9002 16720
rect 9743 16708 9771 16748
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 11333 16779 11391 16785
rect 11333 16776 11345 16779
rect 10928 16748 11345 16776
rect 10928 16736 10934 16748
rect 11333 16745 11345 16748
rect 11379 16745 11391 16779
rect 11333 16739 11391 16745
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 12710 16776 12716 16788
rect 12575 16748 12716 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 12710 16736 12716 16748
rect 12768 16776 12774 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 12768 16748 14105 16776
rect 12768 16736 12774 16748
rect 14093 16745 14105 16748
rect 14139 16776 14151 16779
rect 14458 16776 14464 16788
rect 14139 16748 14464 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 15102 16776 15108 16788
rect 15063 16748 15108 16776
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 15378 16736 15384 16788
rect 15436 16776 15442 16788
rect 16945 16779 17003 16785
rect 16945 16776 16957 16779
rect 15436 16748 16957 16776
rect 15436 16736 15442 16748
rect 16945 16745 16957 16748
rect 16991 16745 17003 16779
rect 18322 16776 18328 16788
rect 18283 16748 18328 16776
rect 16945 16739 17003 16745
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 18874 16776 18880 16788
rect 18835 16748 18880 16776
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 9858 16708 9864 16720
rect 8996 16680 9771 16708
rect 9819 16680 9864 16708
rect 8996 16668 9002 16680
rect 9858 16668 9864 16680
rect 9916 16668 9922 16720
rect 11716 16680 13308 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2130 16640 2136 16652
rect 1443 16612 2136 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 3028 16643 3086 16649
rect 3028 16609 3040 16643
rect 3074 16640 3086 16643
rect 3326 16640 3332 16652
rect 3074 16612 3332 16640
rect 3074 16609 3086 16612
rect 3028 16603 3086 16609
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 4316 16643 4374 16649
rect 4316 16609 4328 16643
rect 4362 16640 4374 16643
rect 4522 16640 4528 16652
rect 4362 16612 4528 16640
rect 4362 16609 4374 16612
rect 4316 16603 4374 16609
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5350 16640 5356 16652
rect 5307 16612 5356 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 6454 16640 6460 16652
rect 5500 16612 6460 16640
rect 5500 16600 5506 16612
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11422 16640 11428 16652
rect 11204 16612 11428 16640
rect 11204 16600 11210 16612
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 11716 16649 11744 16680
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 11664 16612 11713 16640
rect 11664 16600 11670 16612
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 12802 16640 12808 16652
rect 12763 16612 12808 16640
rect 11701 16603 11759 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13280 16649 13308 16680
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 16669 16711 16727 16717
rect 16669 16708 16681 16711
rect 13964 16680 16681 16708
rect 13964 16668 13970 16680
rect 16669 16677 16681 16680
rect 16715 16677 16727 16711
rect 16669 16671 16727 16677
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 19429 16711 19487 16717
rect 19429 16708 19441 16711
rect 17920 16680 19441 16708
rect 17920 16668 17926 16680
rect 19429 16677 19441 16680
rect 19475 16677 19487 16711
rect 19429 16671 19487 16677
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 21085 16711 21143 16717
rect 21085 16708 21097 16711
rect 20772 16680 21097 16708
rect 20772 16668 20778 16680
rect 21085 16677 21097 16680
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 15562 16640 15568 16652
rect 15523 16612 15568 16640
rect 13265 16603 13323 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 16022 16640 16028 16652
rect 15795 16612 16028 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 17276 16612 17325 16640
rect 17276 16600 17282 16612
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16609 18475 16643
rect 18690 16640 18696 16652
rect 18651 16612 18696 16640
rect 18417 16603 18475 16609
rect 385 16575 443 16581
rect 385 16541 397 16575
rect 431 16572 443 16575
rect 2222 16572 2228 16584
rect 431 16544 2228 16572
rect 431 16541 443 16544
rect 385 16535 443 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 6822 16572 6828 16584
rect 4310 16544 6828 16572
rect 3099 16507 3157 16513
rect 3099 16473 3111 16507
rect 3145 16504 3157 16507
rect 4310 16504 4338 16544
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16572 7067 16575
rect 7466 16572 7472 16584
rect 7055 16544 7472 16572
rect 7055 16541 7067 16544
rect 7009 16535 7067 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 9306 16572 9312 16584
rect 8159 16544 9312 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 3145 16476 4338 16504
rect 4387 16507 4445 16513
rect 3145 16473 3157 16476
rect 3099 16467 3157 16473
rect 4387 16473 4399 16507
rect 4433 16504 4445 16507
rect 8128 16504 8156 16535
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 9766 16572 9772 16584
rect 9727 16544 9772 16572
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 12618 16572 12624 16584
rect 10459 16544 12624 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 4433 16476 8156 16504
rect 4433 16473 4445 16476
rect 4387 16467 4445 16473
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 9214 16504 9220 16516
rect 8536 16476 9220 16504
rect 8536 16464 8542 16476
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10428 16504 10456 16535
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 13538 16572 13544 16584
rect 13499 16544 13544 16572
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 14516 16544 15853 16572
rect 14516 16532 14522 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 18432 16572 18460 16603
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 19426 16572 19432 16584
rect 16448 16544 19432 16572
rect 16448 16532 16454 16544
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20864 16544 21005 16572
rect 20864 16532 20870 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 21266 16572 21272 16584
rect 21227 16544 21272 16572
rect 20993 16535 21051 16541
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 9640 16476 10456 16504
rect 9640 16464 9646 16476
rect 11146 16464 11152 16516
rect 11204 16504 11210 16516
rect 14369 16507 14427 16513
rect 14369 16504 14381 16507
rect 11204 16476 14381 16504
rect 11204 16464 11210 16476
rect 14369 16473 14381 16476
rect 14415 16473 14427 16507
rect 14369 16467 14427 16473
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 17865 16507 17923 16513
rect 17865 16504 17877 16507
rect 14884 16476 17877 16504
rect 14884 16464 14890 16476
rect 17865 16473 17877 16476
rect 17911 16504 17923 16507
rect 18509 16507 18567 16513
rect 18509 16504 18521 16507
rect 17911 16476 18521 16504
rect 17911 16473 17923 16476
rect 17865 16467 17923 16473
rect 18509 16473 18521 16476
rect 18555 16473 18567 16507
rect 18509 16467 18567 16473
rect 4154 16396 4160 16448
rect 4212 16436 4218 16448
rect 4709 16439 4767 16445
rect 4709 16436 4721 16439
rect 4212 16408 4721 16436
rect 4212 16396 4218 16408
rect 4709 16405 4721 16408
rect 4755 16405 4767 16439
rect 4709 16399 4767 16405
rect 5169 16439 5227 16445
rect 5169 16405 5181 16439
rect 5215 16436 5227 16439
rect 5718 16436 5724 16448
rect 5215 16408 5724 16436
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 6178 16436 6184 16448
rect 6139 16408 6184 16436
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 6917 16439 6975 16445
rect 6917 16405 6929 16439
rect 6963 16436 6975 16439
rect 7006 16436 7012 16448
rect 6963 16408 7012 16436
rect 6963 16405 6975 16408
rect 6917 16399 6975 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 7708 16408 7849 16436
rect 7708 16396 7714 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 8754 16396 8760 16448
rect 8812 16436 8818 16448
rect 9030 16436 9036 16448
rect 8812 16408 9036 16436
rect 8812 16396 8818 16408
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9306 16436 9312 16448
rect 9171 16408 9312 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 10686 16436 10692 16448
rect 10647 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16436 10750 16448
rect 11057 16439 11115 16445
rect 11057 16436 11069 16439
rect 10744 16408 11069 16436
rect 10744 16396 10750 16408
rect 11057 16405 11069 16408
rect 11103 16405 11115 16439
rect 11057 16399 11115 16405
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 13906 16436 13912 16448
rect 12676 16408 13912 16436
rect 12676 16396 12682 16408
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 15160 16408 16405 16436
rect 15160 16396 15166 16408
rect 16393 16405 16405 16408
rect 16439 16436 16451 16439
rect 17586 16436 17592 16448
rect 16439 16408 17592 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 17586 16396 17592 16408
rect 17644 16436 17650 16448
rect 17770 16436 17776 16448
rect 17644 16408 17776 16436
rect 17644 16396 17650 16408
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 2041 16235 2099 16241
rect 2041 16201 2053 16235
rect 2087 16232 2099 16235
rect 2130 16232 2136 16244
rect 2087 16204 2136 16232
rect 2087 16201 2099 16204
rect 2041 16195 2099 16201
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 3326 16232 3332 16244
rect 2547 16204 3332 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 3326 16192 3332 16204
rect 3384 16232 3390 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 3384 16204 3433 16232
rect 3384 16192 3390 16204
rect 3421 16201 3433 16204
rect 3467 16201 3479 16235
rect 3421 16195 3479 16201
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 3694 16232 3700 16244
rect 3559 16204 3700 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 3694 16192 3700 16204
rect 3752 16232 3758 16244
rect 3752 16204 4267 16232
rect 3752 16192 3758 16204
rect 106 16124 112 16176
rect 164 16164 170 16176
rect 1581 16167 1639 16173
rect 1581 16164 1593 16167
rect 164 16136 1593 16164
rect 164 16124 170 16136
rect 1581 16133 1593 16136
rect 1627 16133 1639 16167
rect 1581 16127 1639 16133
rect 3602 16124 3608 16176
rect 3660 16164 3666 16176
rect 4154 16164 4160 16176
rect 3660 16136 4160 16164
rect 3660 16124 3666 16136
rect 4154 16124 4160 16136
rect 4212 16164 4218 16176
rect 4239 16164 4267 16204
rect 4430 16192 4436 16244
rect 4488 16232 4494 16244
rect 4522 16232 4528 16244
rect 4488 16204 4528 16232
rect 4488 16192 4494 16204
rect 4522 16192 4528 16204
rect 4580 16232 4586 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 4580 16204 5181 16232
rect 4580 16192 4586 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6052 16204 6193 16232
rect 6052 16192 6058 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 6181 16195 6239 16201
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 6656 16204 10456 16232
rect 4295 16167 4353 16173
rect 4295 16164 4307 16167
rect 4212 16136 4307 16164
rect 4212 16124 4218 16136
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 4239 16096 4267 16136
rect 4295 16133 4307 16136
rect 4341 16133 4353 16167
rect 4295 16127 4353 16133
rect 4801 16167 4859 16173
rect 4801 16133 4813 16167
rect 4847 16164 4859 16167
rect 6656 16164 6684 16204
rect 4847 16136 6684 16164
rect 4847 16133 4859 16136
rect 4801 16127 4859 16133
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 8386 16164 8392 16176
rect 6880 16136 8392 16164
rect 6880 16124 6886 16136
rect 7944 16105 7972 16136
rect 8386 16124 8392 16136
rect 8444 16124 8450 16176
rect 8481 16167 8539 16173
rect 8481 16133 8493 16167
rect 8527 16164 8539 16167
rect 8754 16164 8760 16176
rect 8527 16136 8760 16164
rect 8527 16133 8539 16136
rect 8481 16127 8539 16133
rect 8754 16124 8760 16136
rect 8812 16164 8818 16176
rect 9950 16164 9956 16176
rect 8812 16136 9956 16164
rect 8812 16124 8818 16136
rect 4525 16099 4583 16105
rect 4525 16096 4537 16099
rect 2731 16068 4200 16096
rect 4239 16068 4537 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 106 15988 112 16040
rect 164 16028 170 16040
rect 845 16031 903 16037
rect 845 16028 857 16031
rect 164 16000 857 16028
rect 164 15988 170 16000
rect 845 15997 857 16000
rect 891 15997 903 16031
rect 845 15991 903 15997
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1762 16028 1768 16040
rect 1443 16000 1768 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 4172 16028 4200 16068
rect 4525 16065 4537 16068
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 8202 16056 8208 16108
rect 8260 16096 8266 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 8260 16068 9229 16096
rect 8260 16056 8266 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 4614 16028 4620 16040
rect 4172 16000 4620 16028
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 6086 15988 6092 16040
rect 6144 15988 6150 16040
rect 661 15963 719 15969
rect 661 15929 673 15963
rect 707 15960 719 15963
rect 2774 15960 2780 15972
rect 707 15932 2589 15960
rect 2735 15932 2780 15960
rect 707 15929 719 15932
rect 661 15923 719 15929
rect 2561 15892 2589 15932
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 3326 15960 3332 15972
rect 3287 15932 3332 15960
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 4154 15920 4160 15972
rect 4212 15960 4218 15972
rect 6104 15960 6132 15988
rect 4212 15932 4257 15960
rect 5552 15932 6132 15960
rect 4212 15920 4218 15932
rect 3513 15895 3571 15901
rect 3513 15892 3525 15895
rect 2561 15864 3525 15892
rect 3513 15861 3525 15864
rect 3559 15892 3571 15895
rect 3605 15895 3663 15901
rect 3605 15892 3617 15895
rect 3559 15864 3617 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 3605 15861 3617 15864
rect 3651 15861 3663 15895
rect 3605 15855 3663 15861
rect 3694 15852 3700 15904
rect 3752 15892 3758 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3752 15864 3985 15892
rect 3752 15852 3758 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 3973 15855 4031 15861
rect 5074 15852 5080 15904
rect 5132 15892 5138 15904
rect 5552 15901 5580 15932
rect 6362 15920 6368 15972
rect 6420 15960 6426 15972
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 6420 15932 7665 15960
rect 6420 15920 6426 15932
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 7653 15923 7711 15929
rect 8030 15963 8088 15969
rect 8030 15929 8042 15963
rect 8076 15960 8088 15963
rect 8110 15960 8116 15972
rect 8076 15932 8116 15960
rect 8076 15929 8088 15932
rect 8030 15923 8088 15929
rect 5537 15895 5595 15901
rect 5537 15892 5549 15895
rect 5132 15864 5549 15892
rect 5132 15852 5138 15864
rect 5537 15861 5549 15864
rect 5583 15861 5595 15895
rect 5537 15855 5595 15861
rect 5721 15895 5779 15901
rect 5721 15861 5733 15895
rect 5767 15892 5779 15895
rect 6086 15892 6092 15904
rect 5767 15864 6092 15892
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 6825 15895 6883 15901
rect 6825 15861 6837 15895
rect 6871 15892 6883 15895
rect 6914 15892 6920 15904
rect 6871 15864 6920 15892
rect 6871 15861 6883 15864
rect 6825 15855 6883 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 7282 15892 7288 15904
rect 7064 15864 7288 15892
rect 7064 15852 7070 15864
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7668 15892 7696 15923
rect 8110 15920 8116 15932
rect 8168 15960 8174 15972
rect 8849 15963 8907 15969
rect 8849 15960 8861 15963
rect 8168 15932 8861 15960
rect 8168 15920 8174 15932
rect 8849 15929 8861 15932
rect 8895 15929 8907 15963
rect 9122 15960 9128 15972
rect 8849 15923 8907 15929
rect 8956 15932 9128 15960
rect 7834 15892 7840 15904
rect 7668 15864 7840 15892
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8956 15892 8984 15932
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 8444 15864 8984 15892
rect 9232 15892 9260 16059
rect 9324 15960 9352 16136
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 10428 16164 10456 16204
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 11103 16235 11161 16241
rect 11103 16232 11115 16235
rect 10836 16204 11115 16232
rect 10836 16192 10842 16204
rect 11103 16201 11115 16204
rect 11149 16201 11161 16235
rect 11103 16195 11161 16201
rect 11238 16192 11244 16244
rect 11296 16232 11302 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11296 16204 12173 16232
rect 11296 16192 11302 16204
rect 10686 16164 10692 16176
rect 10428 16136 10692 16164
rect 10686 16124 10692 16136
rect 10744 16164 10750 16176
rect 10873 16167 10931 16173
rect 10873 16164 10885 16167
rect 10744 16136 10885 16164
rect 10744 16124 10750 16136
rect 10873 16133 10885 16136
rect 10919 16164 10931 16167
rect 11606 16164 11612 16176
rect 10919 16136 11612 16164
rect 10919 16133 10931 16136
rect 10873 16127 10931 16133
rect 11606 16124 11612 16136
rect 11664 16164 11670 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 11664 16136 11805 16164
rect 11664 16124 11670 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 11992 16164 12020 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15562 16232 15568 16244
rect 15427 16204 15568 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15197 16167 15255 16173
rect 15197 16164 15209 16167
rect 11992 16136 15209 16164
rect 9490 16056 9496 16108
rect 9548 16096 9554 16108
rect 9858 16096 9864 16108
rect 9548 16068 9864 16096
rect 9548 16056 9554 16068
rect 9858 16056 9864 16068
rect 9916 16096 9922 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 9916 16068 10425 16096
rect 9916 16056 9922 16068
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 11422 16096 11428 16108
rect 11383 16068 11428 16096
rect 10413 16059 10471 16065
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10502 16028 10508 16040
rect 10183 16000 10508 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10502 15988 10508 16000
rect 10560 16028 10566 16040
rect 11032 16031 11090 16037
rect 11032 16028 11044 16031
rect 10560 16000 11044 16028
rect 10560 15988 10566 16000
rect 11032 15997 11044 16000
rect 11078 16028 11090 16031
rect 11146 16028 11152 16040
rect 11078 16000 11152 16028
rect 11078 15997 11090 16000
rect 11032 15991 11090 15997
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 11992 16028 12020 16136
rect 15197 16133 15209 16136
rect 15243 16133 15255 16167
rect 15197 16127 15255 16133
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12124 16068 12940 16096
rect 12124 16056 12130 16068
rect 12912 16040 12940 16068
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13044 16068 13578 16096
rect 13044 16056 13050 16068
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 11992 16000 12449 16028
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12894 16028 12900 16040
rect 12855 16000 12900 16028
rect 12437 15991 12495 15997
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 13550 16028 13578 16068
rect 13786 16068 13921 16096
rect 13786 16028 13814 16068
rect 13909 16065 13921 16068
rect 13955 16096 13967 16099
rect 15396 16096 15424 16195
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 17218 16232 17224 16244
rect 16080 16204 17224 16232
rect 16080 16192 16086 16204
rect 17218 16192 17224 16204
rect 17276 16232 17282 16244
rect 17494 16232 17500 16244
rect 17276 16204 17500 16232
rect 17276 16192 17282 16204
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 18748 16204 19073 16232
rect 18748 16192 18754 16204
rect 19061 16201 19073 16204
rect 19107 16232 19119 16235
rect 20254 16232 20260 16244
rect 19107 16204 20260 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 15470 16124 15476 16176
rect 15528 16164 15534 16176
rect 18966 16164 18972 16176
rect 15528 16136 18972 16164
rect 15528 16124 15534 16136
rect 18966 16124 18972 16136
rect 19024 16124 19030 16176
rect 19150 16124 19156 16176
rect 19208 16164 19214 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 19208 16136 19441 16164
rect 19208 16124 19214 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 13955 16068 15424 16096
rect 15948 16068 16865 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 14292 16037 14320 16068
rect 15948 16040 15976 16068
rect 16853 16065 16865 16068
rect 16899 16096 16911 16099
rect 16942 16096 16948 16108
rect 16899 16068 16948 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 17736 16068 18552 16096
rect 17736 16056 17742 16068
rect 13550 16000 13814 16028
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 15102 16028 15108 16040
rect 14599 16000 15108 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 15930 16028 15936 16040
rect 15887 16000 15936 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 9493 15963 9551 15969
rect 9493 15960 9505 15963
rect 9324 15932 9505 15960
rect 9493 15929 9505 15932
rect 9539 15929 9551 15963
rect 9493 15923 9551 15929
rect 9585 15963 9643 15969
rect 9585 15929 9597 15963
rect 9631 15929 9643 15963
rect 9585 15923 9643 15929
rect 9600 15892 9628 15923
rect 11514 15920 11520 15972
rect 11572 15960 11578 15972
rect 15120 15960 15148 15988
rect 15562 15960 15568 15972
rect 11572 15932 14044 15960
rect 15120 15932 15568 15960
rect 11572 15920 11578 15932
rect 9232 15864 9628 15892
rect 8444 15852 8450 15864
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 11054 15892 11060 15904
rect 10744 15864 11060 15892
rect 10744 15852 10750 15864
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12710 15892 12716 15904
rect 12671 15864 12716 15892
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13170 15892 13176 15904
rect 12860 15864 13176 15892
rect 12860 15852 12866 15864
rect 13170 15852 13176 15864
rect 13228 15892 13234 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13228 15864 13461 15892
rect 13228 15852 13234 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 14016 15892 14044 15932
rect 15562 15920 15568 15932
rect 15620 15960 15626 15972
rect 16040 15960 16068 15991
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 18524 16037 18552 16068
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 16724 16000 17877 16028
rect 16724 15988 16730 16000
rect 17865 15997 17877 16000
rect 17911 16028 17923 16031
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17911 16000 18061 16028
rect 17911 15997 17923 16000
rect 17865 15991 17923 15997
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18509 16031 18567 16037
rect 18509 15997 18521 16031
rect 18555 16028 18567 16031
rect 18690 16028 18696 16040
rect 18555 16000 18696 16028
rect 18555 15997 18567 16000
rect 18509 15991 18567 15997
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 19444 16028 19472 16127
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 20772 16068 22017 16096
rect 20772 16056 20778 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 19444 16000 19717 16028
rect 19705 15997 19717 16000
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 19794 15988 19800 16040
rect 19852 16028 19858 16040
rect 21228 16031 21286 16037
rect 21228 16028 21240 16031
rect 19852 16000 21240 16028
rect 19852 15988 19858 16000
rect 21228 15997 21240 16000
rect 21274 15997 21286 16031
rect 21228 15991 21286 15997
rect 21315 16031 21373 16037
rect 21315 15997 21327 16031
rect 21361 16028 21373 16031
rect 21634 16028 21640 16040
rect 21361 16000 21640 16028
rect 21361 15997 21373 16000
rect 21315 15991 21373 15997
rect 15620 15932 16068 15960
rect 16301 15963 16359 15969
rect 15620 15920 15626 15932
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 16390 15960 16396 15972
rect 16347 15932 16396 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 18230 15960 18236 15972
rect 17052 15932 18236 15960
rect 14093 15895 14151 15901
rect 14093 15892 14105 15895
rect 14016 15864 14105 15892
rect 13449 15855 13507 15861
rect 14093 15861 14105 15864
rect 14139 15861 14151 15895
rect 14093 15855 14151 15861
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 17052 15892 17080 15932
rect 18230 15920 18236 15932
rect 18288 15920 18294 15972
rect 18785 15963 18843 15969
rect 18785 15929 18797 15963
rect 18831 15960 18843 15963
rect 18966 15960 18972 15972
rect 18831 15932 18972 15960
rect 18831 15929 18843 15932
rect 18785 15923 18843 15929
rect 18966 15920 18972 15932
rect 19024 15920 19030 15972
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 19613 15963 19671 15969
rect 19613 15960 19625 15963
rect 19392 15932 19625 15960
rect 19392 15920 19398 15932
rect 19613 15929 19625 15932
rect 19659 15929 19671 15963
rect 21243 15960 21271 15991
rect 21634 15988 21640 16000
rect 21692 15988 21698 16040
rect 21243 15932 21496 15960
rect 19613 15923 19671 15929
rect 21468 15904 21496 15932
rect 15243 15864 17080 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 19702 15852 19708 15904
rect 19760 15892 19766 15904
rect 20806 15892 20812 15904
rect 19760 15864 20812 15892
rect 19760 15852 19766 15864
rect 20806 15852 20812 15864
rect 20864 15892 20870 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20864 15864 20913 15892
rect 20864 15852 20870 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 21450 15852 21456 15904
rect 21508 15892 21514 15904
rect 21637 15895 21695 15901
rect 21637 15892 21649 15895
rect 21508 15864 21649 15892
rect 21508 15852 21514 15864
rect 21637 15861 21649 15864
rect 21683 15861 21695 15895
rect 21637 15855 21695 15861
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 1762 15688 1768 15700
rect 1719 15660 1768 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2832 15660 3249 15688
rect 2832 15648 2838 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 4614 15688 4620 15700
rect 4575 15660 4620 15688
rect 3237 15651 3295 15657
rect 845 15623 903 15629
rect 845 15589 857 15623
rect 891 15620 903 15623
rect 2314 15620 2320 15632
rect 891 15592 2320 15620
rect 891 15589 903 15592
rect 845 15583 903 15589
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 2409 15623 2467 15629
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 2590 15620 2596 15632
rect 2455 15592 2596 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 2958 15620 2964 15632
rect 2919 15592 2964 15620
rect 2958 15580 2964 15592
rect 3016 15580 3022 15632
rect 3252 15620 3280 15651
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5350 15688 5356 15700
rect 5311 15660 5356 15688
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5445 15691 5503 15697
rect 5445 15657 5457 15691
rect 5491 15688 5503 15691
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 5491 15660 8953 15688
rect 5491 15657 5503 15660
rect 5445 15651 5503 15657
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 13446 15688 13452 15700
rect 10008 15660 13452 15688
rect 10008 15648 10014 15660
rect 13446 15648 13452 15660
rect 13504 15688 13510 15700
rect 14921 15691 14979 15697
rect 14921 15688 14933 15691
rect 13504 15660 14933 15688
rect 13504 15648 13510 15660
rect 14921 15657 14933 15660
rect 14967 15657 14979 15691
rect 14921 15651 14979 15657
rect 15105 15691 15163 15697
rect 15105 15657 15117 15691
rect 15151 15688 15163 15691
rect 16022 15688 16028 15700
rect 15151 15660 16028 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 18138 15688 18144 15700
rect 17144 15660 18144 15688
rect 3252 15592 4522 15620
rect 1118 15512 1124 15564
rect 1176 15552 1182 15564
rect 1762 15552 1768 15564
rect 1176 15524 1768 15552
rect 1176 15512 1182 15524
rect 1762 15512 1768 15524
rect 1820 15512 1826 15564
rect 3510 15512 3516 15564
rect 3568 15552 3574 15564
rect 3605 15555 3663 15561
rect 3605 15552 3617 15555
rect 3568 15524 3617 15552
rect 3568 15512 3574 15524
rect 3605 15521 3617 15524
rect 3651 15521 3663 15555
rect 3605 15515 3663 15521
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4376 15555 4434 15561
rect 4376 15552 4388 15555
rect 4304 15524 4388 15552
rect 4304 15512 4310 15524
rect 4376 15521 4388 15524
rect 4422 15521 4434 15555
rect 4494 15552 4522 15592
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 5166 15620 5172 15632
rect 4948 15592 5172 15620
rect 4948 15580 4954 15592
rect 5166 15580 5172 15592
rect 5224 15620 5230 15632
rect 5629 15623 5687 15629
rect 5629 15620 5641 15623
rect 5224 15592 5641 15620
rect 5224 15580 5230 15592
rect 5629 15589 5641 15592
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 5994 15580 6000 15632
rect 6052 15620 6058 15632
rect 6457 15623 6515 15629
rect 6457 15620 6469 15623
rect 6052 15592 6469 15620
rect 6052 15580 6058 15592
rect 6457 15589 6469 15592
rect 6503 15589 6515 15623
rect 6457 15583 6515 15589
rect 6638 15580 6644 15632
rect 6696 15620 6702 15632
rect 8113 15623 8171 15629
rect 8113 15620 8125 15623
rect 6696 15592 8125 15620
rect 6696 15580 6702 15592
rect 8113 15589 8125 15592
rect 8159 15620 8171 15623
rect 8386 15620 8392 15632
rect 8159 15592 8392 15620
rect 8159 15589 8171 15592
rect 8113 15583 8171 15589
rect 8386 15580 8392 15592
rect 8444 15580 8450 15632
rect 8478 15580 8484 15632
rect 8536 15620 8542 15632
rect 8665 15623 8723 15629
rect 8665 15620 8677 15623
rect 8536 15592 8677 15620
rect 8536 15580 8542 15592
rect 8665 15589 8677 15592
rect 8711 15620 8723 15623
rect 8754 15620 8760 15632
rect 8711 15592 8760 15620
rect 8711 15589 8723 15592
rect 8665 15583 8723 15589
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9858 15620 9864 15632
rect 9819 15592 9864 15620
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 10962 15580 10968 15632
rect 11020 15620 11026 15632
rect 11146 15620 11152 15632
rect 11020 15592 11152 15620
rect 11020 15580 11026 15592
rect 11146 15580 11152 15592
rect 11204 15620 11210 15632
rect 11425 15623 11483 15629
rect 11425 15620 11437 15623
rect 11204 15592 11437 15620
rect 11204 15580 11210 15592
rect 11425 15589 11437 15592
rect 11471 15589 11483 15623
rect 11425 15583 11483 15589
rect 11977 15623 12035 15629
rect 11977 15589 11989 15623
rect 12023 15620 12035 15623
rect 12618 15620 12624 15632
rect 12023 15592 12624 15620
rect 12023 15589 12035 15592
rect 11977 15583 12035 15589
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 13170 15620 13176 15632
rect 12820 15592 13176 15620
rect 6178 15552 6184 15564
rect 4494 15524 6184 15552
rect 4376 15515 4434 15521
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 12820 15561 12848 15592
rect 13170 15580 13176 15592
rect 13228 15620 13234 15632
rect 13464 15620 13492 15648
rect 13228 15592 13492 15620
rect 13228 15580 13234 15592
rect 14826 15580 14832 15632
rect 14884 15620 14890 15632
rect 17144 15620 17172 15660
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 19426 15688 19432 15700
rect 19387 15660 19432 15688
rect 19426 15648 19432 15660
rect 19484 15688 19490 15700
rect 19484 15660 20944 15688
rect 19484 15648 19490 15660
rect 19978 15620 19984 15632
rect 14884 15592 19984 15620
rect 14884 15580 14890 15592
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 12759 15524 12817 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12805 15521 12817 15524
rect 12851 15521 12863 15555
rect 12805 15515 12863 15521
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 12952 15524 13277 15552
rect 12952 15512 12958 15524
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 14642 15512 14648 15564
rect 14700 15552 14706 15564
rect 15102 15552 15108 15564
rect 14700 15524 15108 15552
rect 14700 15512 14706 15524
rect 15102 15512 15108 15524
rect 15160 15552 15166 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 15160 15524 15301 15552
rect 15160 15512 15166 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15562 15512 15568 15564
rect 15620 15552 15626 15564
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 15620 15524 15761 15552
rect 15620 15512 15626 15524
rect 15749 15521 15761 15524
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 17034 15512 17040 15564
rect 17092 15552 17098 15564
rect 17144 15561 17172 15592
rect 19978 15580 19984 15592
rect 20036 15580 20042 15632
rect 20916 15629 20944 15660
rect 20901 15623 20959 15629
rect 20901 15589 20913 15623
rect 20947 15589 20959 15623
rect 20901 15583 20959 15589
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 17092 15524 17141 15552
rect 17092 15512 17098 15524
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 17494 15552 17500 15564
rect 17451 15524 17500 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 17494 15512 17500 15524
rect 17552 15552 17558 15564
rect 17552 15524 18184 15552
rect 17552 15512 17558 15524
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 2314 15484 2320 15496
rect 1452 15456 2320 15484
rect 1452 15444 1458 15456
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3528 15484 3556 15512
rect 3016 15456 3556 15484
rect 3016 15444 3022 15456
rect 3878 15444 3884 15496
rect 3936 15484 3942 15496
rect 4154 15484 4160 15496
rect 3936 15456 4160 15484
rect 3936 15444 3942 15456
rect 4154 15444 4160 15456
rect 4212 15484 4218 15496
rect 4798 15484 4804 15496
rect 4212 15456 4804 15484
rect 4212 15444 4218 15456
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5040 15456 5457 15484
rect 5040 15444 5046 15456
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 6196 15484 6224 15512
rect 6546 15484 6552 15496
rect 6196 15456 6552 15484
rect 5445 15447 5503 15453
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 7653 15487 7711 15493
rect 7653 15484 7665 15487
rect 6696 15456 7665 15484
rect 6696 15444 6702 15456
rect 7653 15453 7665 15456
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7892 15456 8033 15484
rect 7892 15444 7898 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 8021 15447 8079 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15484 11391 15487
rect 11422 15484 11428 15496
rect 11379 15456 11428 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 12066 15484 12072 15496
rect 11762 15456 12072 15484
rect 750 15376 756 15428
rect 808 15416 814 15428
rect 1118 15416 1124 15428
rect 808 15388 1124 15416
rect 808 15376 814 15388
rect 1118 15376 1124 15388
rect 1176 15376 1182 15428
rect 3050 15376 3056 15428
rect 3108 15416 3114 15428
rect 6181 15419 6239 15425
rect 6181 15416 6193 15419
rect 3108 15388 6193 15416
rect 3108 15376 3114 15388
rect 6181 15385 6193 15388
rect 6227 15416 6239 15419
rect 6270 15416 6276 15428
rect 6227 15388 6276 15416
rect 6227 15385 6239 15388
rect 6181 15379 6239 15385
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 6917 15419 6975 15425
rect 6917 15385 6929 15419
rect 6963 15416 6975 15419
rect 10042 15416 10048 15428
rect 6963 15388 10048 15416
rect 6963 15385 6975 15388
rect 6917 15379 6975 15385
rect 2041 15351 2099 15357
rect 2041 15317 2053 15351
rect 2087 15348 2099 15351
rect 3234 15348 3240 15360
rect 2087 15320 3240 15348
rect 2087 15317 2099 15320
rect 2041 15311 2099 15317
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 3421 15351 3479 15357
rect 3421 15317 3433 15351
rect 3467 15348 3479 15351
rect 3694 15348 3700 15360
rect 3467 15320 3700 15348
rect 3467 15317 3479 15320
rect 3421 15311 3479 15317
rect 3694 15308 3700 15320
rect 3752 15308 3758 15360
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 4154 15348 4160 15360
rect 4028 15320 4160 15348
rect 4028 15308 4034 15320
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 5997 15351 6055 15357
rect 5997 15348 6009 15351
rect 5408 15320 6009 15348
rect 5408 15308 5414 15320
rect 5997 15317 6009 15320
rect 6043 15317 6055 15351
rect 5997 15311 6055 15317
rect 6546 15308 6552 15360
rect 6604 15348 6610 15360
rect 6932 15348 6960 15379
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 10318 15416 10324 15428
rect 10279 15388 10324 15416
rect 10318 15376 10324 15388
rect 10376 15376 10382 15428
rect 10781 15419 10839 15425
rect 10781 15385 10793 15419
rect 10827 15416 10839 15419
rect 11762 15416 11790 15456
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 13446 15484 13452 15496
rect 13407 15456 13452 15484
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15712 15456 15853 15484
rect 15712 15444 15718 15456
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 17586 15484 17592 15496
rect 17547 15456 17592 15484
rect 15841 15447 15899 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 17678 15444 17684 15496
rect 17736 15444 17742 15496
rect 18156 15484 18184 15524
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18288 15524 18429 15552
rect 18288 15512 18294 15524
rect 18417 15521 18429 15524
rect 18463 15552 18475 15555
rect 18874 15552 18880 15564
rect 18463 15524 18880 15552
rect 18463 15521 18475 15524
rect 18417 15515 18475 15521
rect 18874 15512 18880 15524
rect 18932 15512 18938 15564
rect 18969 15555 19027 15561
rect 18969 15521 18981 15555
rect 19015 15552 19027 15555
rect 19150 15552 19156 15564
rect 19015 15524 19156 15552
rect 19015 15521 19027 15524
rect 18969 15515 19027 15521
rect 18984 15484 19012 15515
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 20162 15512 20168 15564
rect 20220 15552 20226 15564
rect 20806 15552 20812 15564
rect 20220 15524 20812 15552
rect 20220 15512 20226 15524
rect 20806 15512 20812 15524
rect 20864 15552 20870 15564
rect 20993 15555 21051 15561
rect 20993 15552 21005 15555
rect 20864 15524 21005 15552
rect 20864 15512 20870 15524
rect 20993 15521 21005 15524
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 19058 15484 19064 15496
rect 18156 15456 19012 15484
rect 19019 15456 19064 15484
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 10827 15388 11790 15416
rect 11992 15388 14381 15416
rect 10827 15385 10839 15388
rect 10781 15379 10839 15385
rect 7282 15348 7288 15360
rect 6604 15320 6960 15348
rect 7243 15320 7288 15348
rect 6604 15308 6610 15320
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8110 15308 8116 15360
rect 8168 15348 8174 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 8168 15320 9321 15348
rect 8168 15308 8174 15320
rect 9309 15317 9321 15320
rect 9355 15317 9367 15351
rect 9674 15348 9680 15360
rect 9309 15311 9367 15317
rect 9646 15308 9680 15348
rect 9732 15308 9738 15360
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11992 15348 12020 15388
rect 14369 15385 14381 15388
rect 14415 15385 14427 15419
rect 14369 15379 14427 15385
rect 14921 15419 14979 15425
rect 14921 15385 14933 15419
rect 14967 15416 14979 15419
rect 17696 15416 17724 15444
rect 18049 15419 18107 15425
rect 18049 15416 18061 15419
rect 14967 15388 18061 15416
rect 14967 15385 14979 15388
rect 14921 15379 14979 15385
rect 18049 15385 18061 15388
rect 18095 15385 18107 15419
rect 18049 15379 18107 15385
rect 18138 15376 18144 15428
rect 18196 15416 18202 15428
rect 19797 15419 19855 15425
rect 19797 15416 19809 15419
rect 18196 15388 19809 15416
rect 18196 15376 18202 15388
rect 19797 15385 19809 15388
rect 19843 15385 19855 15419
rect 19797 15379 19855 15385
rect 11204 15320 12020 15348
rect 12529 15351 12587 15357
rect 11204 15308 11210 15320
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12802 15348 12808 15360
rect 12575 15320 12808 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 14093 15351 14151 15357
rect 14093 15317 14105 15351
rect 14139 15348 14151 15351
rect 15562 15348 15568 15360
rect 14139 15320 15568 15348
rect 14139 15317 14151 15320
rect 14093 15311 14151 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 15930 15308 15936 15360
rect 15988 15348 15994 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 15988 15320 16313 15348
rect 15988 15308 15994 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16666 15348 16672 15360
rect 16627 15320 16672 15348
rect 16301 15311 16359 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17678 15348 17684 15360
rect 16908 15320 17684 15348
rect 16908 15308 16914 15320
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 17770 15308 17776 15360
rect 17828 15348 17834 15360
rect 19426 15348 19432 15360
rect 17828 15320 19432 15348
rect 17828 15308 17834 15320
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 20162 15348 20168 15360
rect 20123 15320 20168 15348
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 20530 15348 20536 15360
rect 20491 15320 20536 15348
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 9646 15280 9674 15308
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 2866 15144 2872 15156
rect 2179 15116 2872 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 3970 15144 3976 15156
rect 3844 15116 3976 15144
rect 3844 15104 3850 15116
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 4246 15104 4252 15156
rect 4304 15144 4310 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 4304 15116 4905 15144
rect 4304 15104 4310 15116
rect 4893 15113 4905 15116
rect 4939 15113 4951 15147
rect 4893 15107 4951 15113
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 6454 15144 6460 15156
rect 6236 15116 6460 15144
rect 6236 15104 6242 15116
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 9646 15144 9674 15184
rect 10502 15144 10508 15156
rect 8496 15116 10508 15144
rect 1578 15076 1584 15088
rect 1539 15048 1584 15076
rect 1578 15036 1584 15048
rect 1636 15036 1642 15088
rect 2038 15036 2044 15088
rect 2096 15076 2102 15088
rect 2096 15048 4562 15076
rect 2096 15036 2102 15048
rect 2222 14968 2228 15020
rect 2280 15008 2286 15020
rect 2685 15011 2743 15017
rect 2685 15008 2697 15011
rect 2280 14980 2697 15008
rect 2280 14968 2286 14980
rect 2685 14977 2697 14980
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3200 14980 3709 15008
rect 3200 14968 3206 14980
rect 3697 14977 3709 14980
rect 3743 15008 3755 15011
rect 3786 15008 3792 15020
rect 3743 14980 3792 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 290 14900 296 14952
rect 348 14940 354 14952
rect 1397 14943 1455 14949
rect 1397 14940 1409 14943
rect 348 14912 1409 14940
rect 348 14900 354 14912
rect 1397 14909 1409 14912
rect 1443 14940 1455 14943
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1443 14912 1961 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1949 14909 1961 14912
rect 1995 14940 2007 14943
rect 2038 14940 2044 14952
rect 1995 14912 2044 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 4534 14940 4562 15048
rect 5166 15036 5172 15088
rect 5224 15076 5230 15088
rect 6822 15076 6828 15088
rect 5224 15048 6828 15076
rect 5224 15036 5230 15048
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 8386 15076 8392 15088
rect 8347 15048 8392 15076
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 15008 5779 15011
rect 7834 15008 7840 15020
rect 5767 14980 7840 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 7834 14968 7840 14980
rect 7892 15008 7898 15020
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7892 14980 7941 15008
rect 7892 14968 7898 14980
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 6270 14940 6276 14952
rect 4534 14912 6276 14940
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 1210 14832 1216 14884
rect 1268 14872 1274 14884
rect 3145 14875 3203 14881
rect 3145 14872 3157 14875
rect 1268 14844 3157 14872
rect 1268 14832 1274 14844
rect 3145 14841 3157 14844
rect 3191 14841 3203 14875
rect 3145 14835 3203 14841
rect 3605 14875 3663 14881
rect 3605 14841 3617 14875
rect 3651 14872 3663 14875
rect 4059 14875 4117 14881
rect 4059 14872 4071 14875
rect 3651 14844 4071 14872
rect 3651 14841 3663 14844
rect 3605 14835 3663 14841
rect 4059 14841 4071 14844
rect 4105 14872 4117 14875
rect 5074 14872 5080 14884
rect 4105 14844 5080 14872
rect 4105 14841 4117 14844
rect 4059 14835 4117 14841
rect 5074 14832 5080 14844
rect 5132 14872 5138 14884
rect 5258 14872 5264 14884
rect 5132 14844 5264 14872
rect 5132 14832 5138 14844
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 6917 14875 6975 14881
rect 6917 14872 6929 14875
rect 6604 14844 6929 14872
rect 6604 14832 6610 14844
rect 6917 14841 6929 14844
rect 6963 14841 6975 14875
rect 6917 14835 6975 14841
rect 7009 14875 7067 14881
rect 7009 14841 7021 14875
rect 7055 14841 7067 14875
rect 7009 14835 7067 14841
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 7607 14844 7741 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 2590 14804 2596 14816
rect 2455 14776 2596 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4488 14776 4629 14804
rect 4488 14764 4494 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 5350 14804 5356 14816
rect 5311 14776 5356 14804
rect 4617 14767 4675 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 6052 14776 6285 14804
rect 6052 14764 6058 14776
rect 6273 14773 6285 14776
rect 6319 14773 6331 14807
rect 6273 14767 6331 14773
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7024 14804 7052 14835
rect 6880 14776 7052 14804
rect 7713 14804 7741 14844
rect 7834 14832 7840 14884
rect 7892 14872 7898 14884
rect 8496 14872 8524 15116
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 8628 15048 8708 15076
rect 8628 15036 8634 15048
rect 8680 15017 8708 15048
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 9646 15076 9674 15116
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 11238 15144 11244 15156
rect 11199 15116 11244 15144
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 12575 15147 12633 15153
rect 12575 15113 12587 15147
rect 12621 15144 12633 15147
rect 14737 15147 14795 15153
rect 14737 15144 14749 15147
rect 12621 15116 13814 15144
rect 12621 15113 12633 15116
rect 12575 15107 12633 15113
rect 9180 15048 9674 15076
rect 9180 15036 9186 15048
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 11977 15079 12035 15085
rect 11977 15076 11989 15079
rect 9824 15048 11989 15076
rect 9824 15036 9830 15048
rect 11977 15045 11989 15048
rect 12023 15045 12035 15079
rect 13786 15076 13814 15116
rect 13924 15116 14749 15144
rect 13924 15076 13952 15116
rect 14737 15113 14749 15116
rect 14783 15113 14795 15147
rect 14737 15107 14795 15113
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15562 15144 15568 15156
rect 15059 15116 15568 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 16206 15104 16212 15156
rect 16264 15144 16270 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 16264 15116 16313 15144
rect 16264 15104 16270 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 16301 15107 16359 15113
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16577 15147 16635 15153
rect 16577 15144 16589 15147
rect 16439 15116 16589 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16577 15113 16589 15116
rect 16623 15144 16635 15147
rect 16942 15144 16948 15156
rect 16623 15116 16948 15144
rect 16623 15113 16635 15116
rect 16577 15107 16635 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17313 15147 17371 15153
rect 17313 15113 17325 15147
rect 17359 15144 17371 15147
rect 17494 15144 17500 15156
rect 17359 15116 17500 15144
rect 17359 15113 17371 15116
rect 17313 15107 17371 15113
rect 17494 15104 17500 15116
rect 17552 15144 17558 15156
rect 17773 15147 17831 15153
rect 17773 15144 17785 15147
rect 17552 15116 17785 15144
rect 17552 15104 17558 15116
rect 17773 15113 17785 15116
rect 17819 15113 17831 15147
rect 17773 15107 17831 15113
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20864 15116 20913 15144
rect 20864 15104 20870 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 21726 15144 21732 15156
rect 21687 15116 21732 15144
rect 20901 15107 20959 15113
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 20622 15076 20628 15088
rect 13786 15048 20628 15076
rect 11977 15039 12035 15045
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 10318 15008 10324 15020
rect 8711 14980 9674 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 9646 14940 9674 14980
rect 10060 14980 10324 15008
rect 10060 14940 10088 14980
rect 10318 14968 10324 14980
rect 10376 15008 10382 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10376 14980 10517 15008
rect 10376 14968 10382 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 12860 14980 13737 15008
rect 12860 14968 12866 14980
rect 13725 14977 13737 14980
rect 13771 15008 13783 15011
rect 13924 15008 13952 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 13771 14980 13952 15008
rect 14001 15011 14059 15017
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 14001 14977 14013 15011
rect 14047 15008 14059 15011
rect 21315 15011 21373 15017
rect 21315 15008 21327 15011
rect 14047 14980 21327 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 21315 14977 21327 14980
rect 21361 15008 21373 15011
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21361 14980 22017 15008
rect 21361 14977 21373 14980
rect 21315 14971 21373 14977
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 9646 14912 10088 14940
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 12158 14940 12164 14952
rect 11296 14912 12164 14940
rect 11296 14900 11302 14912
rect 12158 14900 12164 14912
rect 12216 14940 12222 14952
rect 12472 14943 12530 14949
rect 12472 14940 12484 14943
rect 12216 14912 12484 14940
rect 12216 14900 12222 14912
rect 12472 14909 12484 14912
rect 12518 14940 12530 14943
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12518 14912 12909 14940
rect 12518 14909 12530 14912
rect 12472 14903 12530 14909
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 15160 14912 15301 14940
rect 15160 14900 15166 14912
rect 15289 14909 15301 14912
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14940 15807 14943
rect 15838 14940 15844 14952
rect 15795 14912 15844 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16025 14943 16083 14949
rect 16025 14909 16037 14943
rect 16071 14909 16083 14943
rect 16206 14940 16212 14952
rect 16167 14912 16212 14940
rect 16025 14903 16083 14909
rect 7892 14844 8524 14872
rect 7892 14832 7898 14844
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 8812 14844 8857 14872
rect 8812 14832 8818 14844
rect 9122 14832 9128 14884
rect 9180 14872 9186 14884
rect 9309 14875 9367 14881
rect 9309 14872 9321 14875
rect 9180 14844 9321 14872
rect 9180 14832 9186 14844
rect 9309 14841 9321 14844
rect 9355 14841 9367 14875
rect 9309 14835 9367 14841
rect 9769 14875 9827 14881
rect 9769 14841 9781 14875
rect 9815 14872 9827 14875
rect 9858 14872 9864 14884
rect 9815 14844 9864 14872
rect 9815 14841 9827 14844
rect 9769 14835 9827 14841
rect 9324 14804 9352 14835
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 10229 14875 10287 14881
rect 10229 14841 10241 14875
rect 10275 14841 10287 14875
rect 10229 14835 10287 14841
rect 7713 14776 9352 14804
rect 6880 14764 6886 14776
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 10244 14804 10272 14835
rect 10318 14832 10324 14884
rect 10376 14872 10382 14884
rect 10376 14844 10421 14872
rect 10376 14832 10382 14844
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 11609 14875 11667 14881
rect 11609 14872 11621 14875
rect 11020 14844 11621 14872
rect 11020 14832 11026 14844
rect 11609 14841 11621 14844
rect 11655 14841 11667 14875
rect 11609 14835 11667 14841
rect 14093 14875 14151 14881
rect 14093 14841 14105 14875
rect 14139 14872 14151 14875
rect 14182 14872 14188 14884
rect 14139 14844 14188 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 14645 14875 14703 14881
rect 14645 14841 14657 14875
rect 14691 14872 14703 14875
rect 15010 14872 15016 14884
rect 14691 14844 15016 14872
rect 14691 14841 14703 14844
rect 14645 14835 14703 14841
rect 11146 14804 11152 14816
rect 10008 14776 11152 14804
rect 10008 14764 10014 14776
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 12713 14807 12771 14813
rect 12713 14804 12725 14807
rect 11480 14776 12725 14804
rect 11480 14764 11486 14776
rect 12713 14773 12725 14776
rect 12759 14804 12771 14807
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 12759 14776 13277 14804
rect 12759 14773 12771 14776
rect 12713 14767 12771 14773
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 13998 14764 14004 14816
rect 14056 14804 14062 14816
rect 14660 14804 14688 14835
rect 15010 14832 15016 14844
rect 15068 14832 15074 14884
rect 16040 14872 16068 14903
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 17494 14940 17500 14952
rect 16347 14912 17500 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 19061 14943 19119 14949
rect 19061 14940 19073 14943
rect 18932 14912 19073 14940
rect 18932 14900 18938 14912
rect 19061 14909 19073 14912
rect 19107 14940 19119 14943
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19107 14912 19441 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 19429 14909 19441 14912
rect 19475 14940 19487 14943
rect 19518 14940 19524 14952
rect 19475 14912 19524 14940
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 19518 14900 19524 14912
rect 19576 14940 19582 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19576 14912 19625 14940
rect 19576 14900 19582 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 19978 14900 19984 14952
rect 20036 14940 20042 14952
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 20036 14912 20085 14940
rect 20036 14900 20042 14912
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 20073 14903 20131 14909
rect 21228 14943 21286 14949
rect 21228 14909 21240 14943
rect 21274 14940 21286 14943
rect 21726 14940 21732 14952
rect 21274 14912 21732 14940
rect 21274 14909 21286 14912
rect 21228 14903 21286 14909
rect 21726 14900 21732 14912
rect 21784 14900 21790 14952
rect 16393 14875 16451 14881
rect 16393 14872 16405 14875
rect 15120 14844 16405 14872
rect 14056 14776 14688 14804
rect 14737 14807 14795 14813
rect 14056 14764 14062 14776
rect 14737 14773 14749 14807
rect 14783 14804 14795 14807
rect 15120 14804 15148 14844
rect 16393 14841 16405 14844
rect 16439 14841 16451 14875
rect 18138 14872 18144 14884
rect 16393 14835 16451 14841
rect 16592 14844 17908 14872
rect 18099 14844 18144 14872
rect 14783 14776 15148 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 16592 14804 16620 14844
rect 16850 14804 16856 14816
rect 15896 14776 16620 14804
rect 16811 14776 16856 14804
rect 15896 14764 15902 14776
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17880 14804 17908 14844
rect 18138 14832 18144 14844
rect 18196 14832 18202 14884
rect 18230 14832 18236 14884
rect 18288 14872 18294 14884
rect 18782 14872 18788 14884
rect 18288 14844 18333 14872
rect 18743 14844 18788 14872
rect 18288 14832 18294 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 18892 14844 19748 14872
rect 18892 14804 18920 14844
rect 19720 14813 19748 14844
rect 17880 14776 18920 14804
rect 19705 14807 19763 14813
rect 19705 14773 19717 14807
rect 19751 14773 19763 14807
rect 19705 14767 19763 14773
rect 290 14696 296 14748
rect 348 14736 354 14748
rect 569 14739 627 14745
rect 569 14736 581 14739
rect 348 14708 581 14736
rect 348 14696 354 14708
rect 569 14705 581 14708
rect 615 14705 627 14739
rect 569 14699 627 14705
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 566 14600 572 14612
rect 527 14572 572 14600
rect 566 14560 572 14572
rect 624 14560 630 14612
rect 1535 14603 1593 14609
rect 1535 14569 1547 14603
rect 1581 14600 1593 14603
rect 1854 14600 1860 14612
rect 1581 14572 1860 14600
rect 1581 14569 1593 14572
rect 1535 14563 1593 14569
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2038 14560 2044 14612
rect 2096 14600 2102 14612
rect 3326 14600 3332 14612
rect 2096 14572 3332 14600
rect 2096 14560 2102 14572
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 3786 14600 3792 14612
rect 3747 14572 3792 14600
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4982 14600 4988 14612
rect 3927 14572 4988 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5166 14600 5172 14612
rect 5127 14572 5172 14600
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5316 14572 5666 14600
rect 5316 14560 5322 14572
rect 2590 14532 2596 14544
rect 2551 14504 2596 14532
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 2682 14492 2688 14544
rect 2740 14532 2746 14544
rect 3510 14532 3516 14544
rect 2740 14504 3516 14532
rect 2740 14492 2746 14504
rect 3510 14492 3516 14504
rect 3568 14532 3574 14544
rect 4065 14535 4123 14541
rect 4065 14532 4077 14535
rect 3568 14504 4077 14532
rect 3568 14492 3574 14504
rect 4065 14501 4077 14504
rect 4111 14501 4123 14535
rect 5442 14532 5448 14544
rect 4065 14495 4123 14501
rect 4239 14504 5448 14532
rect 477 14467 535 14473
rect 477 14433 489 14467
rect 523 14464 535 14467
rect 566 14464 572 14476
rect 523 14436 572 14464
rect 523 14433 535 14436
rect 477 14427 535 14433
rect 566 14424 572 14436
rect 624 14424 630 14476
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 1432 14467 1490 14473
rect 1432 14464 1444 14467
rect 1360 14436 1444 14464
rect 1360 14424 1366 14436
rect 1432 14433 1444 14436
rect 1478 14433 1490 14467
rect 1432 14427 1490 14433
rect 3605 14467 3663 14473
rect 3605 14433 3617 14467
rect 3651 14464 3663 14467
rect 3694 14464 3700 14476
rect 3651 14436 3700 14464
rect 3651 14433 3663 14436
rect 3605 14427 3663 14433
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 4239 14396 4267 14504
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 5638 14541 5666 14572
rect 6270 14560 6276 14612
rect 6328 14600 6334 14612
rect 8202 14600 8208 14612
rect 6328 14572 7741 14600
rect 8163 14572 8208 14600
rect 6328 14560 6334 14572
rect 5623 14535 5681 14541
rect 5623 14501 5635 14535
rect 5669 14532 5681 14535
rect 6365 14535 6423 14541
rect 6365 14532 6377 14535
rect 5669 14504 6377 14532
rect 5669 14501 5681 14504
rect 5623 14495 5681 14501
rect 6365 14501 6377 14504
rect 6411 14532 6423 14535
rect 7606 14535 7664 14541
rect 7606 14532 7618 14535
rect 6411 14504 7618 14532
rect 6411 14501 6423 14504
rect 6365 14495 6423 14501
rect 7606 14501 7618 14504
rect 7652 14501 7664 14535
rect 7713 14532 7741 14572
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 8665 14603 8723 14609
rect 8665 14600 8677 14603
rect 8312 14572 8677 14600
rect 8312 14532 8340 14572
rect 8665 14569 8677 14572
rect 8711 14600 8723 14603
rect 8754 14600 8760 14612
rect 8711 14572 8760 14600
rect 8711 14569 8723 14572
rect 8665 14563 8723 14569
rect 7713 14504 8340 14532
rect 7606 14495 7664 14501
rect 8386 14492 8392 14544
rect 8444 14532 8450 14544
rect 8680 14532 8708 14563
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9858 14600 9864 14612
rect 8904 14572 9864 14600
rect 8904 14560 8910 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10410 14560 10416 14612
rect 10468 14600 10474 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 10468 14572 10517 14600
rect 10468 14560 10474 14572
rect 10505 14569 10517 14572
rect 10551 14569 10563 14603
rect 12802 14600 12808 14612
rect 12763 14572 12808 14600
rect 10505 14563 10563 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13357 14603 13415 14609
rect 13357 14569 13369 14603
rect 13403 14600 13415 14603
rect 13906 14600 13912 14612
rect 13403 14572 13912 14600
rect 13403 14569 13415 14572
rect 13357 14563 13415 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14001 14603 14059 14609
rect 14001 14569 14013 14603
rect 14047 14600 14059 14603
rect 14182 14600 14188 14612
rect 14047 14572 14188 14600
rect 14047 14569 14059 14572
rect 14001 14563 14059 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14323 14603 14381 14609
rect 14323 14569 14335 14603
rect 14369 14600 14381 14603
rect 15746 14600 15752 14612
rect 14369 14572 15752 14600
rect 14369 14569 14381 14572
rect 14323 14563 14381 14569
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 17310 14600 17316 14612
rect 15887 14572 17316 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 20349 14603 20407 14609
rect 20349 14600 20361 14603
rect 18104 14572 20361 14600
rect 18104 14560 18110 14572
rect 20349 14569 20361 14572
rect 20395 14569 20407 14603
rect 20349 14563 20407 14569
rect 10137 14535 10195 14541
rect 10137 14532 10149 14535
rect 8444 14504 10149 14532
rect 8444 14492 8450 14504
rect 4387 14467 4445 14473
rect 4387 14433 4399 14467
rect 4433 14464 4445 14467
rect 4433 14436 5580 14464
rect 4433 14433 4445 14436
rect 4387 14427 4445 14433
rect 2547 14368 4267 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 5261 14399 5319 14405
rect 4764 14368 4844 14396
rect 4764 14356 4770 14368
rect 4816 14340 4844 14368
rect 5261 14365 5273 14399
rect 5307 14396 5319 14399
rect 5442 14396 5448 14408
rect 5307 14368 5448 14396
rect 5307 14365 5319 14368
rect 5261 14359 5319 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 5552 14396 5580 14436
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 7285 14467 7343 14473
rect 7285 14464 7297 14467
rect 5960 14436 7297 14464
rect 5960 14424 5966 14436
rect 7285 14433 7297 14436
rect 7331 14464 7343 14467
rect 8570 14464 8576 14476
rect 7331 14436 8576 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 8680 14464 8708 14504
rect 10137 14501 10149 14504
rect 10183 14532 10195 14535
rect 10318 14532 10324 14544
rect 10183 14504 10324 14532
rect 10183 14501 10195 14504
rect 10137 14495 10195 14501
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 11051 14535 11109 14541
rect 11051 14501 11063 14535
rect 11097 14532 11109 14535
rect 12820 14532 12848 14560
rect 14734 14532 14740 14544
rect 11097 14504 12848 14532
rect 14695 14504 14740 14532
rect 11097 14501 11109 14504
rect 11051 14495 11109 14501
rect 14734 14492 14740 14504
rect 14792 14492 14798 14544
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 16301 14535 16359 14541
rect 16301 14532 16313 14535
rect 16080 14504 16313 14532
rect 16080 14492 16086 14504
rect 16301 14501 16313 14504
rect 16347 14532 16359 14535
rect 16482 14532 16488 14544
rect 16347 14504 16488 14532
rect 16347 14501 16359 14504
rect 16301 14495 16359 14501
rect 16482 14492 16488 14504
rect 16540 14492 16546 14544
rect 16850 14492 16856 14544
rect 16908 14532 16914 14544
rect 16945 14535 17003 14541
rect 16945 14532 16957 14535
rect 16908 14504 16957 14532
rect 16908 14492 16914 14504
rect 16945 14501 16957 14504
rect 16991 14532 17003 14535
rect 18506 14532 18512 14544
rect 16991 14504 18512 14532
rect 16991 14501 17003 14504
rect 16945 14495 17003 14501
rect 18506 14492 18512 14504
rect 18564 14492 18570 14544
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 19613 14535 19671 14541
rect 19613 14532 19625 14535
rect 19484 14504 19625 14532
rect 19484 14492 19490 14504
rect 19613 14501 19625 14504
rect 19659 14532 19671 14535
rect 19978 14532 19984 14544
rect 19659 14504 19984 14532
rect 19659 14501 19671 14504
rect 19613 14495 19671 14501
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 20254 14492 20260 14544
rect 20312 14532 20318 14544
rect 20714 14532 20720 14544
rect 20312 14504 20720 14532
rect 20312 14492 20318 14504
rect 20714 14492 20720 14504
rect 20772 14532 20778 14544
rect 20772 14504 21220 14532
rect 20772 14492 20778 14504
rect 9122 14464 9128 14476
rect 8680 14436 9128 14464
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9712 14467 9770 14473
rect 9712 14464 9724 14467
rect 9640 14436 9724 14464
rect 9640 14424 9646 14436
rect 9712 14433 9724 14436
rect 9758 14433 9770 14467
rect 9712 14427 9770 14433
rect 9815 14467 9873 14473
rect 9815 14433 9827 14467
rect 9861 14464 9873 14467
rect 13354 14464 13360 14476
rect 9861 14436 13360 14464
rect 9861 14433 9873 14436
rect 9815 14427 9873 14433
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13630 14424 13636 14476
rect 13688 14464 13694 14476
rect 14252 14467 14310 14473
rect 14252 14464 14264 14467
rect 13688 14436 14264 14464
rect 13688 14424 13694 14436
rect 14252 14433 14264 14436
rect 14298 14464 14310 14467
rect 14550 14464 14556 14476
rect 14298 14436 14556 14464
rect 14298 14433 14310 14436
rect 14252 14427 14310 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 15620 14436 15669 14464
rect 15620 14424 15626 14436
rect 15657 14433 15669 14436
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 15746 14424 15752 14476
rect 15804 14464 15810 14476
rect 16574 14464 16580 14476
rect 15804 14436 16580 14464
rect 15804 14424 15810 14436
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 21192 14473 21220 14504
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20864 14436 20913 14464
rect 20864 14424 20870 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 21177 14467 21235 14473
rect 21177 14433 21189 14467
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 7650 14396 7656 14408
rect 5552 14368 7656 14396
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 7926 14356 7932 14408
rect 7984 14396 7990 14408
rect 8202 14396 8208 14408
rect 7984 14368 8208 14396
rect 7984 14356 7990 14368
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 9950 14396 9956 14408
rect 8444 14368 9956 14396
rect 8444 14356 8450 14368
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 10778 14396 10784 14408
rect 10735 14368 10784 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 10778 14356 10784 14368
rect 10836 14396 10842 14408
rect 12250 14396 12256 14408
rect 10836 14368 12256 14396
rect 10836 14356 10842 14368
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 12434 14396 12440 14408
rect 12395 14368 12440 14396
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 16592 14368 16865 14396
rect 1946 14328 1952 14340
rect 1907 14300 1952 14328
rect 1946 14288 1952 14300
rect 2004 14288 2010 14340
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 2682 14328 2688 14340
rect 2464 14300 2688 14328
rect 2464 14288 2470 14300
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 3053 14331 3111 14337
rect 3053 14297 3065 14331
rect 3099 14328 3111 14331
rect 3694 14328 3700 14340
rect 3099 14300 3700 14328
rect 3099 14297 3111 14300
rect 3053 14291 3111 14297
rect 3694 14288 3700 14300
rect 3752 14288 3758 14340
rect 3878 14328 3884 14340
rect 3839 14300 3884 14328
rect 3878 14288 3884 14300
rect 3936 14288 3942 14340
rect 4798 14288 4804 14340
rect 4856 14288 4862 14340
rect 5902 14288 5908 14340
rect 5960 14328 5966 14340
rect 9309 14331 9367 14337
rect 9309 14328 9321 14331
rect 5960 14300 9321 14328
rect 5960 14288 5966 14300
rect 9309 14297 9321 14300
rect 9355 14297 9367 14331
rect 9309 14291 9367 14297
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 9858 14328 9864 14340
rect 9640 14300 9864 14328
rect 9640 14288 9646 14300
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 11609 14331 11667 14337
rect 11609 14297 11621 14331
rect 11655 14328 11667 14331
rect 15470 14328 15476 14340
rect 11655 14300 15476 14328
rect 11655 14297 11667 14300
rect 11609 14291 11667 14297
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 15565 14331 15623 14337
rect 15565 14297 15577 14331
rect 15611 14328 15623 14331
rect 15930 14328 15936 14340
rect 15611 14300 15936 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 1854 14220 1860 14272
rect 1912 14260 1918 14272
rect 2225 14263 2283 14269
rect 2225 14260 2237 14263
rect 1912 14232 2237 14260
rect 1912 14220 1918 14232
rect 2225 14229 2237 14232
rect 2271 14260 2283 14263
rect 4430 14260 4436 14272
rect 2271 14232 4436 14260
rect 2271 14229 2283 14232
rect 2225 14223 2283 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 6181 14263 6239 14269
rect 6181 14229 6193 14263
rect 6227 14260 6239 14263
rect 6362 14260 6368 14272
rect 6227 14232 6368 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 6546 14260 6552 14272
rect 6507 14232 6552 14260
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 6822 14260 6828 14272
rect 6783 14232 6828 14260
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 7984 14232 8953 14260
rect 7984 14220 7990 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 10686 14260 10692 14272
rect 9272 14232 10692 14260
rect 9272 14220 9278 14232
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11974 14260 11980 14272
rect 11935 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12158 14220 12164 14272
rect 12216 14260 12222 14272
rect 12253 14263 12311 14269
rect 12253 14260 12265 14263
rect 12216 14232 12265 14260
rect 12216 14220 12222 14232
rect 12253 14229 12265 14232
rect 12299 14229 12311 14263
rect 12253 14223 12311 14229
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14792 14232 15025 14260
rect 14792 14220 14798 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16592 14269 16620 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 17310 14396 17316 14408
rect 17271 14368 17316 14396
rect 16853 14359 16911 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 17828 14368 18429 14396
rect 17828 14356 17834 14368
rect 18417 14365 18429 14368
rect 18463 14365 18475 14399
rect 18782 14396 18788 14408
rect 18743 14368 18788 14396
rect 18417 14359 18475 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 19852 14368 21373 14396
rect 19852 14356 19858 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 19981 14331 20039 14337
rect 19981 14328 19993 14331
rect 17000 14300 19993 14328
rect 17000 14288 17006 14300
rect 19981 14297 19993 14300
rect 20027 14297 20039 14331
rect 19981 14291 20039 14297
rect 20438 14288 20444 14340
rect 20496 14328 20502 14340
rect 20993 14331 21051 14337
rect 20993 14328 21005 14331
rect 20496 14300 21005 14328
rect 20496 14288 20502 14300
rect 20993 14297 21005 14300
rect 21039 14297 21051 14331
rect 20993 14291 21051 14297
rect 16577 14263 16635 14269
rect 16577 14260 16589 14263
rect 16540 14232 16589 14260
rect 16540 14220 16546 14232
rect 16577 14229 16589 14232
rect 16623 14229 16635 14263
rect 16577 14223 16635 14229
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 18230 14260 18236 14272
rect 18187 14232 18236 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 21008 14260 21036 14291
rect 21266 14288 21272 14340
rect 21324 14328 21330 14340
rect 22281 14331 22339 14337
rect 22281 14328 22293 14331
rect 21324 14300 22293 14328
rect 21324 14288 21330 14300
rect 22281 14297 22293 14300
rect 22327 14297 22339 14331
rect 22281 14291 22339 14297
rect 21358 14260 21364 14272
rect 21008 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 22002 14260 22008 14272
rect 21963 14232 22008 14260
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 1302 14016 1308 14068
rect 1360 14056 1366 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1360 14028 1593 14056
rect 1360 14016 1366 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2498 14056 2504 14068
rect 2280 14028 2504 14056
rect 2280 14016 2286 14028
rect 2498 14016 2504 14028
rect 2556 14056 2562 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2556 14028 2605 14056
rect 2556 14016 2562 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 7006 14056 7012 14068
rect 3200 14028 7012 14056
rect 3200 14016 3206 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 8754 14056 8760 14068
rect 8435 14028 8760 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 9306 14016 9312 14068
rect 9364 14016 9370 14068
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 10594 14056 10600 14068
rect 9631 14028 10600 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11330 14056 11336 14068
rect 11195 14028 11336 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11330 14016 11336 14028
rect 11388 14056 11394 14068
rect 11606 14056 11612 14068
rect 11388 14028 11612 14056
rect 11388 14016 11394 14028
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12434 14056 12440 14068
rect 12299 14028 12440 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14182 14056 14188 14068
rect 14139 14028 14188 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14461 14059 14519 14065
rect 14461 14025 14473 14059
rect 14507 14056 14519 14059
rect 14550 14056 14556 14068
rect 14507 14028 14556 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 14826 14056 14832 14068
rect 14787 14028 14832 14056
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15059 14059 15117 14065
rect 15059 14025 15071 14059
rect 15105 14056 15117 14059
rect 15286 14056 15292 14068
rect 15105 14028 15292 14056
rect 15105 14025 15117 14028
rect 15059 14019 15117 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 16945 14059 17003 14065
rect 16945 14025 16957 14059
rect 16991 14056 17003 14059
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 16991 14028 17785 14056
rect 16991 14025 17003 14028
rect 16945 14019 17003 14025
rect 17773 14025 17785 14028
rect 17819 14056 17831 14059
rect 18230 14056 18236 14068
rect 17819 14028 18236 14056
rect 17819 14025 17831 14028
rect 17773 14019 17831 14025
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 19150 14056 19156 14068
rect 19111 14028 19156 14056
rect 19150 14016 19156 14028
rect 19208 14056 19214 14068
rect 19208 14028 19334 14056
rect 19208 14016 19214 14028
rect 1903 13991 1961 13997
rect 1903 13957 1915 13991
rect 1949 13988 1961 13991
rect 2314 13988 2320 14000
rect 1949 13960 2320 13988
rect 1949 13957 1961 13960
rect 1903 13951 1961 13957
rect 2314 13948 2320 13960
rect 2372 13948 2378 14000
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 4249 13991 4307 13997
rect 4249 13988 4261 13991
rect 3568 13960 4261 13988
rect 3568 13948 3574 13960
rect 4249 13957 4261 13960
rect 4295 13957 4307 13991
rect 4430 13988 4436 14000
rect 4391 13960 4436 13988
rect 4249 13951 4307 13957
rect 1118 13880 1124 13932
rect 1176 13920 1182 13932
rect 1302 13920 1308 13932
rect 1176 13892 1308 13920
rect 1176 13880 1182 13892
rect 1302 13880 1308 13892
rect 1360 13880 1366 13932
rect 2130 13920 2136 13932
rect 1847 13892 2136 13920
rect 1847 13861 1875 13892
rect 2130 13880 2136 13892
rect 2188 13920 2194 13932
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 2188 13892 2237 13920
rect 2188 13880 2194 13892
rect 2225 13889 2237 13892
rect 2271 13889 2283 13923
rect 4264 13920 4292 13951
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 4709 13991 4767 13997
rect 4709 13957 4721 13991
rect 4755 13988 4767 13991
rect 4798 13988 4804 14000
rect 4755 13960 4804 13988
rect 4755 13957 4767 13960
rect 4709 13951 4767 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 5718 13988 5724 14000
rect 5276 13960 5724 13988
rect 4614 13920 4620 13932
rect 4264 13892 4620 13920
rect 2225 13883 2283 13889
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 1816 13855 1875 13861
rect 1816 13821 1828 13855
rect 1862 13824 1875 13855
rect 1862 13821 1874 13824
rect 1816 13815 1874 13821
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 4816 13861 4844 13948
rect 2904 13855 2962 13861
rect 2904 13852 2916 13855
rect 2832 13824 2916 13852
rect 2832 13812 2838 13824
rect 2904 13821 2916 13824
rect 2950 13852 2962 13855
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 2950 13824 3341 13852
rect 2950 13821 2962 13824
rect 2904 13815 2962 13821
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 4890 13812 4896 13864
rect 4948 13852 4954 13864
rect 5276 13861 5304 13960
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 6457 13991 6515 13997
rect 6236 13960 6408 13988
rect 6236 13948 6242 13960
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5500 13892 5580 13920
rect 5500 13880 5506 13892
rect 5552 13861 5580 13892
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 4948 13824 5273 13852
rect 4948 13812 4954 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 5261 13815 5319 13821
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5583 13824 6193 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 3605 13787 3663 13793
rect 3605 13753 3617 13787
rect 3651 13784 3663 13787
rect 3651 13756 3924 13784
rect 3651 13753 3663 13756
rect 3605 13747 3663 13753
rect 109 13719 167 13725
rect 109 13685 121 13719
rect 155 13716 167 13719
rect 1118 13716 1124 13728
rect 155 13688 1124 13716
rect 155 13685 167 13688
rect 109 13679 167 13685
rect 1118 13676 1124 13688
rect 1176 13676 1182 13728
rect 2038 13676 2044 13728
rect 2096 13716 2102 13728
rect 2133 13719 2191 13725
rect 2133 13716 2145 13719
rect 2096 13688 2145 13716
rect 2096 13676 2102 13688
rect 2133 13685 2145 13688
rect 2179 13685 2191 13719
rect 2133 13679 2191 13685
rect 3007 13719 3065 13725
rect 3007 13685 3019 13719
rect 3053 13716 3065 13719
rect 3510 13716 3516 13728
rect 3053 13688 3516 13716
rect 3053 13685 3065 13688
rect 3007 13679 3065 13685
rect 3510 13676 3516 13688
rect 3568 13676 3574 13728
rect 3694 13716 3700 13728
rect 3655 13688 3700 13716
rect 3694 13676 3700 13688
rect 3752 13676 3758 13728
rect 3896 13648 3924 13756
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 5718 13784 5724 13796
rect 5132 13756 5724 13784
rect 5132 13744 5138 13756
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 6380 13784 6408 13960
rect 6457 13957 6469 13991
rect 6503 13988 6515 13991
rect 6503 13960 8242 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13920 6699 13923
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 6687 13892 7481 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 7469 13889 7481 13892
rect 7515 13920 7527 13923
rect 7558 13920 7564 13932
rect 7515 13892 7564 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 7834 13920 7840 13932
rect 7668 13892 7840 13920
rect 6328 13756 6408 13784
rect 6328 13744 6334 13756
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 7558 13784 7564 13796
rect 7064 13756 7564 13784
rect 7064 13744 7070 13756
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 7668 13728 7696 13892
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 8214 13920 8242 13960
rect 8570 13948 8576 14000
rect 8628 13988 8634 14000
rect 8665 13991 8723 13997
rect 8665 13988 8677 13991
rect 8628 13960 8677 13988
rect 8628 13948 8634 13960
rect 8665 13957 8677 13960
rect 8711 13957 8723 13991
rect 8665 13951 8723 13957
rect 8938 13948 8944 14000
rect 8996 13988 9002 14000
rect 9324 13988 9352 14016
rect 9674 13988 9680 14000
rect 8996 13960 9680 13988
rect 8996 13948 9002 13960
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8214 13892 9045 13920
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9324 13920 9352 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 14844 13988 14872 14016
rect 13188 13960 14872 13988
rect 9355 13923 9413 13929
rect 9355 13920 9367 13923
rect 9324 13892 9367 13920
rect 9033 13883 9091 13889
rect 9355 13889 9367 13892
rect 9401 13889 9413 13923
rect 9355 13883 9413 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10410 13920 10416 13932
rect 10275 13892 10416 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 13188 13929 13216 13960
rect 16758 13948 16764 14000
rect 16816 13988 16822 14000
rect 17402 13988 17408 14000
rect 16816 13960 17408 13988
rect 16816 13948 16822 13960
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19306 13988 19334 14028
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20864 14028 20913 14056
rect 20864 14016 20870 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 22189 14059 22247 14065
rect 22189 14056 22201 14059
rect 20901 14019 20959 14025
rect 21227 14028 22201 14056
rect 18748 13960 18920 13988
rect 19306 13960 20208 13988
rect 18748 13948 18754 13960
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 16942 13920 16948 13932
rect 15160 13892 16948 13920
rect 15160 13880 15166 13892
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 18417 13923 18475 13929
rect 18417 13920 18429 13923
rect 17368 13892 18429 13920
rect 17368 13880 17374 13892
rect 18417 13889 18429 13892
rect 18463 13889 18475 13923
rect 18892 13920 18920 13960
rect 20180 13920 20208 13960
rect 20990 13920 20996 13932
rect 18892 13892 19334 13920
rect 18417 13883 18475 13889
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9252 13855 9310 13861
rect 9252 13852 9264 13855
rect 9180 13824 9264 13852
rect 9180 13812 9186 13824
rect 9252 13821 9264 13824
rect 9298 13852 9310 13855
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9298 13824 9781 13852
rect 9298 13821 9310 13824
rect 9252 13815 9310 13821
rect 9769 13821 9781 13824
rect 9815 13852 9827 13855
rect 11882 13852 11888 13864
rect 9815 13824 11888 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 11882 13812 11888 13824
rect 11940 13852 11946 13864
rect 12894 13852 12900 13864
rect 11940 13824 12900 13852
rect 11940 13812 11946 13824
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14826 13852 14832 13864
rect 14240 13824 14832 13852
rect 14240 13812 14246 13824
rect 14826 13812 14832 13824
rect 14884 13852 14890 13864
rect 14956 13855 15014 13861
rect 14956 13852 14968 13855
rect 14884 13824 14968 13852
rect 14884 13812 14890 13824
rect 14956 13821 14968 13824
rect 15002 13852 15014 13855
rect 15381 13855 15439 13861
rect 15381 13852 15393 13855
rect 15002 13824 15393 13852
rect 15002 13821 15014 13824
rect 14956 13815 15014 13821
rect 15381 13821 15393 13824
rect 15427 13821 15439 13855
rect 16022 13852 16028 13864
rect 15983 13824 16028 13852
rect 15381 13815 15439 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 17862 13852 17868 13864
rect 16632 13824 17868 13852
rect 16632 13812 16638 13824
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 19306 13852 19334 13892
rect 20180 13892 20996 13920
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19306 13824 19533 13852
rect 19521 13821 19533 13824
rect 19567 13852 19579 13855
rect 19794 13852 19800 13864
rect 19567 13824 19800 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 20180 13861 20208 13892
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 21227 13861 21255 14028
rect 22189 14025 22201 14028
rect 22235 14056 22247 14059
rect 23474 14056 23480 14068
rect 22235 14028 23480 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 21361 13991 21419 13997
rect 21361 13957 21373 13991
rect 21407 13988 21419 13991
rect 23566 13988 23572 14000
rect 21407 13960 23572 13988
rect 21407 13957 21419 13960
rect 21361 13951 21419 13957
rect 23566 13948 23572 13960
rect 23624 13948 23630 14000
rect 20165 13855 20223 13861
rect 20165 13821 20177 13855
rect 20211 13821 20223 13855
rect 20165 13815 20223 13821
rect 21177 13855 21255 13861
rect 21177 13821 21189 13855
rect 21223 13824 21255 13855
rect 21223 13821 21235 13824
rect 21177 13815 21235 13821
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 21729 13855 21787 13861
rect 21729 13852 21741 13855
rect 21416 13824 21741 13852
rect 21416 13812 21422 13824
rect 21729 13821 21741 13824
rect 21775 13821 21787 13855
rect 21729 13815 21787 13821
rect 7790 13787 7848 13793
rect 7790 13784 7802 13787
rect 7760 13756 7802 13784
rect 4433 13719 4491 13725
rect 4433 13685 4445 13719
rect 4479 13716 4491 13719
rect 5442 13716 5448 13728
rect 4479 13688 5448 13716
rect 4479 13685 4491 13688
rect 4433 13679 4491 13685
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 5813 13719 5871 13725
rect 5813 13716 5825 13719
rect 5552 13688 5825 13716
rect 5552 13648 5580 13688
rect 5813 13685 5825 13688
rect 5859 13716 5871 13719
rect 6365 13719 6423 13725
rect 6365 13716 6377 13719
rect 5859 13688 6377 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 6365 13685 6377 13688
rect 6411 13716 6423 13719
rect 6454 13716 6460 13728
rect 6411 13688 6460 13716
rect 6411 13685 6423 13688
rect 6365 13679 6423 13685
rect 6454 13676 6460 13688
rect 6512 13716 6518 13728
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 6512 13688 7297 13716
rect 6512 13676 6518 13688
rect 7285 13685 7297 13688
rect 7331 13716 7343 13719
rect 7374 13716 7380 13728
rect 7331 13688 7380 13716
rect 7331 13685 7343 13688
rect 7285 13679 7343 13685
rect 7374 13676 7380 13688
rect 7432 13716 7438 13728
rect 7650 13716 7656 13728
rect 7432 13688 7656 13716
rect 7432 13676 7438 13688
rect 7650 13676 7656 13688
rect 7708 13716 7714 13728
rect 7760 13716 7788 13756
rect 7790 13753 7802 13756
rect 7836 13753 7848 13787
rect 7790 13747 7848 13753
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 9398 13784 9404 13796
rect 8904 13756 9404 13784
rect 8904 13744 8910 13756
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 10550 13787 10608 13793
rect 10550 13784 10562 13787
rect 10428 13756 10562 13784
rect 10428 13728 10456 13756
rect 10550 13753 10562 13756
rect 10596 13753 10608 13787
rect 10550 13747 10608 13753
rect 10686 13744 10692 13796
rect 10744 13784 10750 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 10744 13756 11805 13784
rect 10744 13744 10750 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 13494 13787 13552 13793
rect 13494 13753 13506 13787
rect 13540 13753 13552 13787
rect 13494 13747 13552 13753
rect 7708 13688 7788 13716
rect 7708 13676 7714 13688
rect 8202 13676 8208 13728
rect 8260 13716 8266 13728
rect 8478 13716 8484 13728
rect 8260 13688 8484 13716
rect 8260 13676 8266 13688
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 9674 13716 9680 13728
rect 9631 13688 9680 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 10137 13719 10195 13725
rect 10137 13685 10149 13719
rect 10183 13716 10195 13719
rect 10410 13716 10416 13728
rect 10183 13688 10416 13716
rect 10183 13685 10195 13688
rect 10137 13679 10195 13685
rect 10410 13676 10416 13688
rect 10468 13716 10474 13728
rect 11425 13719 11483 13725
rect 11425 13716 11437 13719
rect 10468 13688 11437 13716
rect 10468 13676 10474 13688
rect 11425 13685 11437 13688
rect 11471 13716 11483 13719
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 11471 13688 12633 13716
rect 11471 13685 11483 13688
rect 11425 13679 11483 13685
rect 12621 13685 12633 13688
rect 12667 13716 12679 13719
rect 12802 13716 12808 13728
rect 12667 13688 12808 13716
rect 12667 13685 12679 13688
rect 12621 13679 12679 13685
rect 12802 13676 12808 13688
rect 12860 13716 12866 13728
rect 12989 13719 13047 13725
rect 12989 13716 13001 13719
rect 12860 13688 13001 13716
rect 12860 13676 12866 13688
rect 12989 13685 13001 13688
rect 13035 13716 13047 13719
rect 13170 13716 13176 13728
rect 13035 13688 13176 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 13170 13676 13176 13688
rect 13228 13716 13234 13728
rect 13509 13716 13537 13747
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 15841 13787 15899 13793
rect 15841 13784 15853 13787
rect 15620 13756 15853 13784
rect 15620 13744 15626 13756
rect 15841 13753 15853 13756
rect 15887 13784 15899 13787
rect 18141 13787 18199 13793
rect 15887 13756 17816 13784
rect 15887 13753 15899 13756
rect 15841 13747 15899 13753
rect 13228 13688 13537 13716
rect 13228 13676 13234 13688
rect 14734 13676 14740 13728
rect 14792 13716 14798 13728
rect 15470 13716 15476 13728
rect 14792 13688 15476 13716
rect 14792 13676 14798 13688
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 17221 13719 17279 13725
rect 17221 13716 17233 13719
rect 16908 13688 17233 13716
rect 16908 13676 16914 13688
rect 17221 13685 17233 13688
rect 17267 13685 17279 13719
rect 17788 13716 17816 13756
rect 18141 13753 18153 13787
rect 18187 13753 18199 13787
rect 18141 13747 18199 13753
rect 17862 13716 17868 13728
rect 17788 13688 17868 13716
rect 17221 13679 17279 13685
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 18156 13716 18184 13747
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 18288 13756 18333 13784
rect 18288 13744 18294 13756
rect 18322 13716 18328 13728
rect 18156 13688 18328 13716
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 19705 13719 19763 13725
rect 19705 13716 19717 13719
rect 19392 13688 19717 13716
rect 19392 13676 19398 13688
rect 19705 13685 19717 13688
rect 19751 13685 19763 13719
rect 19705 13679 19763 13685
rect 1104 13626 22816 13648
rect 477 13583 535 13589
rect 477 13549 489 13583
rect 523 13580 535 13583
rect 845 13583 903 13589
rect 845 13580 857 13583
rect 523 13552 857 13580
rect 523 13549 535 13552
rect 477 13543 535 13549
rect 845 13549 857 13552
rect 891 13549 903 13583
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 845 13543 903 13549
rect 753 13515 811 13521
rect 753 13481 765 13515
rect 799 13512 811 13515
rect 1029 13515 1087 13521
rect 1029 13512 1041 13515
rect 799 13484 1041 13512
rect 799 13481 811 13484
rect 753 13475 811 13481
rect 1029 13481 1041 13484
rect 1075 13481 1087 13515
rect 1029 13475 1087 13481
rect 1118 13472 1124 13524
rect 1176 13512 1182 13524
rect 2590 13512 2596 13524
rect 1176 13484 2596 13512
rect 1176 13472 1182 13484
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 3896 13456 3924 13552
rect 845 13447 903 13453
rect 845 13413 857 13447
rect 891 13444 903 13447
rect 2317 13447 2375 13453
rect 2317 13444 2329 13447
rect 891 13416 2329 13444
rect 891 13413 903 13416
rect 845 13407 903 13413
rect 2317 13413 2329 13416
rect 2363 13444 2375 13447
rect 2498 13444 2504 13456
rect 2363 13416 2504 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 2498 13404 2504 13416
rect 2556 13444 2562 13456
rect 3513 13447 3571 13453
rect 3513 13444 3525 13447
rect 2556 13416 3525 13444
rect 2556 13404 2562 13416
rect 3513 13413 3525 13416
rect 3559 13444 3571 13447
rect 3694 13444 3700 13456
rect 3559 13416 3700 13444
rect 3559 13413 3571 13416
rect 3513 13407 3571 13413
rect 3694 13404 3700 13416
rect 3752 13404 3758 13456
rect 3878 13404 3884 13456
rect 3936 13404 3942 13456
rect 4890 13404 4896 13456
rect 4948 13444 4954 13456
rect 5490 13447 5548 13453
rect 5490 13444 5502 13447
rect 4948 13416 5502 13444
rect 4948 13404 4954 13416
rect 5490 13413 5502 13416
rect 5536 13444 5548 13447
rect 5552 13444 5580 13552
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 6052 13484 6101 13512
rect 6052 13472 6058 13484
rect 6089 13481 6101 13484
rect 6135 13512 6147 13515
rect 7055 13515 7113 13521
rect 6135 13484 6868 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 5536 13416 5580 13444
rect 5536 13413 5548 13416
rect 5490 13407 5548 13413
rect 5626 13404 5632 13456
rect 5684 13444 5690 13456
rect 6733 13447 6791 13453
rect 6733 13444 6745 13447
rect 5684 13416 6745 13444
rect 5684 13404 5690 13416
rect 6733 13413 6745 13416
rect 6779 13413 6791 13447
rect 6840 13444 6868 13484
rect 7055 13481 7067 13515
rect 7101 13512 7113 13515
rect 8386 13512 8392 13524
rect 7101 13484 8392 13512
rect 7101 13481 7113 13484
rect 7055 13475 7113 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 10778 13472 10784 13524
rect 10836 13512 10842 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10836 13484 10885 13512
rect 10836 13472 10842 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11112 13484 12204 13512
rect 11112 13472 11118 13484
rect 8113 13447 8171 13453
rect 8113 13444 8125 13447
rect 6840 13416 8125 13444
rect 6733 13407 6791 13413
rect 8113 13413 8125 13416
rect 8159 13444 8171 13447
rect 8754 13444 8760 13456
rect 8159 13416 8760 13444
rect 8159 13413 8171 13416
rect 8113 13407 8171 13413
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 10039 13447 10097 13453
rect 10039 13413 10051 13447
rect 10085 13444 10097 13447
rect 10410 13444 10416 13456
rect 10085 13416 10416 13444
rect 10085 13413 10097 13416
rect 10039 13407 10097 13413
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 11609 13447 11667 13453
rect 11609 13413 11621 13447
rect 11655 13444 11667 13447
rect 11882 13444 11888 13456
rect 11655 13416 11888 13444
rect 11655 13413 11667 13416
rect 11609 13407 11667 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 12176 13444 12204 13484
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12437 13515 12495 13521
rect 12437 13512 12449 13515
rect 12308 13484 12449 13512
rect 12308 13472 12314 13484
rect 12437 13481 12449 13484
rect 12483 13481 12495 13515
rect 12437 13475 12495 13481
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 15930 13512 15936 13524
rect 13955 13484 15936 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18104 13484 18368 13512
rect 18104 13472 18110 13484
rect 12342 13444 12348 13456
rect 12032 13416 12348 13444
rect 12032 13404 12038 13416
rect 109 13379 167 13385
rect 109 13345 121 13379
rect 155 13376 167 13379
rect 1486 13376 1492 13388
rect 155 13348 1492 13376
rect 155 13345 167 13348
rect 109 13339 167 13345
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 1854 13376 1860 13388
rect 1636 13348 1860 13376
rect 1636 13336 1642 13348
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 4224 13379 4282 13385
rect 4224 13345 4236 13379
rect 4270 13376 4282 13379
rect 4338 13376 4344 13388
rect 4270 13348 4344 13376
rect 4270 13345 4282 13348
rect 4224 13339 4282 13345
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 4430 13336 4436 13388
rect 4488 13376 4494 13388
rect 7006 13385 7012 13388
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 4488 13348 5181 13376
rect 4488 13336 4494 13348
rect 5169 13345 5181 13348
rect 5215 13376 5227 13379
rect 6365 13379 6423 13385
rect 6365 13376 6377 13379
rect 5215 13348 6377 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 6365 13345 6377 13348
rect 6411 13345 6423 13379
rect 6365 13339 6423 13345
rect 6984 13379 7012 13385
rect 6984 13345 6996 13379
rect 6984 13339 7012 13345
rect 7006 13336 7012 13339
rect 7064 13336 7070 13388
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7432 13348 7481 13376
rect 7432 13336 7438 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 12176 13376 12204 13416
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 13310 13447 13368 13453
rect 13310 13444 13322 13447
rect 13228 13416 13322 13444
rect 13228 13404 13234 13416
rect 13310 13413 13322 13416
rect 13356 13444 13368 13447
rect 15749 13447 15807 13453
rect 15749 13444 15761 13447
rect 13356 13416 15761 13444
rect 13356 13413 13368 13416
rect 13310 13407 13368 13413
rect 13924 13388 13952 13416
rect 15749 13413 15761 13416
rect 15795 13444 15807 13447
rect 16025 13447 16083 13453
rect 16025 13444 16037 13447
rect 15795 13416 16037 13444
rect 15795 13413 15807 13416
rect 15749 13407 15807 13413
rect 16025 13413 16037 13416
rect 16071 13444 16083 13447
rect 16117 13447 16175 13453
rect 16117 13444 16129 13447
rect 16071 13416 16129 13444
rect 16071 13413 16083 13416
rect 16025 13407 16083 13413
rect 16117 13413 16129 13416
rect 16163 13444 16175 13447
rect 16393 13447 16451 13453
rect 16393 13444 16405 13447
rect 16163 13416 16405 13444
rect 16163 13413 16175 13416
rect 16117 13407 16175 13413
rect 16393 13413 16405 13416
rect 16439 13413 16451 13447
rect 16666 13444 16672 13456
rect 16627 13416 16672 13444
rect 16393 13407 16451 13413
rect 16666 13404 16672 13416
rect 16724 13404 16730 13456
rect 18230 13444 18236 13456
rect 18191 13416 18236 13444
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 18340 13444 18368 13484
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 19061 13515 19119 13521
rect 19061 13512 19073 13515
rect 18564 13484 19073 13512
rect 18564 13472 18570 13484
rect 19061 13481 19073 13484
rect 19107 13481 19119 13515
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 19061 13475 19119 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 20898 13472 20904 13524
rect 20956 13512 20962 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 20956 13484 21005 13512
rect 20956 13472 20962 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 20257 13447 20315 13453
rect 20257 13444 20269 13447
rect 18340 13416 20269 13444
rect 20257 13413 20269 13416
rect 20303 13413 20315 13447
rect 20257 13407 20315 13413
rect 12434 13376 12440 13388
rect 12176 13348 12440 13376
rect 7469 13339 7527 13345
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13906 13336 13912 13388
rect 13964 13336 13970 13388
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 15356 13379 15414 13385
rect 14424 13348 14688 13376
rect 14424 13336 14430 13348
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 2314 13308 2320 13320
rect 2271 13280 2320 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 2866 13308 2872 13320
rect 2827 13280 2872 13308
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 6454 13308 6460 13320
rect 4126 13280 6460 13308
rect 382 13200 388 13252
rect 440 13240 446 13252
rect 753 13243 811 13249
rect 753 13240 765 13243
rect 440 13212 765 13240
rect 440 13200 446 13212
rect 753 13209 765 13212
rect 799 13209 811 13243
rect 753 13203 811 13209
rect 1118 13200 1124 13252
rect 1176 13240 1182 13252
rect 1949 13243 2007 13249
rect 1949 13240 1961 13243
rect 1176 13212 1961 13240
rect 1176 13200 1182 13212
rect 1949 13209 1961 13212
rect 1995 13209 2007 13243
rect 1949 13203 2007 13209
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 2498 13240 2504 13252
rect 2096 13212 2504 13240
rect 2096 13200 2102 13212
rect 2498 13200 2504 13212
rect 2556 13240 2562 13252
rect 4126 13240 4154 13280
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13308 8079 13311
rect 9582 13308 9588 13320
rect 8067 13280 9588 13308
rect 8067 13277 8079 13280
rect 8021 13271 8079 13277
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9950 13308 9956 13320
rect 9723 13280 9956 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 12158 13308 12164 13320
rect 11563 13280 12164 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12308 13280 13001 13308
rect 12308 13268 12314 13280
rect 12989 13277 13001 13280
rect 13035 13308 13047 13311
rect 13262 13308 13268 13320
rect 13035 13280 13268 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 2556 13212 4154 13240
rect 2556 13200 2562 13212
rect 4614 13200 4620 13252
rect 4672 13240 4678 13252
rect 4982 13240 4988 13252
rect 4672 13212 4988 13240
rect 4672 13200 4678 13212
rect 4982 13200 4988 13212
rect 5040 13200 5046 13252
rect 8570 13240 8576 13252
rect 8531 13212 8576 13240
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 12066 13240 12072 13252
rect 8680 13212 11468 13240
rect 11979 13212 12072 13240
rect 1029 13175 1087 13181
rect 1029 13172 1041 13175
rect 952 13144 1041 13172
rect 952 12968 980 13144
rect 1029 13141 1041 13144
rect 1075 13141 1087 13175
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1029 13135 1087 13141
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 2314 13132 2320 13184
rect 2372 13172 2378 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 2372 13144 3157 13172
rect 2372 13132 2378 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 3145 13135 3203 13141
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3602 13172 3608 13184
rect 3384 13144 3608 13172
rect 3384 13132 3390 13144
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 4295 13175 4353 13181
rect 4295 13141 4307 13175
rect 4341 13172 4353 13175
rect 4430 13172 4436 13184
rect 4341 13144 4436 13172
rect 4341 13141 4353 13144
rect 4295 13135 4353 13141
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 4801 13175 4859 13181
rect 4801 13172 4813 13175
rect 4764 13144 4813 13172
rect 4764 13132 4770 13144
rect 4801 13141 4813 13144
rect 4847 13141 4859 13175
rect 4801 13135 4859 13141
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8018 13172 8024 13184
rect 7708 13144 8024 13172
rect 7708 13132 7714 13144
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 8680 13172 8708 13212
rect 8444 13144 8708 13172
rect 8444 13132 8450 13144
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 8904 13144 8953 13172
rect 8904 13132 8910 13144
rect 8941 13141 8953 13144
rect 8987 13141 8999 13175
rect 9306 13172 9312 13184
rect 9267 13144 9312 13172
rect 8941 13135 8999 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 11238 13172 11244 13184
rect 11199 13144 11244 13172
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 11440 13172 11468 13212
rect 12066 13200 12072 13212
rect 12124 13240 12130 13252
rect 12434 13240 12440 13252
rect 12124 13212 12440 13240
rect 12124 13200 12130 13212
rect 12434 13200 12440 13212
rect 12492 13200 12498 13252
rect 14660 13184 14688 13348
rect 15356 13345 15368 13379
rect 15402 13376 15414 13379
rect 15562 13376 15568 13388
rect 15402 13348 15568 13376
rect 15402 13345 15414 13348
rect 15356 13339 15414 13345
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 18874 13336 18880 13388
rect 18932 13376 18938 13388
rect 19426 13376 19432 13388
rect 18932 13348 19432 13376
rect 18932 13336 18938 13348
rect 19426 13336 19432 13348
rect 19484 13376 19490 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19484 13348 19717 13376
rect 19484 13336 19490 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20864 13348 20913 13376
rect 20864 13336 20870 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 20990 13336 20996 13388
rect 21048 13376 21054 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 21048 13348 21465 13376
rect 21048 13336 21054 13348
rect 21453 13345 21465 13348
rect 21499 13376 21511 13379
rect 22094 13376 22100 13388
rect 21499 13348 22100 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 15212 13280 16589 13308
rect 15212 13184 15240 13280
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13308 17279 13311
rect 17310 13308 17316 13320
rect 17267 13280 17316 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17310 13268 17316 13280
rect 17368 13308 17374 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17368 13280 18153 13308
rect 17368 13268 17374 13280
rect 18141 13277 18153 13280
rect 18187 13308 18199 13311
rect 18506 13308 18512 13320
rect 18187 13280 18512 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 18656 13280 18701 13308
rect 18656 13268 18662 13280
rect 17589 13243 17647 13249
rect 15442 13212 16620 13240
rect 12805 13175 12863 13181
rect 12805 13172 12817 13175
rect 11440 13144 12817 13172
rect 12805 13141 12817 13144
rect 12851 13141 12863 13175
rect 14550 13172 14556 13184
rect 14511 13144 14556 13172
rect 12805 13135 12863 13141
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 15105 13175 15163 13181
rect 15105 13141 15117 13175
rect 15151 13172 15163 13175
rect 15194 13172 15200 13184
rect 15151 13144 15200 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 15442 13181 15470 13212
rect 16592 13184 16620 13212
rect 17589 13209 17601 13243
rect 17635 13240 17647 13243
rect 18322 13240 18328 13252
rect 17635 13212 18328 13240
rect 17635 13209 17647 13212
rect 17589 13203 17647 13209
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 19889 13243 19947 13249
rect 19889 13209 19901 13243
rect 19935 13240 19947 13243
rect 22554 13240 22560 13252
rect 19935 13212 22560 13240
rect 19935 13209 19947 13212
rect 19889 13203 19947 13209
rect 22554 13200 22560 13212
rect 22612 13200 22618 13252
rect 15427 13175 15485 13181
rect 15427 13172 15439 13175
rect 15344 13144 15439 13172
rect 15344 13132 15350 13144
rect 15427 13141 15439 13144
rect 15473 13141 15485 13175
rect 16022 13172 16028 13184
rect 15983 13144 16028 13172
rect 15427 13135 15485 13141
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16574 13132 16580 13184
rect 16632 13132 16638 13184
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 17770 13172 17776 13184
rect 16908 13144 17776 13172
rect 16908 13132 16914 13144
rect 17770 13132 17776 13144
rect 17828 13172 17834 13184
rect 17865 13175 17923 13181
rect 17865 13172 17877 13175
rect 17828 13144 17877 13172
rect 17828 13132 17834 13144
rect 17865 13141 17877 13144
rect 17911 13141 17923 13175
rect 17865 13135 17923 13141
rect 18414 13132 18420 13184
rect 18472 13172 18478 13184
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 18472 13144 19441 13172
rect 18472 13132 18478 13144
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 21910 13172 21916 13184
rect 21871 13144 21916 13172
rect 19429 13135 19487 13141
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 22278 13172 22284 13184
rect 22239 13144 22284 13172
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 1578 12968 1584 12980
rect 952 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 4111 12971 4169 12977
rect 4111 12968 4123 12971
rect 1820 12940 4123 12968
rect 1820 12928 1826 12940
rect 4111 12937 4123 12940
rect 4157 12937 4169 12971
rect 4111 12931 4169 12937
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 5810 12968 5816 12980
rect 4488 12940 5816 12968
rect 4488 12928 4494 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6822 12968 6828 12980
rect 5951 12940 6828 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 8754 12968 8760 12980
rect 8527 12940 8760 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9582 12968 9588 12980
rect 9272 12940 9588 12968
rect 9272 12928 9278 12940
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 10594 12968 10600 12980
rect 10555 12940 10600 12968
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 12066 12968 12072 12980
rect 11440 12940 12072 12968
rect 2958 12860 2964 12912
rect 3016 12900 3022 12912
rect 3418 12900 3424 12912
rect 3016 12872 3424 12900
rect 3016 12860 3022 12872
rect 3418 12860 3424 12872
rect 3476 12860 3482 12912
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 5442 12900 5448 12912
rect 3936 12872 5448 12900
rect 3936 12860 3942 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 7101 12903 7159 12909
rect 7101 12900 7113 12903
rect 7064 12872 7113 12900
rect 7064 12860 7070 12872
rect 7101 12869 7113 12872
rect 7147 12900 7159 12903
rect 7650 12900 7656 12912
rect 7147 12872 7656 12900
rect 7147 12869 7159 12872
rect 7101 12863 7159 12869
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 8113 12903 8171 12909
rect 8113 12869 8125 12903
rect 8159 12900 8171 12903
rect 9306 12900 9312 12912
rect 8159 12872 9312 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 11440 12909 11468 12940
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12250 12968 12256 12980
rect 12211 12940 12256 12968
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 13906 12968 13912 12980
rect 13863 12940 13912 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 13906 12928 13912 12940
rect 13964 12968 13970 12980
rect 14090 12968 14096 12980
rect 13964 12940 14096 12968
rect 13964 12928 13970 12940
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 16942 12968 16948 12980
rect 16715 12940 16948 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 20901 12971 20959 12977
rect 20901 12968 20913 12971
rect 20864 12940 20913 12968
rect 20864 12928 20870 12940
rect 20901 12937 20913 12940
rect 20947 12937 20959 12971
rect 20901 12931 20959 12937
rect 21361 12971 21419 12977
rect 21361 12937 21373 12971
rect 21407 12968 21419 12971
rect 21542 12968 21548 12980
rect 21407 12940 21548 12968
rect 21407 12937 21419 12940
rect 21361 12931 21419 12937
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 22094 12968 22100 12980
rect 22055 12940 22100 12968
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 11425 12903 11483 12909
rect 11425 12900 11437 12903
rect 10560 12872 11437 12900
rect 10560 12860 10566 12872
rect 11425 12869 11437 12872
rect 11471 12869 11483 12903
rect 11425 12863 11483 12869
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 11974 12900 11980 12912
rect 11756 12872 11980 12900
rect 11756 12860 11762 12872
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 12084 12900 12112 12928
rect 14366 12900 14372 12912
rect 12084 12872 14372 12900
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 14829 12903 14887 12909
rect 14829 12869 14841 12903
rect 14875 12900 14887 12903
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 14875 12872 17417 12900
rect 14875 12869 14887 12872
rect 14829 12863 14887 12869
rect 17405 12869 17417 12872
rect 17451 12900 17463 12903
rect 18230 12900 18236 12912
rect 17451 12872 18236 12900
rect 17451 12869 17463 12872
rect 17405 12863 17463 12869
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 21450 12900 21456 12912
rect 18340 12872 21456 12900
rect 14 12792 20 12844
rect 72 12832 78 12844
rect 1673 12835 1731 12841
rect 72 12804 1475 12832
rect 72 12792 78 12804
rect 1447 12773 1475 12804
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 1762 12832 1768 12844
rect 1719 12804 1768 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 3142 12832 3148 12844
rect 2547 12804 3148 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3510 12832 3516 12844
rect 3292 12804 3516 12832
rect 3292 12792 3298 12804
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5626 12832 5632 12844
rect 5031 12804 5632 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 6604 12804 7205 12832
rect 6604 12792 6610 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7374 12792 7380 12844
rect 7432 12792 7438 12844
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9398 12832 9404 12844
rect 9079 12804 9404 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9858 12832 9864 12844
rect 9723 12804 9864 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 13630 12832 13636 12844
rect 10520 12804 13636 12832
rect 1432 12767 1490 12773
rect 1432 12733 1444 12767
rect 1478 12764 1490 12767
rect 1857 12767 1915 12773
rect 1857 12764 1869 12767
rect 1478 12736 1869 12764
rect 1478 12733 1490 12736
rect 1432 12727 1490 12733
rect 1857 12733 1869 12736
rect 1903 12733 1915 12767
rect 1857 12727 1915 12733
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3384 12736 3801 12764
rect 3384 12724 3390 12736
rect 3789 12733 3801 12736
rect 3835 12764 3847 12767
rect 3878 12764 3884 12776
rect 3835 12736 3884 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 4040 12767 4098 12773
rect 4040 12733 4052 12767
rect 4086 12764 4098 12767
rect 4086 12736 4292 12764
rect 4086 12733 4098 12736
rect 4040 12727 4098 12733
rect 1946 12656 1952 12708
rect 2004 12696 2010 12708
rect 2593 12699 2651 12705
rect 2004 12668 2452 12696
rect 2004 12656 2010 12668
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 2225 12631 2283 12637
rect 2225 12628 2237 12631
rect 1728 12600 2237 12628
rect 1728 12588 1734 12600
rect 2225 12597 2237 12600
rect 2271 12597 2283 12631
rect 2424 12628 2452 12668
rect 2593 12665 2605 12699
rect 2639 12665 2651 12699
rect 3142 12696 3148 12708
rect 3103 12668 3148 12696
rect 2593 12659 2651 12665
rect 2608 12628 2636 12659
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 4264 12696 4292 12736
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 4525 12767 4583 12773
rect 4525 12764 4537 12767
rect 4396 12736 4537 12764
rect 4396 12724 4402 12736
rect 4525 12733 4537 12736
rect 4571 12764 4583 12767
rect 7392 12764 7420 12792
rect 4571 12736 8892 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 4798 12696 4804 12708
rect 3292 12668 4154 12696
rect 4264 12668 4804 12696
rect 3292 12656 3298 12668
rect 3970 12628 3976 12640
rect 2424 12600 3976 12628
rect 2225 12591 2283 12597
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4126 12628 4154 12668
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5306 12699 5364 12705
rect 5306 12696 5318 12699
rect 4948 12668 5318 12696
rect 4948 12656 4954 12668
rect 5306 12665 5318 12668
rect 5352 12665 5364 12699
rect 5306 12659 5364 12665
rect 5718 12656 5724 12708
rect 5776 12696 5782 12708
rect 6822 12696 6828 12708
rect 5776 12668 6828 12696
rect 5776 12656 5782 12668
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 7392 12696 7420 12736
rect 7514 12699 7572 12705
rect 7514 12696 7526 12699
rect 7392 12668 7526 12696
rect 7514 12665 7526 12668
rect 7560 12665 7572 12699
rect 7514 12659 7572 12665
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 8202 12696 8208 12708
rect 7800 12668 8208 12696
rect 7800 12656 7806 12668
rect 8202 12656 8208 12668
rect 8260 12656 8266 12708
rect 5626 12628 5632 12640
rect 4126 12600 5632 12628
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 6052 12600 6193 12628
rect 6052 12588 6058 12600
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 6181 12591 6239 12597
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 8570 12628 8576 12640
rect 7432 12600 8576 12628
rect 7432 12588 7438 12600
rect 8570 12588 8576 12600
rect 8628 12628 8634 12640
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8628 12600 8769 12628
rect 8628 12588 8634 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 8864 12628 8892 12736
rect 9125 12699 9183 12705
rect 9125 12665 9137 12699
rect 9171 12696 9183 12699
rect 9306 12696 9312 12708
rect 9171 12668 9312 12696
rect 9171 12665 9183 12668
rect 9125 12659 9183 12665
rect 9306 12656 9312 12668
rect 9364 12656 9370 12708
rect 10520 12696 10548 12804
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 16758 12832 16764 12844
rect 15703 12804 16764 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 18340 12832 18368 12872
rect 21450 12860 21456 12872
rect 21508 12900 21514 12912
rect 22646 12900 22652 12912
rect 21508 12872 22652 12900
rect 21508 12860 21514 12872
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 18782 12832 18788 12844
rect 16868 12804 18368 12832
rect 18743 12804 18788 12832
rect 12472 12767 12530 12773
rect 12472 12764 12484 12767
rect 11761 12736 12484 12764
rect 10870 12696 10876 12708
rect 9416 12668 10548 12696
rect 10831 12668 10876 12696
rect 9416 12628 9444 12668
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 10965 12699 11023 12705
rect 10965 12665 10977 12699
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 8864 12600 9444 12628
rect 10045 12631 10103 12637
rect 8757 12591 8815 12597
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10410 12628 10416 12640
rect 10091 12600 10416 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10410 12588 10416 12600
rect 10468 12628 10474 12640
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 10468 12600 10517 12628
rect 10468 12588 10474 12600
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 10505 12591 10563 12597
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 10980 12628 11008 12659
rect 10652 12600 11008 12628
rect 10652 12588 10658 12600
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11761 12628 11789 12736
rect 12472 12733 12484 12736
rect 12518 12764 12530 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12518 12736 12909 12764
rect 12518 12733 12530 12736
rect 12472 12727 12530 12733
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 13906 12764 13912 12776
rect 13867 12736 13912 12764
rect 12897 12727 12955 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14148 12736 14274 12764
rect 14148 12724 14154 12736
rect 14246 12705 14274 12736
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 15286 12764 15292 12776
rect 14424 12736 15292 12764
rect 14424 12724 14430 12736
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15381 12767 15439 12773
rect 15381 12733 15393 12767
rect 15427 12764 15439 12767
rect 15562 12764 15568 12776
rect 15427 12736 15568 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15562 12724 15568 12736
rect 15620 12764 15626 12776
rect 16868 12764 16896 12804
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 15620 12736 16896 12764
rect 19889 12767 19947 12773
rect 15620 12724 15626 12736
rect 19889 12733 19901 12767
rect 19935 12733 19947 12767
rect 20162 12764 20168 12776
rect 20123 12736 20168 12764
rect 19889 12727 19947 12733
rect 14231 12699 14289 12705
rect 14231 12665 14243 12699
rect 14277 12665 14289 12699
rect 14231 12659 14289 12665
rect 14918 12656 14924 12708
rect 14976 12696 14982 12708
rect 16022 12705 16028 12708
rect 16019 12696 16028 12705
rect 14976 12668 15469 12696
rect 15983 12668 16028 12696
rect 14976 12656 14982 12668
rect 11882 12628 11888 12640
rect 11480 12600 11789 12628
rect 11843 12600 11888 12628
rect 11480 12588 11486 12600
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 12575 12631 12633 12637
rect 12575 12628 12587 12631
rect 12400 12600 12587 12628
rect 12400 12588 12406 12600
rect 12575 12597 12587 12600
rect 12621 12597 12633 12631
rect 12575 12591 12633 12597
rect 13357 12631 13415 12637
rect 13357 12597 13369 12631
rect 13403 12628 13415 12631
rect 14090 12628 14096 12640
rect 13403 12600 14096 12628
rect 13403 12597 13415 12600
rect 13357 12591 13415 12597
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 15441 12628 15469 12668
rect 16019 12659 16028 12668
rect 16022 12656 16028 12659
rect 16080 12656 16086 12708
rect 17862 12656 17868 12708
rect 17920 12696 17926 12708
rect 18141 12699 18199 12705
rect 18141 12696 18153 12699
rect 17920 12668 18153 12696
rect 17920 12656 17926 12668
rect 18141 12665 18153 12668
rect 18187 12665 18199 12699
rect 18141 12659 18199 12665
rect 18233 12699 18291 12705
rect 18233 12665 18245 12699
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 19153 12699 19211 12705
rect 19153 12665 19165 12699
rect 19199 12696 19211 12699
rect 19242 12696 19248 12708
rect 19199 12668 19248 12696
rect 19199 12665 19211 12668
rect 19153 12659 19211 12665
rect 16574 12628 16580 12640
rect 15441 12600 16580 12628
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 16724 12600 16865 12628
rect 16724 12588 16730 12600
rect 16853 12597 16865 12600
rect 16899 12628 16911 12631
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 16899 12600 17785 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17773 12597 17785 12600
rect 17819 12628 17831 12631
rect 18248 12628 18276 12659
rect 19242 12656 19248 12668
rect 19300 12696 19306 12708
rect 19904 12696 19932 12727
rect 20162 12724 20168 12736
rect 20220 12724 20226 12776
rect 20530 12724 20536 12776
rect 20588 12764 20594 12776
rect 21177 12767 21235 12773
rect 21177 12764 21189 12767
rect 20588 12736 21189 12764
rect 20588 12724 20594 12736
rect 21177 12733 21189 12736
rect 21223 12764 21235 12767
rect 21729 12767 21787 12773
rect 21729 12764 21741 12767
rect 21223 12736 21741 12764
rect 21223 12733 21235 12736
rect 21177 12727 21235 12733
rect 21729 12733 21741 12736
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 20714 12696 20720 12708
rect 19300 12668 20720 12696
rect 19300 12656 19306 12668
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 17819 12600 18276 12628
rect 17819 12597 17831 12600
rect 17773 12591 17831 12597
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 19705 12631 19763 12637
rect 19705 12628 19717 12631
rect 18748 12600 19717 12628
rect 18748 12588 18754 12600
rect 19705 12597 19717 12600
rect 19751 12597 19763 12631
rect 19705 12591 19763 12597
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 937 12427 995 12433
rect 937 12393 949 12427
rect 983 12424 995 12427
rect 1627 12427 1685 12433
rect 1627 12424 1639 12427
rect 983 12396 1639 12424
rect 983 12393 995 12396
rect 937 12387 995 12393
rect 1627 12393 1639 12396
rect 1673 12393 1685 12427
rect 1627 12387 1685 12393
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2639 12427 2697 12433
rect 2639 12393 2651 12427
rect 2685 12424 2697 12427
rect 3234 12424 3240 12436
rect 2685 12396 3240 12424
rect 2685 12393 2697 12396
rect 2639 12387 2697 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 6512 12396 7205 12424
rect 6512 12384 6518 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 7653 12427 7711 12433
rect 7653 12393 7665 12427
rect 7699 12424 7711 12427
rect 8018 12424 8024 12436
rect 7699 12396 8024 12424
rect 7699 12393 7711 12396
rect 7653 12387 7711 12393
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 8570 12424 8576 12436
rect 8220 12396 8576 12424
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 4154 12356 4160 12368
rect 2924 12328 4160 12356
rect 2924 12316 2930 12328
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4249 12359 4307 12365
rect 4249 12325 4261 12359
rect 4295 12356 4307 12359
rect 5994 12356 6000 12368
rect 4295 12328 6000 12356
rect 4295 12325 4307 12328
rect 4249 12319 4307 12325
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 6270 12356 6276 12368
rect 6231 12328 6276 12356
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 6365 12359 6423 12365
rect 6365 12325 6377 12359
rect 6411 12356 6423 12359
rect 7006 12356 7012 12368
rect 6411 12328 7012 12356
rect 6411 12325 6423 12328
rect 6365 12319 6423 12325
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 7742 12356 7748 12368
rect 7064 12328 7748 12356
rect 7064 12316 7070 12328
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 8220 12365 8248 12396
rect 8570 12384 8576 12396
rect 8628 12424 8634 12436
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 8628 12396 11345 12424
rect 8628 12384 8634 12396
rect 11333 12393 11345 12396
rect 11379 12393 11391 12427
rect 11698 12424 11704 12436
rect 11659 12396 11704 12424
rect 11333 12387 11391 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12170 12396 12541 12424
rect 8205 12359 8263 12365
rect 8205 12325 8217 12359
rect 8251 12325 8263 12359
rect 8205 12319 8263 12325
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 9858 12356 9864 12368
rect 8803 12328 9864 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 12170 12356 12198 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 13446 12424 13452 12436
rect 12529 12387 12587 12393
rect 12636 12396 13124 12424
rect 13407 12396 13452 12424
rect 12636 12356 12664 12396
rect 12986 12356 12992 12368
rect 9968 12328 12664 12356
rect 12912 12328 12992 12356
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1524 12291 1582 12297
rect 1524 12288 1536 12291
rect 1452 12260 1536 12288
rect 1452 12248 1458 12260
rect 1524 12257 1536 12260
rect 1570 12257 1582 12291
rect 1524 12251 1582 12257
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2568 12291 2626 12297
rect 2568 12288 2580 12291
rect 2464 12260 2580 12288
rect 2464 12248 2470 12260
rect 2568 12257 2580 12260
rect 2614 12288 2626 12291
rect 3142 12288 3148 12300
rect 2614 12260 3148 12288
rect 2614 12257 2626 12260
rect 2568 12251 2626 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 7101 12291 7159 12297
rect 4856 12260 6107 12288
rect 4856 12248 4862 12260
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4338 12220 4344 12232
rect 4212 12192 4344 12220
rect 4212 12180 4218 12192
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4890 12220 4896 12232
rect 4724 12192 4896 12220
rect 2406 12112 2412 12164
rect 2464 12152 2470 12164
rect 2464 12124 3464 12152
rect 2464 12112 2470 12124
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 2188 12056 2329 12084
rect 2188 12044 2194 12056
rect 2317 12053 2329 12056
rect 2363 12053 2375 12087
rect 2317 12047 2375 12053
rect 3053 12087 3111 12093
rect 3053 12053 3065 12087
rect 3099 12084 3111 12087
rect 3234 12084 3240 12096
rect 3099 12056 3240 12084
rect 3099 12053 3111 12056
rect 3053 12047 3111 12053
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3436 12093 3464 12124
rect 3421 12087 3479 12093
rect 3421 12053 3433 12087
rect 3467 12084 3479 12087
rect 3697 12087 3755 12093
rect 3697 12084 3709 12087
rect 3467 12056 3709 12084
rect 3467 12053 3479 12056
rect 3421 12047 3479 12053
rect 3697 12053 3709 12056
rect 3743 12053 3755 12087
rect 3697 12047 3755 12053
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 4246 12084 4252 12096
rect 3936 12056 4252 12084
rect 3936 12044 3942 12056
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4522 12044 4528 12096
rect 4580 12084 4586 12096
rect 4724 12084 4752 12192
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5718 12220 5724 12232
rect 5592 12192 5724 12220
rect 5592 12180 5598 12192
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 6079 12220 6107 12260
rect 7101 12257 7113 12291
rect 7147 12288 7159 12291
rect 7466 12288 7472 12300
rect 7147 12260 7472 12288
rect 7147 12257 7159 12260
rect 7101 12251 7159 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 8938 12248 8944 12300
rect 8996 12288 9002 12300
rect 9968 12288 9996 12328
rect 11054 12288 11060 12300
rect 8996 12260 11060 12288
rect 8996 12248 9002 12260
rect 6270 12220 6276 12232
rect 6079 12192 6276 12220
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 8110 12220 8116 12232
rect 6972 12192 8116 12220
rect 6972 12180 6978 12192
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9030 12220 9036 12232
rect 8444 12192 9036 12220
rect 8444 12180 8450 12192
rect 9030 12180 9036 12192
rect 9088 12220 9094 12232
rect 9968 12220 9996 12260
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 12170 12288 12198 12328
rect 11756 12260 12198 12288
rect 11756 12248 11762 12260
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 12912 12297 12940 12328
rect 12986 12316 12992 12328
rect 13044 12316 13050 12368
rect 13096 12356 13124 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14001 12427 14059 12433
rect 14001 12424 14013 12427
rect 13964 12396 14013 12424
rect 13964 12384 13970 12396
rect 14001 12393 14013 12396
rect 14047 12424 14059 12427
rect 15381 12427 15439 12433
rect 15381 12424 15393 12427
rect 14047 12396 15393 12424
rect 14047 12393 14059 12396
rect 14001 12387 14059 12393
rect 15381 12393 15393 12396
rect 15427 12393 15439 12427
rect 15381 12387 15439 12393
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 16669 12427 16727 12433
rect 16669 12424 16681 12427
rect 16172 12396 16681 12424
rect 16172 12384 16178 12396
rect 16669 12393 16681 12396
rect 16715 12393 16727 12427
rect 16669 12387 16727 12393
rect 17175 12427 17233 12433
rect 17175 12393 17187 12427
rect 17221 12424 17233 12427
rect 18138 12424 18144 12436
rect 17221 12396 18144 12424
rect 17221 12393 17233 12396
rect 17175 12387 17233 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 19751 12427 19809 12433
rect 19751 12424 19763 12427
rect 18380 12396 19763 12424
rect 18380 12384 18386 12396
rect 19751 12393 19763 12396
rect 19797 12393 19809 12427
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 19751 12387 19809 12393
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 20993 12427 21051 12433
rect 20993 12424 21005 12427
rect 20496 12396 21005 12424
rect 20496 12384 20502 12396
rect 20993 12393 21005 12396
rect 21039 12393 21051 12427
rect 20993 12387 21051 12393
rect 14645 12359 14703 12365
rect 14645 12356 14657 12359
rect 13096 12328 14657 12356
rect 14645 12325 14657 12328
rect 14691 12325 14703 12359
rect 14645 12319 14703 12325
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 15562 12356 15568 12368
rect 15068 12328 15568 12356
rect 15068 12316 15074 12328
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 12400 12260 12449 12288
rect 12400 12248 12406 12260
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12257 12955 12291
rect 13722 12288 13728 12300
rect 12897 12251 12955 12257
rect 13004 12260 13728 12288
rect 9088 12192 9996 12220
rect 9088 12180 9094 12192
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10100 12192 10149 12220
rect 10100 12180 10106 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 13004 12220 13032 12260
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 15488 12297 15516 12328
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16393 12359 16451 12365
rect 16393 12325 16405 12359
rect 16439 12356 16451 12359
rect 16758 12356 16764 12368
rect 16439 12328 16764 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 16758 12316 16764 12328
rect 16816 12316 16822 12368
rect 17494 12316 17500 12368
rect 17552 12356 17558 12368
rect 18233 12359 18291 12365
rect 18233 12356 18245 12359
rect 17552 12328 18245 12356
rect 17552 12316 17558 12328
rect 18233 12325 18245 12328
rect 18279 12325 18291 12359
rect 20180 12356 20208 12384
rect 20180 12328 21404 12356
rect 18233 12319 18291 12325
rect 14252 12291 14310 12297
rect 14252 12257 14264 12291
rect 14298 12288 14310 12291
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 14298 12260 14473 12288
rect 14298 12257 14310 12260
rect 14252 12251 14310 12257
rect 14461 12257 14473 12260
rect 14507 12257 14519 12291
rect 14461 12251 14519 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 15930 12288 15936 12300
rect 15887 12260 15936 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 17104 12291 17162 12297
rect 17104 12257 17116 12291
rect 17150 12288 17162 12291
rect 17218 12288 17224 12300
rect 17150 12260 17224 12288
rect 17150 12257 17162 12260
rect 17104 12251 17162 12257
rect 17218 12248 17224 12260
rect 17276 12288 17282 12300
rect 17770 12288 17776 12300
rect 17276 12260 17776 12288
rect 17276 12248 17282 12260
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19648 12291 19706 12297
rect 19648 12288 19660 12291
rect 19484 12260 19660 12288
rect 19484 12248 19490 12260
rect 19648 12257 19660 12260
rect 19694 12257 19706 12291
rect 19648 12251 19706 12257
rect 19794 12248 19800 12300
rect 19852 12288 19858 12300
rect 20806 12288 20812 12300
rect 19852 12260 20812 12288
rect 19852 12248 19858 12260
rect 20806 12248 20812 12260
rect 20864 12288 20870 12300
rect 21376 12297 21404 12328
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20864 12260 20913 12288
rect 20864 12248 20870 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 21361 12291 21419 12297
rect 21361 12257 21373 12291
rect 21407 12288 21419 12291
rect 21450 12288 21456 12300
rect 21407 12260 21456 12288
rect 21407 12257 21419 12260
rect 21361 12251 21419 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 10928 12192 13032 12220
rect 13280 12192 15025 12220
rect 10928 12180 10934 12192
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 5905 12155 5963 12161
rect 5905 12152 5917 12155
rect 4856 12124 5917 12152
rect 4856 12112 4862 12124
rect 5905 12121 5917 12124
rect 5951 12121 5963 12155
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 5905 12115 5963 12121
rect 6999 12124 9413 12152
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 4580 12056 5181 12084
rect 4580 12044 4586 12056
rect 5169 12053 5181 12056
rect 5215 12053 5227 12087
rect 5534 12084 5540 12096
rect 5495 12056 5540 12084
rect 5169 12047 5227 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6999 12084 7027 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 11330 12112 11336 12164
rect 11388 12152 11394 12164
rect 13280 12152 13308 12192
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17586 12220 17592 12232
rect 17460 12192 17592 12220
rect 17460 12180 17466 12192
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12220 18199 12223
rect 19061 12223 19119 12229
rect 19061 12220 19073 12223
rect 18187 12192 19073 12220
rect 18187 12189 18199 12192
rect 18141 12183 18199 12189
rect 19061 12189 19073 12192
rect 19107 12189 19119 12223
rect 19061 12183 19119 12189
rect 11388 12124 13308 12152
rect 11388 12112 11394 12124
rect 13630 12112 13636 12164
rect 13688 12152 13694 12164
rect 13906 12152 13912 12164
rect 13688 12124 13912 12152
rect 13688 12112 13694 12124
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 14323 12155 14381 12161
rect 14323 12121 14335 12155
rect 14369 12152 14381 12155
rect 18156 12152 18184 12183
rect 14369 12124 18184 12152
rect 14369 12121 14381 12124
rect 14323 12115 14381 12121
rect 18506 12112 18512 12164
rect 18564 12152 18570 12164
rect 18693 12155 18751 12161
rect 18693 12152 18705 12155
rect 18564 12124 18705 12152
rect 18564 12112 18570 12124
rect 18693 12121 18705 12124
rect 18739 12152 18751 12155
rect 19429 12155 19487 12161
rect 19429 12152 19441 12155
rect 18739 12124 19441 12152
rect 18739 12121 18751 12124
rect 18693 12115 18751 12121
rect 19429 12121 19441 12124
rect 19475 12121 19487 12155
rect 19429 12115 19487 12121
rect 6788 12056 7027 12084
rect 6788 12044 6794 12056
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 7800 12056 9045 12084
rect 7800 12044 7806 12056
rect 9033 12053 9045 12056
rect 9079 12084 9091 12087
rect 9306 12084 9312 12096
rect 9079 12056 9312 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9950 12084 9956 12096
rect 9863 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12084 10014 12096
rect 10686 12084 10692 12096
rect 10008 12056 10692 12084
rect 10008 12044 10014 12056
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11054 12084 11060 12096
rect 11015 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11204 12056 12081 12084
rect 11204 12044 11210 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 14461 12087 14519 12093
rect 14461 12053 14473 12087
rect 14507 12084 14519 12087
rect 14642 12084 14648 12096
rect 14507 12056 14648 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 17586 12084 17592 12096
rect 17547 12056 17592 12084
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 17862 12084 17868 12096
rect 17823 12056 17868 12084
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 19576 12056 20453 12084
rect 19576 12044 19582 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 21634 12044 21640 12096
rect 21692 12084 21698 12096
rect 21913 12087 21971 12093
rect 21913 12084 21925 12087
rect 21692 12056 21925 12084
rect 21692 12044 21698 12056
rect 21913 12053 21925 12056
rect 21959 12053 21971 12087
rect 22278 12084 22284 12096
rect 22239 12056 22284 12084
rect 21913 12047 21971 12053
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4154 11880 4160 11892
rect 4028 11852 4160 11880
rect 4028 11840 4034 11852
rect 4154 11840 4160 11852
rect 4212 11880 4218 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 4212 11852 6193 11880
rect 4212 11840 4218 11852
rect 6181 11849 6193 11852
rect 6227 11849 6239 11883
rect 6181 11843 6239 11849
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6914 11880 6920 11892
rect 6328 11852 6920 11880
rect 6328 11840 6334 11852
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8110 11880 8116 11892
rect 8071 11852 8116 11880
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 9490 11880 9496 11892
rect 9451 11852 9496 11880
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 14001 11883 14059 11889
rect 14001 11880 14013 11883
rect 11940 11852 14013 11880
rect 11940 11840 11946 11852
rect 14001 11849 14013 11852
rect 14047 11849 14059 11883
rect 14182 11880 14188 11892
rect 14001 11843 14059 11849
rect 14108 11852 14188 11880
rect 14 11772 20 11824
rect 72 11812 78 11824
rect 5445 11815 5503 11821
rect 5445 11812 5457 11815
rect 72 11784 5457 11812
rect 72 11772 78 11784
rect 5445 11781 5457 11784
rect 5491 11781 5503 11815
rect 5445 11775 5503 11781
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 7926 11812 7932 11824
rect 6420 11784 7932 11812
rect 6420 11772 6426 11784
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 12342 11772 12348 11824
rect 12400 11812 12406 11824
rect 14108 11812 14136 11852
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15059 11883 15117 11889
rect 15059 11849 15071 11883
rect 15105 11880 15117 11883
rect 16482 11880 16488 11892
rect 15105 11852 16488 11880
rect 15105 11849 15117 11852
rect 15059 11843 15117 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17552 11852 17785 11880
rect 17552 11840 17558 11852
rect 17773 11849 17785 11852
rect 17819 11880 17831 11883
rect 18230 11880 18236 11892
rect 17819 11852 18236 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 18230 11840 18236 11852
rect 18288 11880 18294 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 18288 11852 19073 11880
rect 18288 11840 18294 11852
rect 19061 11849 19073 11852
rect 19107 11849 19119 11883
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19061 11843 19119 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 19610 11840 19616 11892
rect 19668 11880 19674 11892
rect 19668 11852 20760 11880
rect 19668 11840 19674 11852
rect 16853 11815 16911 11821
rect 12400 11784 14136 11812
rect 14200 11784 16298 11812
rect 12400 11772 12406 11784
rect 198 11704 204 11756
rect 256 11744 262 11756
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 256 11716 1961 11744
rect 256 11704 262 11716
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 1964 11676 1992 11707
rect 2590 11704 2596 11756
rect 2648 11744 2654 11756
rect 4522 11744 4528 11756
rect 2648 11716 4528 11744
rect 2648 11704 2654 11716
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 6454 11744 6460 11756
rect 5137 11716 6460 11744
rect 1964 11648 3556 11676
rect 934 11568 940 11620
rect 992 11608 998 11620
rect 1394 11608 1400 11620
rect 992 11580 1400 11608
rect 992 11568 998 11580
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 2270 11611 2328 11617
rect 2270 11577 2282 11611
rect 2316 11577 2328 11611
rect 3528 11608 3556 11648
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3732 11679 3790 11685
rect 3732 11676 3744 11679
rect 3660 11648 3744 11676
rect 3660 11636 3666 11648
rect 3732 11645 3744 11648
rect 3778 11676 3790 11679
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 3778 11648 4169 11676
rect 3778 11645 3790 11648
rect 3732 11639 3790 11645
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 5137 11676 5165 11716
rect 6454 11704 6460 11716
rect 6512 11744 6518 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6512 11716 6561 11744
rect 6512 11704 6518 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 4396 11648 5165 11676
rect 5261 11679 5319 11685
rect 4396 11636 4402 11648
rect 5261 11645 5273 11679
rect 5307 11676 5319 11679
rect 5442 11676 5448 11688
rect 5307 11648 5448 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 5442 11636 5448 11648
rect 5500 11676 5506 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5500 11648 5825 11676
rect 5500 11636 5506 11648
rect 5813 11645 5825 11648
rect 5859 11645 5871 11679
rect 5813 11639 5871 11645
rect 3528 11580 4016 11608
rect 2270 11571 2328 11577
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11540 1826 11552
rect 2285 11540 2313 11571
rect 2866 11540 2872 11552
rect 1820 11512 2313 11540
rect 2827 11512 2872 11540
rect 1820 11500 1826 11512
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3142 11540 3148 11552
rect 3103 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3878 11549 3884 11552
rect 3835 11543 3884 11549
rect 3835 11540 3847 11543
rect 3660 11512 3847 11540
rect 3660 11500 3666 11512
rect 3835 11509 3847 11512
rect 3881 11509 3884 11543
rect 3835 11503 3884 11509
rect 3878 11500 3884 11503
rect 3936 11500 3942 11552
rect 3988 11540 4016 11580
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 4525 11611 4583 11617
rect 4525 11608 4537 11611
rect 4120 11580 4537 11608
rect 4120 11568 4126 11580
rect 4525 11577 4537 11580
rect 4571 11577 4583 11611
rect 4890 11608 4896 11620
rect 4851 11580 4896 11608
rect 4525 11571 4583 11577
rect 4890 11568 4896 11580
rect 4948 11568 4954 11620
rect 6564 11608 6592 11707
rect 6730 11704 6736 11756
rect 6788 11744 6794 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6788 11716 6837 11744
rect 6788 11704 6794 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8846 11744 8852 11756
rect 8619 11716 8852 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 9861 11747 9919 11753
rect 9861 11744 9873 11747
rect 9824 11716 9873 11744
rect 9824 11704 9830 11716
rect 9861 11713 9873 11716
rect 9907 11744 9919 11747
rect 12253 11747 12311 11753
rect 9907 11716 11192 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 8909 11648 10149 11676
rect 8909 11617 8937 11648
rect 10137 11645 10149 11648
rect 10183 11676 10195 11679
rect 10410 11676 10416 11688
rect 10183 11648 10416 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10870 11676 10876 11688
rect 10831 11648 10876 11676
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 11164 11685 11192 11716
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12802 11744 12808 11756
rect 12299 11716 12808 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13446 11744 13452 11756
rect 13127 11716 13452 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11645 11207 11679
rect 11149 11639 11207 11645
rect 7146 11611 7204 11617
rect 7146 11608 7158 11611
rect 6564 11580 7158 11608
rect 7146 11577 7158 11580
rect 7192 11608 7204 11611
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 7192 11580 8217 11608
rect 7192 11577 7204 11580
rect 7146 11571 7204 11577
rect 8205 11577 8217 11580
rect 8251 11608 8263 11611
rect 8389 11611 8447 11617
rect 8389 11608 8401 11611
rect 8251 11580 8401 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8389 11577 8401 11580
rect 8435 11608 8447 11611
rect 8894 11611 8952 11617
rect 8894 11608 8906 11611
rect 8435 11580 8906 11608
rect 8435 11577 8447 11580
rect 8389 11571 8447 11577
rect 8894 11577 8906 11580
rect 8940 11577 8952 11611
rect 10318 11608 10324 11620
rect 8894 11571 8952 11577
rect 9692 11580 10324 11608
rect 4798 11540 4804 11552
rect 3988 11512 4804 11540
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6270 11540 6276 11552
rect 5960 11512 6276 11540
rect 5960 11500 5966 11512
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9692 11540 9720 11580
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 11164 11608 11192 11639
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 14200 11676 14228 11784
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 14884 11716 15393 11744
rect 14884 11704 14890 11716
rect 15003 11685 15031 11716
rect 15381 11713 15393 11716
rect 15427 11744 15439 11747
rect 15562 11744 15568 11756
rect 15427 11716 15568 11744
rect 15427 11713 15439 11716
rect 15381 11707 15439 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16114 11744 16120 11756
rect 15979 11716 16120 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16270 11744 16298 11784
rect 16853 11781 16865 11815
rect 16899 11812 16911 11815
rect 19794 11812 19800 11824
rect 16899 11784 19800 11812
rect 16899 11781 16911 11784
rect 16853 11775 16911 11781
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 18414 11744 18420 11756
rect 16270 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 18782 11744 18788 11756
rect 18743 11716 18788 11744
rect 18782 11704 18788 11716
rect 18840 11744 18846 11756
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 18840 11716 19717 11744
rect 18840 11704 18846 11716
rect 19705 11713 19717 11716
rect 19751 11744 19763 11747
rect 20162 11744 20168 11756
rect 19751 11716 20168 11744
rect 19751 11713 19763 11716
rect 19705 11707 19763 11713
rect 20162 11704 20168 11716
rect 20220 11704 20226 11756
rect 20732 11744 20760 11852
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20864 11852 20913 11880
rect 20864 11840 20870 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 21358 11880 21364 11892
rect 21319 11852 21364 11880
rect 20901 11843 20959 11849
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 21726 11840 21732 11892
rect 21784 11880 21790 11892
rect 22097 11883 22155 11889
rect 22097 11880 22109 11883
rect 21784 11852 22109 11880
rect 21784 11840 21790 11852
rect 22097 11849 22109 11852
rect 22143 11849 22155 11883
rect 22097 11843 22155 11849
rect 21450 11772 21456 11824
rect 21508 11812 21514 11824
rect 21821 11815 21879 11821
rect 21821 11812 21833 11815
rect 21508 11784 21833 11812
rect 21508 11772 21514 11784
rect 21821 11781 21833 11784
rect 21867 11781 21879 11815
rect 21821 11775 21879 11781
rect 21358 11744 21364 11756
rect 20732 11716 21364 11744
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 14988 11679 15046 11685
rect 14988 11676 15000 11679
rect 11940 11648 14228 11676
rect 14966 11648 15000 11676
rect 11940 11636 11946 11648
rect 14988 11645 15000 11648
rect 15034 11645 15046 11679
rect 17218 11676 17224 11688
rect 17179 11648 17224 11676
rect 14988 11639 15046 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 21177 11679 21235 11685
rect 21177 11645 21189 11679
rect 21223 11676 21235 11679
rect 21726 11676 21732 11688
rect 21223 11648 21732 11676
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 21726 11636 21732 11648
rect 21784 11636 21790 11688
rect 13078 11608 13084 11620
rect 11164 11580 13084 11608
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 13443 11611 13501 11617
rect 13443 11577 13455 11611
rect 13489 11608 13501 11611
rect 14090 11608 14096 11620
rect 13489 11580 14096 11608
rect 13489 11577 13501 11580
rect 13443 11571 13501 11577
rect 13648 11552 13676 11580
rect 14090 11568 14096 11580
rect 14148 11608 14154 11620
rect 15749 11611 15807 11617
rect 15749 11608 15761 11611
rect 14148 11580 15761 11608
rect 14148 11568 14154 11580
rect 15749 11577 15761 11580
rect 15795 11608 15807 11611
rect 16114 11608 16120 11620
rect 15795 11580 16120 11608
rect 15795 11577 15807 11580
rect 15749 11571 15807 11577
rect 16114 11568 16120 11580
rect 16172 11608 16178 11620
rect 16254 11611 16312 11617
rect 16254 11608 16266 11611
rect 16172 11580 16266 11608
rect 16172 11568 16178 11580
rect 16254 11577 16266 11580
rect 16300 11577 16312 11611
rect 16254 11571 16312 11577
rect 17586 11568 17592 11620
rect 17644 11608 17650 11620
rect 18138 11608 18144 11620
rect 17644 11580 18144 11608
rect 17644 11568 17650 11580
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 18288 11580 18333 11608
rect 18288 11568 18294 11580
rect 19794 11568 19800 11620
rect 19852 11608 19858 11620
rect 20349 11611 20407 11617
rect 19852 11580 19897 11608
rect 19852 11568 19858 11580
rect 20349 11577 20361 11611
rect 20395 11577 20407 11611
rect 20349 11571 20407 11577
rect 10686 11540 10692 11552
rect 8536 11512 9720 11540
rect 10647 11512 10692 11540
rect 8536 11500 8542 11512
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12434 11540 12440 11552
rect 11931 11512 12440 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 12989 11543 13047 11549
rect 12989 11509 13001 11543
rect 13035 11540 13047 11543
rect 13630 11540 13636 11552
rect 13035 11512 13636 11540
rect 13035 11509 13047 11512
rect 12989 11503 13047 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 14369 11543 14427 11549
rect 14369 11509 14381 11543
rect 14415 11540 14427 11543
rect 14642 11540 14648 11552
rect 14415 11512 14648 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 14829 11543 14887 11549
rect 14829 11509 14841 11543
rect 14875 11540 14887 11543
rect 15010 11540 15016 11552
rect 14875 11512 15016 11540
rect 14875 11509 14887 11512
rect 14829 11503 14887 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 20364 11540 20392 11571
rect 18656 11512 20392 11540
rect 18656 11500 18662 11512
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 17 11339 75 11345
rect 17 11305 29 11339
rect 63 11336 75 11339
rect 842 11336 848 11348
rect 63 11308 848 11336
rect 63 11305 75 11308
rect 17 11299 75 11305
rect 842 11296 848 11308
rect 900 11296 906 11348
rect 3510 11336 3516 11348
rect 2884 11308 3516 11336
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 2546 11271 2604 11277
rect 2546 11268 2558 11271
rect 1820 11240 2558 11268
rect 1820 11228 1826 11240
rect 2546 11237 2558 11240
rect 2592 11237 2604 11271
rect 2546 11231 2604 11237
rect 198 11160 204 11212
rect 256 11200 262 11212
rect 2884 11200 2912 11308
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4338 11336 4344 11348
rect 3936 11308 4344 11336
rect 3936 11296 3942 11308
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 4948 11308 5641 11336
rect 4948 11296 4954 11308
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 5629 11299 5687 11305
rect 5828 11308 7113 11336
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 4249 11271 4307 11277
rect 4249 11268 4261 11271
rect 4120 11240 4261 11268
rect 4120 11228 4126 11240
rect 4249 11237 4261 11240
rect 4295 11237 4307 11271
rect 5828 11268 5856 11308
rect 7101 11305 7113 11308
rect 7147 11305 7159 11339
rect 7101 11299 7159 11305
rect 7190 11296 7196 11348
rect 7248 11296 7254 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 7742 11336 7748 11348
rect 7699 11308 7748 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8628 11308 8769 11336
rect 8628 11296 8634 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 9364 11308 9413 11336
rect 9364 11296 9370 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9858 11336 9864 11348
rect 9819 11308 9864 11336
rect 9401 11299 9459 11305
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 10689 11339 10747 11345
rect 10689 11305 10701 11339
rect 10735 11336 10747 11339
rect 10870 11336 10876 11348
rect 10735 11308 10876 11336
rect 10735 11305 10747 11308
rect 10689 11299 10747 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11974 11336 11980 11348
rect 10980 11308 11980 11336
rect 4249 11231 4307 11237
rect 4310 11240 5856 11268
rect 4310 11212 4338 11240
rect 5902 11228 5908 11280
rect 5960 11268 5966 11280
rect 5997 11271 6055 11277
rect 5997 11268 6009 11271
rect 5960 11240 6009 11268
rect 5960 11228 5966 11240
rect 5997 11237 6009 11240
rect 6043 11268 6055 11271
rect 6546 11268 6552 11280
rect 6043 11240 6552 11268
rect 6043 11237 6055 11240
rect 5997 11231 6055 11237
rect 6546 11228 6552 11240
rect 6604 11228 6610 11280
rect 256 11172 2912 11200
rect 3145 11203 3203 11209
rect 256 11160 262 11172
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 4310 11200 4344 11212
rect 3191 11172 4344 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 4338 11160 4344 11172
rect 4396 11200 4402 11212
rect 5258 11200 5264 11212
rect 4396 11172 5264 11200
rect 4396 11160 4402 11172
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 4246 11132 4252 11144
rect 2271 11104 4252 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 3513 11067 3571 11073
rect 3513 11033 3525 11067
rect 3559 11064 3571 11067
rect 4448 11064 4476 11172
rect 4632 11141 4660 11172
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5905 11135 5963 11141
rect 4764 11104 4809 11132
rect 4764 11092 4770 11104
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 7208 11132 7236 11296
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9214 11268 9220 11280
rect 9088 11240 9220 11268
rect 9088 11228 9094 11240
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 10980 11268 11008 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12066 11296 12072 11348
rect 12124 11296 12130 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 13446 11336 13452 11348
rect 13136 11308 13452 11336
rect 13136 11296 13142 11308
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 14231 11339 14289 11345
rect 14231 11336 14243 11339
rect 13780 11308 14243 11336
rect 13780 11296 13786 11308
rect 14231 11305 14243 11308
rect 14277 11305 14289 11339
rect 14918 11336 14924 11348
rect 14879 11308 14924 11336
rect 14231 11299 14289 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16114 11336 16120 11348
rect 16075 11308 16120 11336
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16666 11336 16672 11348
rect 16627 11308 16672 11336
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 17635 11339 17693 11345
rect 17635 11305 17647 11339
rect 17681 11336 17693 11339
rect 17862 11336 17868 11348
rect 17681 11308 17868 11336
rect 17681 11305 17693 11308
rect 17635 11299 17693 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 19705 11339 19763 11345
rect 19705 11305 19717 11339
rect 19751 11336 19763 11339
rect 19794 11336 19800 11348
rect 19751 11308 19800 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 20162 11296 20168 11348
rect 20220 11336 20226 11348
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 20220 11308 20361 11336
rect 20220 11296 20226 11308
rect 20349 11305 20361 11308
rect 20395 11305 20407 11339
rect 20349 11299 20407 11305
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20680 11308 21005 11336
rect 20680 11296 20686 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 10842 11240 11008 11268
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 8904 11172 9689 11200
rect 8904 11160 8910 11172
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 10410 11200 10416 11212
rect 9723 11172 10416 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 7742 11132 7748 11144
rect 5951 11104 7748 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 10842 11132 10870 11240
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 11149 11271 11207 11277
rect 11149 11268 11161 11271
rect 11112 11240 11161 11268
rect 11112 11228 11118 11240
rect 11149 11237 11161 11240
rect 11195 11237 11207 11271
rect 11149 11231 11207 11237
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11200 11759 11203
rect 12084 11200 12112 11296
rect 12618 11268 12624 11280
rect 12579 11240 12624 11268
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 12713 11271 12771 11277
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 12802 11268 12808 11280
rect 12759 11240 12808 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 12952 11240 13308 11268
rect 12952 11228 12958 11240
rect 11747 11172 12112 11200
rect 13280 11200 13308 11240
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 14553 11271 14611 11277
rect 14553 11268 14565 11271
rect 13412 11240 14565 11268
rect 13412 11228 13418 11240
rect 14553 11237 14565 11240
rect 14599 11237 14611 11271
rect 14553 11231 14611 11237
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 18693 11271 18751 11277
rect 18693 11268 18705 11271
rect 17828 11240 18705 11268
rect 17828 11228 17834 11240
rect 18693 11237 18705 11240
rect 18739 11268 18751 11271
rect 18874 11268 18880 11280
rect 18739 11240 18880 11268
rect 18739 11237 18751 11240
rect 18693 11231 18751 11237
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 19886 11228 19892 11280
rect 19944 11268 19950 11280
rect 19944 11240 21404 11268
rect 19944 11228 19950 11240
rect 14090 11200 14096 11212
rect 13280 11172 14096 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 15746 11200 15752 11212
rect 15707 11172 15752 11200
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11200 17555 11203
rect 17586 11200 17592 11212
rect 17543 11172 17592 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 21376 11209 21404 11240
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20864 11172 20913 11200
rect 20864 11160 20870 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 21361 11203 21419 11209
rect 21361 11169 21373 11203
rect 21407 11200 21419 11203
rect 21726 11200 21732 11212
rect 21407 11172 21732 11200
rect 21407 11169 21419 11172
rect 21361 11163 21419 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 7883 11104 10870 11132
rect 11057 11135 11115 11141
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 11057 11101 11069 11135
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 3559 11036 4476 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 4522 11024 4528 11076
rect 4580 11064 4586 11076
rect 4798 11064 4804 11076
rect 4580 11036 4804 11064
rect 4580 11024 4586 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5258 11064 5264 11076
rect 5219 11036 5264 11064
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 6457 11067 6515 11073
rect 6457 11033 6469 11067
rect 6503 11064 6515 11067
rect 6730 11064 6736 11076
rect 6503 11036 6736 11064
rect 6503 11033 6515 11036
rect 6457 11027 6515 11033
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 7984 11036 10548 11064
rect 7984 11024 7990 11036
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 1762 10996 1768 11008
rect 1719 10968 1768 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 1762 10956 1768 10968
rect 1820 10996 1826 11008
rect 1949 10999 2007 11005
rect 1949 10996 1961 10999
rect 1820 10968 1961 10996
rect 1820 10956 1826 10968
rect 1949 10965 1961 10968
rect 1995 10965 2007 10999
rect 1949 10959 2007 10965
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 3881 10999 3939 11005
rect 3881 10996 3893 10999
rect 3752 10968 3893 10996
rect 3752 10956 3758 10968
rect 3881 10965 3893 10968
rect 3927 10996 3939 10999
rect 4387 10999 4445 11005
rect 4387 10996 4399 10999
rect 3927 10968 4399 10996
rect 3927 10965 3939 10968
rect 3881 10959 3939 10965
rect 4172 10928 4200 10968
rect 4387 10965 4399 10968
rect 4433 10965 4445 10999
rect 4387 10959 4445 10965
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 6825 10999 6883 11005
rect 6825 10996 6837 10999
rect 5776 10968 6837 10996
rect 5776 10956 5782 10968
rect 6825 10965 6837 10968
rect 6871 10965 6883 10999
rect 7098 10996 7104 11008
rect 7011 10968 7104 10996
rect 6825 10959 6883 10965
rect 7098 10956 7104 10968
rect 7156 10996 7162 11008
rect 7285 10999 7343 11005
rect 7285 10996 7297 10999
rect 7156 10968 7297 10996
rect 7156 10956 7162 10968
rect 7285 10965 7297 10968
rect 7331 10996 7343 10999
rect 8110 10996 8116 11008
rect 7331 10968 8116 10996
rect 7331 10965 7343 10968
rect 7285 10959 7343 10965
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 9030 10996 9036 11008
rect 8991 10968 9036 10996
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9490 10996 9496 11008
rect 9364 10968 9496 10996
rect 9364 10956 9370 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 10042 10956 10048 11008
rect 10100 10996 10106 11008
rect 10229 10999 10287 11005
rect 10229 10996 10241 10999
rect 10100 10968 10241 10996
rect 10100 10956 10106 10968
rect 10229 10965 10241 10968
rect 10275 10965 10287 10999
rect 10520 10996 10548 11036
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 11072 11064 11100 11095
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13320 11104 13553 11132
rect 13320 11092 13326 11104
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 15344 11104 15485 11132
rect 15344 11092 15350 11104
rect 15473 11101 15485 11104
rect 15519 11132 15531 11135
rect 15930 11132 15936 11144
rect 15519 11104 15936 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 18598 11132 18604 11144
rect 18559 11104 18604 11132
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 10928 11036 11100 11064
rect 10928 11024 10934 11036
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 13170 11064 13176 11076
rect 11388 11036 13176 11064
rect 11388 11024 11394 11036
rect 13170 11024 13176 11036
rect 13228 11064 13234 11076
rect 18892 11064 18920 11095
rect 13228 11036 18920 11064
rect 13228 11024 13234 11036
rect 12345 10999 12403 11005
rect 12345 10996 12357 10999
rect 10520 10968 12357 10996
rect 10229 10959 10287 10965
rect 12345 10965 12357 10968
rect 12391 10965 12403 10999
rect 12345 10959 12403 10965
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13909 10999 13967 11005
rect 13909 10996 13921 10999
rect 13412 10968 13921 10996
rect 13412 10956 13418 10968
rect 13909 10965 13921 10968
rect 13955 10965 13967 10999
rect 16942 10996 16948 11008
rect 16903 10968 16948 10996
rect 13909 10959 13967 10965
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17310 10996 17316 11008
rect 17271 10968 17316 10996
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 18141 10999 18199 11005
rect 18141 10965 18153 10999
rect 18187 10996 18199 10999
rect 18230 10996 18236 11008
rect 18187 10968 18236 10996
rect 18187 10965 18199 10968
rect 18141 10959 18199 10965
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 19981 10999 20039 11005
rect 19981 10996 19993 10999
rect 18656 10968 19993 10996
rect 18656 10956 18662 10968
rect 19981 10965 19993 10968
rect 20027 10965 20039 10999
rect 19981 10959 20039 10965
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 21913 10999 21971 11005
rect 21913 10996 21925 10999
rect 20772 10968 21925 10996
rect 20772 10956 20778 10968
rect 21913 10965 21925 10968
rect 21959 10965 21971 10999
rect 22278 10996 22284 11008
rect 22239 10968 22284 10996
rect 21913 10959 21971 10965
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 4172 10804 4200 10832
rect 1210 10752 1216 10804
rect 1268 10792 1274 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1268 10764 1593 10792
rect 1268 10752 1274 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2682 10792 2688 10804
rect 2455 10764 2688 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2516 10597 2544 10764
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 4154 10752 4160 10804
rect 4212 10752 4218 10804
rect 4338 10792 4344 10804
rect 4299 10764 4344 10792
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 5902 10792 5908 10804
rect 5767 10764 5908 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8754 10792 8760 10804
rect 7800 10764 8760 10792
rect 7800 10752 7806 10764
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 9398 10792 9404 10804
rect 9263 10764 9404 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11112 10764 11345 10792
rect 11112 10752 11118 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 11974 10792 11980 10804
rect 11756 10764 11980 10792
rect 11756 10752 11762 10764
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 13354 10752 13360 10804
rect 13412 10792 13418 10804
rect 13906 10792 13912 10804
rect 13412 10764 13912 10792
rect 13412 10752 13418 10764
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14090 10792 14096 10804
rect 14051 10764 14096 10792
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 15841 10795 15899 10801
rect 15841 10761 15853 10795
rect 15887 10792 15899 10795
rect 16114 10792 16120 10804
rect 15887 10764 16120 10792
rect 15887 10761 15899 10764
rect 15841 10755 15899 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 17586 10792 17592 10804
rect 17499 10764 17592 10792
rect 17586 10752 17592 10764
rect 17644 10792 17650 10804
rect 18322 10792 18328 10804
rect 17644 10764 18328 10792
rect 17644 10752 17650 10764
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 19061 10795 19119 10801
rect 19061 10792 19073 10795
rect 18932 10764 19073 10792
rect 18932 10752 18938 10764
rect 19061 10761 19073 10764
rect 19107 10761 19119 10795
rect 19061 10755 19119 10761
rect 19610 10752 19616 10804
rect 19668 10792 19674 10804
rect 19751 10795 19809 10801
rect 19751 10792 19763 10795
rect 19668 10764 19763 10792
rect 19668 10752 19674 10764
rect 19751 10761 19763 10764
rect 19797 10761 19809 10795
rect 19751 10755 19809 10761
rect 20254 10752 20260 10804
rect 20312 10792 20318 10804
rect 20533 10795 20591 10801
rect 20533 10792 20545 10795
rect 20312 10764 20545 10792
rect 20312 10752 20318 10764
rect 20533 10761 20545 10764
rect 20579 10761 20591 10795
rect 20533 10755 20591 10761
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 4028 10696 6377 10724
rect 4028 10684 4034 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 9030 10724 9036 10736
rect 6365 10687 6423 10693
rect 7024 10696 9036 10724
rect 7024 10656 7052 10696
rect 9030 10684 9036 10696
rect 9088 10684 9094 10736
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 10870 10724 10876 10736
rect 9548 10696 10876 10724
rect 9548 10684 9554 10696
rect 10870 10684 10876 10696
rect 10928 10724 10934 10736
rect 10965 10727 11023 10733
rect 10965 10724 10977 10727
rect 10928 10696 10977 10724
rect 10928 10684 10934 10696
rect 10965 10693 10977 10696
rect 11011 10693 11023 10727
rect 13446 10724 13452 10736
rect 10965 10687 11023 10693
rect 11440 10696 13452 10724
rect 7558 10656 7564 10668
rect 4816 10628 7052 10656
rect 7519 10628 7564 10656
rect 937 10591 995 10597
rect 937 10557 949 10591
rect 983 10588 995 10591
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 983 10560 1409 10588
rect 983 10557 995 10560
rect 937 10551 995 10557
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10557 2559 10591
rect 2501 10551 2559 10557
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10588 2743 10591
rect 2731 10560 3464 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 385 10523 443 10529
rect 385 10489 397 10523
rect 431 10520 443 10523
rect 431 10492 2820 10520
rect 431 10489 443 10492
rect 385 10483 443 10489
rect 2516 10464 2544 10492
rect 1762 10452 1768 10464
rect 1675 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10452 1826 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1820 10424 1961 10452
rect 1820 10412 1826 10424
rect 1949 10421 1961 10424
rect 1995 10421 2007 10455
rect 1949 10415 2007 10421
rect 2498 10412 2504 10464
rect 2556 10412 2562 10464
rect 2792 10461 2820 10492
rect 3436 10464 3464 10560
rect 3878 10548 3884 10600
rect 3936 10548 3942 10600
rect 4522 10548 4528 10600
rect 4580 10588 4586 10600
rect 4816 10597 4844 10628
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 8168 10628 8309 10656
rect 8168 10616 8174 10628
rect 8297 10625 8309 10628
rect 8343 10656 8355 10659
rect 9122 10656 9128 10668
rect 8343 10628 9128 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 9824 10628 9904 10656
rect 9824 10616 9830 10628
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4580 10560 4813 10588
rect 4580 10548 4586 10560
rect 4801 10557 4813 10560
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5442 10588 5448 10600
rect 5132 10560 5448 10588
rect 5132 10548 5138 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8478 10588 8484 10600
rect 8435 10560 8484 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 9398 10588 9404 10600
rect 9359 10560 9404 10588
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 9876 10597 9904 10628
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11440 10656 11468 10696
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 17678 10684 17684 10736
rect 17736 10724 17742 10736
rect 20438 10724 20444 10736
rect 17736 10696 20444 10724
rect 17736 10684 17742 10696
rect 20438 10684 20444 10696
rect 20496 10684 20502 10736
rect 12802 10656 12808 10668
rect 10468 10628 11468 10656
rect 11761 10628 12808 10656
rect 10468 10616 10474 10628
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 10042 10588 10048 10600
rect 10003 10560 10048 10588
rect 9861 10551 9919 10557
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 3896 10520 3924 10548
rect 6917 10523 6975 10529
rect 3712 10492 4752 10520
rect 3712 10464 3740 10492
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10421 2835 10455
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 2777 10415 2835 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3694 10452 3700 10464
rect 3655 10424 3700 10452
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 4338 10452 4344 10464
rect 3936 10424 4344 10452
rect 3936 10412 3942 10424
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4724 10461 4752 10492
rect 6917 10489 6929 10523
rect 6963 10489 6975 10523
rect 6917 10483 6975 10489
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 5166 10452 5172 10464
rect 4755 10424 5172 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 5500 10424 6009 10452
rect 5500 10412 5506 10424
rect 5997 10421 6009 10424
rect 6043 10421 6055 10455
rect 6932 10452 6960 10483
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7064 10492 7109 10520
rect 7064 10480 7070 10492
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 11761 10520 11789 10628
rect 12802 10616 12808 10628
rect 12860 10656 12866 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12860 10628 13553 10656
rect 12860 10616 12866 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 14550 10656 14556 10668
rect 14511 10628 14556 10656
rect 13541 10619 13599 10625
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 14826 10656 14832 10668
rect 14787 10628 14832 10656
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16206 10656 16212 10668
rect 16071 10628 16212 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 18012 10628 18153 10656
rect 18012 10616 18018 10628
rect 18141 10625 18153 10628
rect 18187 10656 18199 10659
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 18187 10628 19441 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 19429 10625 19441 10628
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 15344 10560 16957 10588
rect 15344 10548 15350 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 19648 10591 19706 10597
rect 19648 10588 19660 10591
rect 16945 10551 17003 10557
rect 18892 10560 19660 10588
rect 9824 10492 11789 10520
rect 12253 10523 12311 10529
rect 9824 10480 9830 10492
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12526 10520 12532 10532
rect 12299 10492 12532 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12630 10523 12688 10529
rect 12630 10489 12642 10523
rect 12676 10520 12688 10523
rect 12894 10520 12900 10532
rect 12676 10492 12900 10520
rect 12676 10489 12688 10492
rect 12630 10483 12688 10489
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 13170 10520 13176 10532
rect 13131 10492 13176 10520
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 14642 10480 14648 10532
rect 14700 10520 14706 10532
rect 14700 10492 14745 10520
rect 14700 10480 14706 10492
rect 16114 10480 16120 10532
rect 16172 10520 16178 10532
rect 16346 10523 16404 10529
rect 16346 10520 16358 10523
rect 16172 10492 16358 10520
rect 16172 10480 16178 10492
rect 16346 10489 16358 10492
rect 16392 10520 16404 10523
rect 16574 10520 16580 10532
rect 16392 10492 16580 10520
rect 16392 10489 16404 10492
rect 16346 10483 16404 10489
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 18230 10520 18236 10532
rect 18191 10492 18236 10520
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 18782 10520 18788 10532
rect 18743 10492 18788 10520
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 7742 10452 7748 10464
rect 6932 10424 7748 10452
rect 5997 10415 6055 10421
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 8573 10455 8631 10461
rect 8573 10452 8585 10455
rect 8536 10424 8585 10452
rect 8536 10412 8542 10424
rect 8573 10421 8585 10424
rect 8619 10452 8631 10455
rect 10042 10452 10048 10464
rect 8619 10424 10048 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10870 10452 10876 10464
rect 10459 10424 10876 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 11793 10455 11851 10461
rect 11793 10452 11805 10455
rect 11756 10424 11805 10452
rect 11756 10412 11762 10424
rect 11793 10421 11805 10424
rect 11839 10421 11851 10455
rect 11793 10415 11851 10421
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 18892 10452 18920 10560
rect 19648 10557 19660 10560
rect 19694 10588 19706 10591
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 19694 10560 20085 10588
rect 19694 10557 19706 10560
rect 19648 10551 19706 10557
rect 20073 10557 20085 10560
rect 20119 10557 20131 10591
rect 20548 10588 20576 10755
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20864 10764 20913 10792
rect 20864 10752 20870 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 21726 10792 21732 10804
rect 21687 10764 21732 10792
rect 20901 10755 20959 10761
rect 21726 10752 21732 10764
rect 21784 10752 21790 10804
rect 21361 10727 21419 10733
rect 21361 10693 21373 10727
rect 21407 10724 21419 10727
rect 23474 10724 23480 10736
rect 21407 10696 23480 10724
rect 21407 10693 21419 10696
rect 21361 10687 21419 10693
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 20548 10560 21189 10588
rect 20073 10551 20131 10557
rect 21177 10557 21189 10560
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 20088 10520 20116 10551
rect 20530 10520 20536 10532
rect 20088 10492 20536 10520
rect 20530 10480 20536 10492
rect 20588 10480 20594 10532
rect 22094 10452 22100 10464
rect 17828 10424 18920 10452
rect 22055 10424 22100 10452
rect 17828 10412 17834 10424
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 201 10387 259 10393
rect 201 10353 213 10387
rect 247 10384 259 10387
rect 385 10387 443 10393
rect 385 10384 397 10387
rect 247 10356 397 10384
rect 247 10353 259 10356
rect 201 10347 259 10353
rect 385 10353 397 10356
rect 431 10353 443 10387
rect 385 10347 443 10353
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 1811 10220 2605 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 2593 10217 2605 10220
rect 2639 10248 2651 10251
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2639 10220 2973 10248
rect 2639 10217 2651 10220
rect 2593 10211 2651 10217
rect 2961 10217 2973 10220
rect 3007 10248 3019 10251
rect 3329 10251 3387 10257
rect 3329 10248 3341 10251
rect 3007 10220 3341 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 3329 10217 3341 10220
rect 3375 10248 3387 10251
rect 3694 10248 3700 10260
rect 3375 10220 3700 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4341 10251 4399 10257
rect 4212 10220 4257 10248
rect 4212 10208 4218 10220
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 4614 10248 4620 10260
rect 4387 10220 4620 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 5442 10248 5448 10260
rect 4856 10220 5448 10248
rect 4856 10208 4862 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6546 10248 6552 10260
rect 6144 10220 6552 10248
rect 6144 10208 6150 10220
rect 6546 10208 6552 10220
rect 6604 10248 6610 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 6604 10220 7205 10248
rect 6604 10208 6610 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7739 10251 7797 10257
rect 7739 10248 7751 10251
rect 7193 10211 7251 10217
rect 7392 10220 7751 10248
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 4522 10180 4528 10192
rect 3568 10152 4528 10180
rect 3568 10140 3574 10152
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 5166 10140 5172 10192
rect 5224 10180 5230 10192
rect 5991 10183 6049 10189
rect 5991 10180 6003 10183
rect 5224 10152 6003 10180
rect 5224 10140 5230 10152
rect 5991 10149 6003 10152
rect 6037 10180 6049 10183
rect 7392 10180 7420 10220
rect 7739 10217 7751 10220
rect 7785 10217 7797 10251
rect 7739 10211 7797 10217
rect 7834 10208 7840 10260
rect 7892 10248 7898 10260
rect 9815 10251 9873 10257
rect 9815 10248 9827 10251
rect 7892 10220 9827 10248
rect 7892 10208 7898 10220
rect 9815 10217 9827 10220
rect 9861 10217 9873 10251
rect 9815 10211 9873 10217
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10594 10248 10600 10260
rect 10008 10220 10600 10248
rect 10008 10208 10014 10220
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 11514 10248 11520 10260
rect 11287 10220 11520 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 12253 10251 12311 10257
rect 12253 10217 12265 10251
rect 12299 10248 12311 10251
rect 12434 10248 12440 10260
rect 12299 10220 12440 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13170 10248 13176 10260
rect 12728 10220 13176 10248
rect 6037 10152 7420 10180
rect 6037 10149 6049 10152
rect 5991 10143 6049 10149
rect 8570 10140 8576 10192
rect 8628 10180 8634 10192
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 8628 10152 8953 10180
rect 8628 10140 8634 10152
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 8941 10143 8999 10149
rect 9306 10140 9312 10192
rect 9364 10180 9370 10192
rect 10321 10183 10379 10189
rect 10321 10180 10333 10183
rect 9364 10152 10333 10180
rect 9364 10140 9370 10152
rect 10321 10149 10333 10152
rect 10367 10149 10379 10183
rect 10321 10143 10379 10149
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 12728 10180 12756 10220
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13504 10220 13921 10248
rect 13504 10208 13510 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 14553 10251 14611 10257
rect 14553 10217 14565 10251
rect 14599 10248 14611 10251
rect 14642 10248 14648 10260
rect 14599 10220 14648 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 15746 10248 15752 10260
rect 15703 10220 15752 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16025 10251 16083 10257
rect 16025 10217 16037 10251
rect 16071 10248 16083 10251
rect 16206 10248 16212 10260
rect 16071 10220 16212 10248
rect 16071 10217 16083 10220
rect 16025 10211 16083 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16574 10248 16580 10260
rect 16535 10220 16580 10248
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 16816 10220 17816 10248
rect 16816 10208 16822 10220
rect 11204 10152 12756 10180
rect 11204 10140 11210 10152
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 13034 10183 13092 10189
rect 13034 10180 13046 10183
rect 12860 10152 13046 10180
rect 12860 10140 12866 10152
rect 13034 10149 13046 10152
rect 13080 10180 13092 10183
rect 13630 10180 13636 10192
rect 13080 10152 13636 10180
rect 13080 10149 13092 10152
rect 13034 10143 13092 10149
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 13786 10152 14044 10180
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 2774 10112 2780 10124
rect 1443 10084 2780 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4652 10115 4710 10121
rect 4652 10112 4664 10115
rect 4212 10084 4664 10112
rect 4212 10072 4218 10084
rect 4652 10081 4664 10084
rect 4698 10081 4710 10115
rect 4652 10075 4710 10081
rect 4755 10115 4813 10121
rect 4755 10081 4767 10115
rect 4801 10112 4813 10115
rect 5810 10112 5816 10124
rect 4801 10084 5816 10112
rect 4801 10081 4813 10084
rect 4755 10075 4813 10081
rect 5810 10072 5816 10084
rect 5868 10112 5874 10124
rect 6914 10112 6920 10124
rect 5868 10084 6920 10112
rect 5868 10072 5874 10084
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7374 10112 7380 10124
rect 7335 10084 7380 10112
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 8665 10115 8723 10121
rect 8665 10081 8677 10115
rect 8711 10112 8723 10115
rect 8754 10112 8760 10124
rect 8711 10084 8760 10112
rect 8711 10081 8723 10084
rect 8665 10075 8723 10081
rect 8754 10072 8760 10084
rect 8812 10072 8818 10124
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9674 10112 9680 10124
rect 9631 10084 9680 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10152 10084 10517 10112
rect 3878 10044 3884 10056
rect 2516 10016 3884 10044
rect 566 9936 572 9988
rect 624 9976 630 9988
rect 2317 9979 2375 9985
rect 2317 9976 2329 9979
rect 624 9948 2329 9976
rect 624 9936 630 9948
rect 2317 9945 2329 9948
rect 2363 9945 2375 9979
rect 2317 9939 2375 9945
rect 661 9911 719 9917
rect 661 9908 673 9911
rect 571 9880 673 9908
rect 661 9877 673 9880
rect 707 9908 719 9911
rect 2516 9908 2544 10016
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 5258 10004 5264 10056
rect 5316 10044 5322 10056
rect 5442 10044 5448 10056
rect 5316 10016 5448 10044
rect 5316 10004 5322 10016
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 8018 10044 8024 10056
rect 5675 10016 8024 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 8018 10004 8024 10016
rect 8076 10044 8082 10056
rect 10152 10044 10180 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10686 10112 10692 10124
rect 10647 10084 10692 10112
rect 10505 10075 10563 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 10870 10072 10876 10124
rect 10928 10112 10934 10124
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 10928 10084 11529 10112
rect 10928 10072 10934 10084
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 11752 10115 11810 10121
rect 11752 10081 11764 10115
rect 11798 10112 11810 10115
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11798 10084 11989 10112
rect 11798 10081 11810 10084
rect 11752 10075 11810 10081
rect 11977 10081 11989 10084
rect 12023 10081 12035 10115
rect 12710 10112 12716 10124
rect 12671 10084 12716 10112
rect 11977 10075 12035 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 13786 10112 13814 10152
rect 13228 10084 13814 10112
rect 13228 10072 13234 10084
rect 8076 10016 10180 10044
rect 8076 10004 8082 10016
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 11839 10047 11897 10053
rect 11839 10044 11851 10047
rect 10468 10016 11851 10044
rect 10468 10004 10474 10016
rect 11839 10013 11851 10016
rect 11885 10044 11897 10047
rect 12250 10044 12256 10056
rect 11885 10016 12256 10044
rect 11885 10013 11897 10016
rect 11839 10007 11897 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 13446 10044 13452 10056
rect 12452 10016 13452 10044
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 4062 9976 4068 9988
rect 2832 9948 4068 9976
rect 2832 9936 2838 9948
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 5074 9976 5080 9988
rect 4667 9948 5080 9976
rect 707 9880 2544 9908
rect 707 9877 719 9880
rect 661 9871 719 9877
rect 385 9775 443 9781
rect 385 9741 397 9775
rect 431 9772 443 9775
rect 566 9772 572 9784
rect 431 9744 572 9772
rect 431 9741 443 9744
rect 385 9735 443 9741
rect 566 9732 572 9744
rect 624 9732 630 9784
rect 566 9634 572 9686
rect 624 9674 630 9686
rect 676 9674 704 9871
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 4667 9908 4695 9948
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 6549 9979 6607 9985
rect 5215 9948 5672 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 5644 9920 5672 9948
rect 6549 9945 6561 9979
rect 6595 9976 6607 9979
rect 9766 9976 9772 9988
rect 6595 9948 9772 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 10321 9979 10379 9985
rect 10321 9945 10333 9979
rect 10367 9976 10379 9979
rect 12452 9976 12480 10016
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 14016 10044 14044 10152
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 14826 10180 14832 10192
rect 14148 10152 14832 10180
rect 14148 10140 14154 10152
rect 14826 10140 14832 10152
rect 14884 10180 14890 10192
rect 17402 10180 17408 10192
rect 14884 10152 17264 10180
rect 17363 10152 17408 10180
rect 14884 10140 14890 10152
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 15930 10112 15936 10124
rect 14792 10084 15936 10112
rect 14792 10072 14798 10084
rect 15930 10072 15936 10084
rect 15988 10112 15994 10124
rect 16152 10115 16210 10121
rect 16152 10112 16164 10115
rect 15988 10084 16164 10112
rect 15988 10072 15994 10084
rect 16152 10081 16164 10084
rect 16198 10081 16210 10115
rect 16152 10075 16210 10081
rect 16255 10115 16313 10121
rect 16255 10081 16267 10115
rect 16301 10112 16313 10115
rect 16850 10112 16856 10124
rect 16301 10084 16856 10112
rect 16301 10081 16313 10084
rect 16255 10075 16313 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17236 10112 17264 10152
rect 17402 10140 17408 10152
rect 17460 10140 17466 10192
rect 17788 10124 17816 10220
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 18104 10220 19717 10248
rect 18104 10208 18110 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 20438 10248 20444 10260
rect 20399 10220 20444 10248
rect 19705 10211 19763 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20993 10251 21051 10257
rect 20993 10248 21005 10251
rect 20588 10220 21005 10248
rect 20588 10208 20594 10220
rect 20993 10217 21005 10220
rect 21039 10217 21051 10251
rect 20993 10211 21051 10217
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 18782 10180 18788 10192
rect 17920 10152 18788 10180
rect 17920 10140 17926 10152
rect 18782 10140 18788 10152
rect 18840 10140 18846 10192
rect 18877 10183 18935 10189
rect 18877 10149 18889 10183
rect 18923 10180 18935 10183
rect 19058 10180 19064 10192
rect 18923 10152 19064 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 17586 10112 17592 10124
rect 17236 10084 17592 10112
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17770 10121 17776 10124
rect 17748 10115 17776 10121
rect 17748 10081 17760 10115
rect 17828 10112 17834 10124
rect 17828 10084 17921 10112
rect 17748 10075 17776 10081
rect 17770 10072 17776 10075
rect 17828 10072 17834 10084
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20806 10112 20812 10124
rect 20036 10084 20812 10112
rect 20036 10072 20042 10084
rect 20806 10072 20812 10084
rect 20864 10112 20870 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20864 10084 20913 10112
rect 20864 10072 20870 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 21453 10115 21511 10121
rect 21453 10081 21465 10115
rect 21499 10112 21511 10115
rect 21726 10112 21732 10124
rect 21499 10084 21732 10112
rect 21499 10081 21511 10084
rect 21453 10075 21511 10081
rect 21726 10072 21732 10084
rect 21784 10072 21790 10124
rect 14829 10047 14887 10053
rect 14829 10044 14841 10047
rect 14016 10016 14841 10044
rect 14829 10013 14841 10016
rect 14875 10013 14887 10047
rect 18782 10044 18788 10056
rect 18743 10016 18788 10044
rect 14829 10007 14887 10013
rect 18782 10004 18788 10016
rect 18840 10044 18846 10056
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 18840 10016 20085 10044
rect 18840 10004 18846 10016
rect 20073 10013 20085 10016
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 10367 9948 12480 9976
rect 10367 9945 10379 9948
rect 10321 9939 10379 9945
rect 12986 9936 12992 9988
rect 13044 9936 13050 9988
rect 13630 9976 13636 9988
rect 13591 9948 13636 9976
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 18690 9976 18696 9988
rect 16908 9948 18696 9976
rect 16908 9936 16914 9948
rect 18690 9936 18696 9948
rect 18748 9936 18754 9988
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 19337 9979 19395 9985
rect 19337 9976 19349 9979
rect 18932 9948 19349 9976
rect 18932 9936 18938 9948
rect 19337 9945 19349 9948
rect 19383 9945 19395 9979
rect 19337 9939 19395 9945
rect 20162 9936 20168 9988
rect 20220 9976 20226 9988
rect 22281 9979 22339 9985
rect 22281 9976 22293 9979
rect 20220 9948 22293 9976
rect 20220 9936 20226 9948
rect 22281 9945 22293 9948
rect 22327 9945 22339 9979
rect 22281 9939 22339 9945
rect 3568 9880 4695 9908
rect 3568 9868 3574 9880
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 6454 9868 6460 9920
rect 6512 9908 6518 9920
rect 6638 9908 6644 9920
rect 6512 9880 6644 9908
rect 6512 9868 6518 9880
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6788 9880 6837 9908
rect 6788 9868 6794 9880
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 6825 9871 6883 9877
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 8018 9908 8024 9920
rect 7064 9880 8024 9908
rect 7064 9868 7070 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8294 9908 8300 9920
rect 8207 9880 8300 9908
rect 8294 9868 8300 9880
rect 8352 9908 8358 9920
rect 8478 9908 8484 9920
rect 8352 9880 8484 9908
rect 8352 9868 8358 9880
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 9088 9880 9413 9908
rect 9088 9868 9094 9880
rect 9401 9877 9413 9880
rect 9447 9908 9459 9911
rect 9858 9908 9864 9920
rect 9447 9880 9864 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10137 9911 10195 9917
rect 10137 9908 10149 9911
rect 10100 9880 10149 9908
rect 10100 9868 10106 9880
rect 10137 9877 10149 9880
rect 10183 9877 10195 9911
rect 10137 9871 10195 9877
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 10827 9911 10885 9917
rect 10827 9908 10839 9911
rect 10744 9880 10839 9908
rect 10744 9868 10750 9880
rect 10827 9877 10839 9880
rect 10873 9877 10885 9911
rect 10827 9871 10885 9877
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13004 9908 13032 9936
rect 12492 9880 13032 9908
rect 12492 9868 12498 9880
rect 15102 9868 15108 9920
rect 15160 9908 15166 9920
rect 15286 9908 15292 9920
rect 15160 9880 15292 9908
rect 15160 9868 15166 9880
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16816 9880 16957 9908
rect 16816 9868 16822 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 17954 9908 17960 9920
rect 17915 9880 17960 9908
rect 16945 9871 17003 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 18230 9908 18236 9920
rect 18191 9880 18236 9908
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18506 9908 18512 9920
rect 18467 9880 18512 9908
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 21910 9908 21916 9920
rect 21871 9880 21916 9908
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 2314 9704 2320 9716
rect 2275 9676 2320 9704
rect 624 9646 704 9674
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 3559 9707 3617 9713
rect 3559 9704 3571 9707
rect 3108 9676 3571 9704
rect 3108 9664 3114 9676
rect 3559 9673 3571 9676
rect 3605 9673 3617 9707
rect 3559 9667 3617 9673
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 4062 9704 4068 9716
rect 3752 9676 4068 9704
rect 3752 9664 3758 9676
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 4614 9704 4620 9716
rect 4488 9676 4620 9704
rect 4488 9664 4494 9676
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 5718 9704 5724 9716
rect 5276 9676 5724 9704
rect 5276 9648 5304 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 7653 9707 7711 9713
rect 6696 9676 7604 9704
rect 6696 9664 6702 9676
rect 624 9634 630 9646
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 2556 9608 2773 9636
rect 2556 9596 2562 9608
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 1762 9528 1768 9580
rect 1820 9568 1826 9580
rect 2038 9568 2044 9580
rect 1820 9540 2044 9568
rect 1820 9528 1826 9540
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2590 9568 2596 9580
rect 2551 9540 2596 9568
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 2745 9568 2773 9608
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 4338 9636 4344 9648
rect 3476 9608 4344 9636
rect 3476 9596 3482 9608
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 4706 9636 4712 9648
rect 4667 9608 4712 9636
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 5258 9596 5264 9648
rect 5316 9596 5322 9648
rect 6089 9639 6147 9645
rect 6089 9605 6101 9639
rect 6135 9636 6147 9639
rect 7098 9636 7104 9648
rect 6135 9608 7104 9636
rect 6135 9605 6147 9608
rect 6089 9599 6147 9605
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7466 9636 7472 9648
rect 7427 9608 7472 9636
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 7576 9636 7604 9676
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 9030 9704 9036 9716
rect 7699 9676 9036 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9674 9704 9680 9716
rect 9635 9676 9680 9704
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 10367 9707 10425 9713
rect 10367 9673 10379 9707
rect 10413 9704 10425 9707
rect 10502 9704 10508 9716
rect 10413 9676 10508 9704
rect 10413 9673 10425 9676
rect 10367 9667 10425 9673
rect 10382 9636 10410 9667
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13081 9707 13139 9713
rect 13081 9704 13093 9707
rect 12768 9676 13093 9704
rect 12768 9664 12774 9676
rect 13081 9673 13093 9676
rect 13127 9673 13139 9707
rect 13081 9667 13139 9673
rect 13722 9664 13728 9716
rect 13780 9704 13786 9716
rect 13906 9704 13912 9716
rect 13780 9676 13912 9704
rect 13780 9664 13786 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 14700 9676 15301 9704
rect 14700 9664 14706 9676
rect 15289 9673 15301 9676
rect 15335 9704 15347 9707
rect 16298 9704 16304 9716
rect 15335 9676 16304 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 17126 9704 17132 9716
rect 17087 9676 17132 9704
rect 17126 9664 17132 9676
rect 17184 9664 17190 9716
rect 17770 9704 17776 9716
rect 17731 9676 17776 9704
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 18138 9664 18144 9716
rect 18196 9704 18202 9716
rect 19751 9707 19809 9713
rect 19751 9704 19763 9707
rect 18196 9676 19763 9704
rect 18196 9664 18202 9676
rect 19751 9673 19763 9676
rect 19797 9673 19809 9707
rect 19751 9667 19809 9673
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20864 9676 20913 9704
rect 20864 9664 20870 9676
rect 20901 9673 20913 9676
rect 20947 9673 20959 9707
rect 20901 9667 20959 9673
rect 21361 9707 21419 9713
rect 21361 9673 21373 9707
rect 21407 9704 21419 9707
rect 22002 9704 22008 9716
rect 21407 9676 22008 9704
rect 21407 9673 21419 9676
rect 21361 9667 21419 9673
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 11379 9639 11437 9645
rect 11379 9636 11391 9639
rect 7576 9608 10410 9636
rect 10933 9608 11391 9636
rect 4430 9568 4436 9580
rect 2745 9540 4436 9568
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5626 9568 5632 9580
rect 4847 9540 5632 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5626 9528 5632 9540
rect 5684 9568 5690 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5684 9540 6193 9568
rect 5684 9528 5690 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 10933 9568 10961 9608
rect 11379 9605 11391 9608
rect 11425 9636 11437 9639
rect 11882 9636 11888 9648
rect 11425 9608 11888 9636
rect 11425 9605 11437 9608
rect 11379 9599 11437 9605
rect 11882 9596 11888 9608
rect 11940 9596 11946 9648
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 14734 9636 14740 9648
rect 12216 9608 14740 9636
rect 12216 9596 12222 9608
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 15381 9639 15439 9645
rect 15381 9605 15393 9639
rect 15427 9636 15439 9639
rect 20530 9636 20536 9648
rect 15427 9608 20536 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 20625 9639 20683 9645
rect 20625 9605 20637 9639
rect 20671 9636 20683 9639
rect 21726 9636 21732 9648
rect 20671 9608 21732 9636
rect 20671 9605 20683 9608
rect 20625 9599 20683 9605
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 11054 9568 11060 9580
rect 8260 9540 10961 9568
rect 11015 9540 11060 9568
rect 8260 9528 8266 9540
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 13495 9571 13553 9577
rect 13495 9537 13507 9571
rect 13541 9568 13553 9571
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 13541 9540 16221 9568
rect 13541 9537 13553 9540
rect 13495 9531 13553 9537
rect 16209 9537 16221 9540
rect 16255 9568 16267 9571
rect 17310 9568 17316 9580
rect 16255 9540 17316 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 17644 9540 18429 9568
rect 17644 9528 17650 9540
rect 18417 9537 18429 9540
rect 18463 9568 18475 9571
rect 18598 9568 18604 9580
rect 18463 9540 18604 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 20036 9540 22109 9568
rect 20036 9528 20042 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 3456 9503 3514 9509
rect 3456 9500 3468 9503
rect 1544 9472 3468 9500
rect 1544 9460 1550 9472
rect 3456 9469 3468 9472
rect 3502 9500 3514 9503
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3502 9472 3893 9500
rect 3502 9469 3514 9472
rect 3456 9463 3514 9469
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4580 9503 4638 9509
rect 4580 9500 4592 9503
rect 4203 9472 4592 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4580 9469 4592 9472
rect 4626 9500 4638 9503
rect 4626 9472 4844 9500
rect 4626 9469 4638 9472
rect 4580 9463 4638 9469
rect 4816 9444 4844 9472
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5132 9472 5457 9500
rect 5132 9460 5138 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6270 9500 6276 9512
rect 6144 9472 6276 9500
rect 6144 9460 6150 9472
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 8570 9500 8576 9512
rect 8076 9472 8576 9500
rect 8076 9460 8082 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9674 9500 9680 9512
rect 9447 9472 9680 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10296 9503 10354 9509
rect 10296 9469 10308 9503
rect 10342 9500 10354 9503
rect 11308 9503 11366 9509
rect 10342 9472 10824 9500
rect 10342 9469 10354 9472
rect 10296 9463 10354 9469
rect 1759 9435 1817 9441
rect 1759 9401 1771 9435
rect 1805 9432 1817 9435
rect 1805 9404 4016 9432
rect 1805 9401 1817 9404
rect 1759 9395 1817 9401
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 2961 9367 3019 9373
rect 2961 9364 2973 9367
rect 2556 9336 2973 9364
rect 2556 9324 2562 9336
rect 2961 9333 2973 9336
rect 3007 9333 3019 9367
rect 3988 9364 4016 9404
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4120 9404 4338 9432
rect 4120 9392 4126 9404
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 3988 9336 4169 9364
rect 2961 9327 3019 9333
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 4310 9364 4338 9404
rect 4430 9392 4436 9444
rect 4488 9432 4494 9444
rect 4488 9404 4533 9432
rect 4488 9392 4494 9404
rect 4798 9392 4804 9444
rect 4856 9392 4862 9444
rect 5169 9435 5227 9441
rect 5169 9401 5181 9435
rect 5215 9432 5227 9435
rect 6914 9432 6920 9444
rect 5215 9404 6684 9432
rect 6875 9404 6920 9432
rect 5215 9401 5227 9404
rect 5169 9395 5227 9401
rect 5184 9364 5212 9395
rect 4310 9336 5212 9364
rect 5905 9367 5963 9373
rect 4157 9327 4215 9333
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 5951 9336 6101 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6089 9333 6101 9336
rect 6135 9333 6147 9367
rect 6089 9327 6147 9333
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6328 9336 6561 9364
rect 6328 9324 6334 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6656 9364 6684 9404
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 7024 9364 7052 9395
rect 7098 9392 7104 9444
rect 7156 9432 7162 9444
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7156 9404 7849 9432
rect 7156 9392 7162 9404
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 8757 9435 8815 9441
rect 8757 9432 8769 9435
rect 8352 9404 8769 9432
rect 8352 9392 8358 9404
rect 8757 9401 8769 9404
rect 8803 9401 8815 9435
rect 8757 9395 8815 9401
rect 8849 9435 8907 9441
rect 8849 9401 8861 9435
rect 8895 9401 8907 9435
rect 10594 9432 10600 9444
rect 8849 9395 8907 9401
rect 9692 9404 10600 9432
rect 7653 9367 7711 9373
rect 7653 9364 7665 9367
rect 6656 9336 7665 9364
rect 6549 9327 6607 9333
rect 7024 9296 7052 9336
rect 7653 9333 7665 9336
rect 7699 9333 7711 9367
rect 7653 9327 7711 9333
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 8076 9336 8401 9364
rect 8076 9324 8082 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 8864 9364 8892 9395
rect 9692 9364 9720 9404
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 10796 9441 10824 9472
rect 11308 9469 11320 9503
rect 11354 9500 11366 9503
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11354 9472 11529 9500
rect 11354 9469 11366 9472
rect 11308 9463 11366 9469
rect 11517 9469 11529 9472
rect 11563 9500 11575 9503
rect 13392 9503 13450 9509
rect 13392 9500 13404 9503
rect 11563 9472 13404 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 13392 9469 13404 9472
rect 13438 9500 13450 9503
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13438 9472 13829 9500
rect 13438 9469 13450 9472
rect 13392 9463 13450 9469
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14458 9500 14464 9512
rect 14415 9472 14464 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 14458 9460 14464 9472
rect 14516 9500 14522 9512
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 14516 9472 15393 9500
rect 14516 9460 14522 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15930 9500 15936 9512
rect 15891 9472 15936 9500
rect 15381 9463 15439 9469
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 16942 9500 16948 9512
rect 16899 9472 16948 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 16942 9460 16948 9472
rect 17000 9500 17006 9512
rect 17862 9500 17868 9512
rect 17000 9472 17868 9500
rect 17000 9460 17006 9472
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 19680 9503 19738 9509
rect 19680 9469 19692 9503
rect 19726 9469 19738 9503
rect 19680 9463 19738 9469
rect 10781 9435 10839 9441
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 15102 9432 15108 9444
rect 10827 9404 15108 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 18138 9432 18144 9444
rect 16356 9404 16401 9432
rect 18099 9404 18144 9432
rect 16356 9392 16362 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18230 9392 18236 9444
rect 18288 9432 18294 9444
rect 18288 9404 18381 9432
rect 18288 9392 18294 9404
rect 18414 9392 18420 9444
rect 18472 9432 18478 9444
rect 18874 9432 18880 9444
rect 18472 9404 18880 9432
rect 18472 9392 18478 9404
rect 18874 9392 18880 9404
rect 18932 9392 18938 9444
rect 19695 9432 19723 9463
rect 19794 9460 19800 9512
rect 19852 9500 19858 9512
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 19852 9472 21189 9500
rect 19852 9460 19858 9472
rect 21177 9469 21189 9472
rect 21223 9500 21235 9503
rect 21223 9472 21864 9500
rect 21223 9469 21235 9472
rect 21177 9463 21235 9469
rect 19695 9404 20208 9432
rect 10042 9364 10048 9376
rect 8619 9336 9720 9364
rect 10003 9336 10048 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 10560 9336 11529 9364
rect 10560 9324 10566 9336
rect 11517 9333 11529 9336
rect 11563 9364 11575 9367
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11563 9336 11713 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 11701 9327 11759 9333
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12158 9364 12164 9376
rect 12023 9336 12164 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12710 9364 12716 9376
rect 12671 9336 12716 9364
rect 12710 9324 12716 9336
rect 12768 9364 12774 9376
rect 14185 9367 14243 9373
rect 14185 9364 14197 9367
rect 12768 9336 14197 9364
rect 12768 9324 12774 9336
rect 14185 9333 14197 9336
rect 14231 9364 14243 9367
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14231 9336 14749 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 15562 9364 15568 9376
rect 15523 9336 15568 9364
rect 14737 9327 14795 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 18248 9364 18276 9392
rect 19058 9364 19064 9376
rect 17920 9336 18276 9364
rect 19019 9336 19064 9364
rect 17920 9324 17926 9336
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20180 9373 20208 9404
rect 20990 9392 20996 9444
rect 21048 9432 21054 9444
rect 21542 9432 21548 9444
rect 21048 9404 21548 9432
rect 21048 9392 21054 9404
rect 21542 9392 21548 9404
rect 21600 9392 21606 9444
rect 21836 9441 21864 9472
rect 21821 9435 21879 9441
rect 21821 9401 21833 9435
rect 21867 9432 21879 9435
rect 22002 9432 22008 9444
rect 21867 9404 22008 9432
rect 21867 9401 21879 9404
rect 21821 9395 21879 9401
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 20165 9367 20223 9373
rect 20165 9333 20177 9367
rect 20211 9364 20223 9367
rect 20254 9364 20260 9376
rect 20211 9336 20260 9364
rect 20211 9333 20223 9336
rect 20165 9327 20223 9333
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 1535 9163 1593 9169
rect 1535 9160 1547 9163
rect 1360 9132 1547 9160
rect 1360 9120 1366 9132
rect 1535 9129 1547 9132
rect 1581 9129 1593 9163
rect 1535 9123 1593 9129
rect 1733 9132 2452 9160
rect 1210 9052 1216 9104
rect 1268 9092 1274 9104
rect 1733 9092 1761 9132
rect 1268 9064 1761 9092
rect 1811 9095 1869 9101
rect 1268 9052 1274 9064
rect 1447 9033 1475 9064
rect 1811 9061 1823 9095
rect 1857 9092 1869 9095
rect 2038 9092 2044 9104
rect 1857 9064 2044 9092
rect 1857 9061 1869 9064
rect 1811 9055 1869 9061
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 2133 9095 2191 9101
rect 2133 9061 2145 9095
rect 2179 9092 2191 9095
rect 2314 9092 2320 9104
rect 2179 9064 2320 9092
rect 2179 9061 2191 9064
rect 2133 9055 2191 9061
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 2424 9092 2452 9132
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 3292 9132 4154 9160
rect 3292 9120 3298 9132
rect 3697 9095 3755 9101
rect 3697 9092 3709 9095
rect 2424 9064 3709 9092
rect 3697 9061 3709 9064
rect 3743 9061 3755 9095
rect 4126 9092 4154 9132
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 5442 9160 5448 9172
rect 4488 9132 5448 9160
rect 4488 9120 4494 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5626 9160 5632 9172
rect 5539 9132 5632 9160
rect 5626 9120 5632 9132
rect 5684 9160 5690 9172
rect 7024 9160 7052 9200
rect 7929 9163 7987 9169
rect 5684 9132 7788 9160
rect 5684 9120 5690 9132
rect 4890 9092 4896 9104
rect 4126 9064 4896 9092
rect 3697 9055 3755 9061
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 6178 9092 6184 9104
rect 5040 9064 5085 9092
rect 5137 9064 6184 9092
rect 5040 9052 5046 9064
rect 1432 9027 1490 9033
rect 1432 8993 1444 9027
rect 1478 8993 1490 9027
rect 1432 8987 1490 8993
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 1708 9027 1766 9033
rect 1708 9024 1720 9027
rect 1636 8996 1720 9024
rect 1636 8984 1642 8996
rect 1708 8993 1720 8996
rect 1754 8993 1766 9027
rect 1708 8987 1766 8993
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 4709 9027 4767 9033
rect 2740 8996 2785 9024
rect 2740 8984 2746 8996
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 5137 9024 5165 9064
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 6656 9101 6684 9132
rect 6641 9095 6699 9101
rect 6641 9061 6653 9095
rect 6687 9061 6699 9095
rect 6822 9092 6828 9104
rect 6641 9055 6699 9061
rect 6748 9064 6828 9092
rect 4755 8996 5165 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 5994 9024 6000 9036
rect 5500 8996 6000 9024
rect 5500 8984 5506 8996
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 106 8956 112 8968
rect 67 8928 112 8956
rect 106 8916 112 8928
rect 164 8916 170 8968
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 937 8891 995 8897
rect 937 8857 949 8891
rect 983 8888 995 8891
rect 1026 8888 1032 8900
rect 983 8860 1032 8888
rect 983 8857 995 8860
rect 937 8851 995 8857
rect 1026 8848 1032 8860
rect 1084 8848 1090 8900
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 2056 8888 2084 8919
rect 2314 8916 2320 8968
rect 2372 8956 2378 8968
rect 3142 8956 3148 8968
rect 2372 8928 3148 8956
rect 2372 8916 2378 8928
rect 3142 8916 3148 8928
rect 3200 8956 3206 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3200 8928 3341 8956
rect 3200 8916 3206 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 4982 8956 4988 8968
rect 3329 8919 3387 8925
rect 4724 8928 4988 8956
rect 1820 8860 2084 8888
rect 1820 8848 1826 8860
rect 4724 8832 4752 8928
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6638 8956 6644 8968
rect 6595 8928 6644 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 6270 8888 6276 8900
rect 4856 8860 6276 8888
rect 4856 8848 4862 8860
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 2958 8820 2964 8832
rect 1452 8792 2964 8820
rect 1452 8780 1458 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3234 8820 3240 8832
rect 3099 8792 3240 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4706 8820 4712 8832
rect 4203 8792 4712 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4706 8780 4712 8792
rect 4764 8820 4770 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 4764 8792 5917 8820
rect 4764 8780 4770 8792
rect 5905 8789 5917 8792
rect 5951 8820 5963 8823
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5951 8792 6101 8820
rect 5951 8789 5963 8792
rect 5905 8783 5963 8789
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 6089 8783 6147 8789
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 6748 8820 6776 9064
rect 6822 9052 6828 9064
rect 6880 9092 6886 9104
rect 7024 9092 7052 9132
rect 6880 9064 7052 9092
rect 7193 9095 7251 9101
rect 6880 9052 6886 9064
rect 7193 9061 7205 9095
rect 7239 9092 7251 9095
rect 7558 9092 7564 9104
rect 7239 9064 7564 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 7760 9092 7788 9132
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8018 9160 8024 9172
rect 7975 9132 8024 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8205 9163 8263 9169
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8662 9160 8668 9172
rect 8251 9132 8668 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 10192 9132 10241 9160
rect 10192 9120 10198 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 10318 9120 10324 9172
rect 10376 9160 10382 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10376 9132 10425 9160
rect 10376 9120 10382 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10870 9160 10876 9172
rect 10413 9123 10471 9129
rect 10520 9132 10876 9160
rect 10520 9092 10548 9132
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11241 9163 11299 9169
rect 11241 9129 11253 9163
rect 11287 9160 11299 9163
rect 12710 9160 12716 9172
rect 11287 9132 12716 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 13354 9160 13360 9172
rect 12912 9132 13360 9160
rect 11698 9092 11704 9104
rect 7760 9064 10548 9092
rect 11624 9064 11704 9092
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 8168 8996 8585 9024
rect 8168 8984 8174 8996
rect 8573 8993 8585 8996
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 8812 8996 9689 9024
rect 8812 8984 8818 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 6880 8928 8953 8956
rect 6880 8916 6886 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 8987 8928 9321 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9692 8956 9720 8987
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10284 8996 10885 9024
rect 10284 8984 10290 8996
rect 10873 8993 10885 8996
rect 10919 9024 10931 9027
rect 11624 9024 11652 9064
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 12912 9101 12940 9132
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14458 9160 14464 9172
rect 13780 9120 13814 9160
rect 14419 9132 14464 9160
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 15427 9163 15485 9169
rect 15427 9160 15439 9163
rect 14608 9132 15439 9160
rect 14608 9120 14614 9132
rect 15427 9129 15439 9132
rect 15473 9129 15485 9163
rect 15427 9123 15485 9129
rect 16209 9163 16267 9169
rect 16209 9129 16221 9163
rect 16255 9160 16267 9163
rect 16298 9160 16304 9172
rect 16255 9132 16304 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 19058 9160 19064 9172
rect 17828 9132 19064 9160
rect 17828 9120 17834 9132
rect 12897 9095 12955 9101
rect 12897 9061 12909 9095
rect 12943 9061 12955 9095
rect 13786 9092 13814 9120
rect 14826 9092 14832 9104
rect 13786 9064 14832 9092
rect 12897 9055 12955 9061
rect 14826 9052 14832 9064
rect 14884 9052 14890 9104
rect 16574 9052 16580 9104
rect 16632 9092 16638 9104
rect 16714 9095 16772 9101
rect 16714 9092 16726 9095
rect 16632 9064 16726 9092
rect 16632 9052 16638 9064
rect 16714 9061 16726 9064
rect 16760 9061 16772 9095
rect 18046 9092 18052 9104
rect 18007 9064 18052 9092
rect 16714 9055 16772 9061
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 18340 9101 18368 9132
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 19242 9120 19248 9172
rect 19300 9160 19306 9172
rect 19843 9163 19901 9169
rect 19843 9160 19855 9163
rect 19300 9132 19855 9160
rect 19300 9120 19306 9132
rect 19843 9129 19855 9132
rect 19889 9160 19901 9163
rect 21910 9160 21916 9172
rect 19889 9132 21916 9160
rect 19889 9129 19901 9132
rect 19843 9123 19901 9129
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 18325 9095 18383 9101
rect 18325 9061 18337 9095
rect 18371 9061 18383 9095
rect 18325 9055 18383 9061
rect 18598 9052 18604 9104
rect 18656 9092 18662 9104
rect 19334 9092 19340 9104
rect 18656 9064 19340 9092
rect 18656 9052 18662 9064
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 20533 9095 20591 9101
rect 20533 9092 20545 9095
rect 19668 9064 20545 9092
rect 19668 9052 19674 9064
rect 20533 9061 20545 9064
rect 20579 9061 20591 9095
rect 20990 9092 20996 9104
rect 20951 9064 20996 9092
rect 20533 9055 20591 9061
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 21082 9052 21088 9104
rect 21140 9092 21146 9104
rect 21140 9064 21185 9092
rect 21140 9052 21146 9064
rect 10919 8996 11652 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 13906 9024 13912 9036
rect 13688 8996 13912 9024
rect 13688 8984 13694 8996
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 15356 9027 15414 9033
rect 15356 8993 15368 9027
rect 15402 8993 15414 9027
rect 15356 8987 15414 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 16850 9024 16856 9036
rect 16439 8996 16856 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 9766 8956 9772 8968
rect 9692 8928 9772 8956
rect 9309 8919 9367 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 12032 8928 12173 8956
rect 12032 8916 12038 8928
rect 12161 8925 12173 8928
rect 12207 8956 12219 8959
rect 12250 8956 12256 8968
rect 12207 8928 12256 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12802 8956 12808 8968
rect 12763 8928 12808 8956
rect 12802 8916 12808 8928
rect 12860 8956 12866 8968
rect 13262 8956 13268 8968
rect 12860 8928 13268 8956
rect 12860 8916 12866 8928
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 14642 8956 14648 8968
rect 14332 8928 14648 8956
rect 14332 8916 14338 8928
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15371 8956 15399 8987
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 9024 18935 9027
rect 19058 9024 19064 9036
rect 18923 8996 19064 9024
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 19058 8984 19064 8996
rect 19116 9024 19122 9036
rect 19518 9024 19524 9036
rect 19116 8996 19524 9024
rect 19116 8984 19122 8996
rect 19518 8984 19524 8996
rect 19576 8984 19582 9036
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 19794 9024 19800 9036
rect 19751 8996 19800 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 15160 8928 17816 8956
rect 15160 8916 15166 8928
rect 7466 8888 7472 8900
rect 7427 8860 7472 8888
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 7742 8848 7748 8900
rect 7800 8888 7806 8900
rect 12437 8891 12495 8897
rect 12437 8888 12449 8891
rect 7800 8860 12449 8888
rect 7800 8848 7806 8860
rect 12437 8857 12449 8860
rect 12483 8857 12495 8891
rect 12437 8851 12495 8857
rect 13357 8891 13415 8897
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 13630 8888 13636 8900
rect 13403 8860 13636 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 17589 8891 17647 8897
rect 17589 8888 17601 8891
rect 14516 8860 17601 8888
rect 14516 8848 14522 8860
rect 17589 8857 17601 8860
rect 17635 8857 17647 8891
rect 17788 8888 17816 8928
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18012 8928 18245 8956
rect 18012 8916 18018 8928
rect 18233 8925 18245 8928
rect 18279 8956 18291 8959
rect 18279 8928 19472 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18690 8888 18696 8900
rect 17788 8860 18696 8888
rect 17589 8851 17647 8857
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 19444 8888 19472 8928
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 19668 8928 20177 8956
rect 19668 8916 19674 8928
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 22281 8959 22339 8965
rect 22281 8956 22293 8959
rect 20165 8919 20223 8925
rect 21100 8928 22293 8956
rect 21100 8888 21128 8928
rect 22281 8925 22293 8928
rect 22327 8925 22339 8959
rect 22281 8919 22339 8925
rect 19444 8860 21128 8888
rect 21545 8891 21603 8897
rect 21545 8857 21557 8891
rect 21591 8888 21603 8891
rect 21634 8888 21640 8900
rect 21591 8860 21640 8888
rect 21591 8857 21603 8860
rect 21545 8851 21603 8857
rect 21634 8848 21640 8860
rect 21692 8848 21698 8900
rect 6696 8792 6776 8820
rect 8757 8823 8815 8829
rect 6696 8780 6702 8792
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9122 8820 9128 8832
rect 8803 8792 9128 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9858 8820 9864 8832
rect 9819 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10413 8823 10471 8829
rect 10413 8820 10425 8823
rect 10284 8792 10425 8820
rect 10284 8780 10290 8792
rect 10413 8789 10425 8792
rect 10459 8820 10471 8823
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10459 8792 10609 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 11793 8823 11851 8829
rect 11793 8789 11805 8823
rect 11839 8820 11851 8823
rect 12158 8820 12164 8832
rect 11839 8792 12164 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 13722 8820 13728 8832
rect 13683 8792 13728 8820
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14829 8823 14887 8829
rect 14829 8789 14841 8823
rect 14875 8820 14887 8823
rect 15010 8820 15016 8832
rect 14875 8792 15016 8820
rect 14875 8789 14887 8792
rect 14829 8783 14887 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 17310 8820 17316 8832
rect 17271 8792 17316 8820
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 18322 8780 18328 8832
rect 18380 8820 18386 8832
rect 19153 8823 19211 8829
rect 19153 8820 19165 8823
rect 18380 8792 19165 8820
rect 18380 8780 18386 8792
rect 19153 8789 19165 8792
rect 19199 8789 19211 8823
rect 19610 8820 19616 8832
rect 19571 8792 19616 8820
rect 19153 8783 19211 8789
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 20530 8820 20536 8832
rect 19944 8792 20536 8820
rect 19944 8780 19950 8792
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 21910 8820 21916 8832
rect 21871 8792 21916 8820
rect 21910 8780 21916 8792
rect 21968 8780 21974 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1535 8619 1593 8625
rect 1535 8616 1547 8619
rect 1452 8588 1547 8616
rect 1452 8576 1458 8588
rect 1535 8585 1547 8588
rect 1581 8585 1593 8619
rect 1535 8579 1593 8585
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 3234 8616 3240 8628
rect 2004 8588 3240 8616
rect 2004 8576 2010 8588
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3510 8616 3516 8628
rect 3467 8588 3516 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3844 8588 3985 8616
rect 3844 8576 3850 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 6089 8619 6147 8625
rect 3973 8579 4031 8585
rect 4126 8588 5948 8616
rect 106 8508 112 8560
rect 164 8548 170 8560
rect 4126 8548 4154 8588
rect 164 8520 4154 8548
rect 164 8508 170 8520
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 4985 8551 5043 8557
rect 4985 8548 4997 8551
rect 4764 8520 4997 8548
rect 4764 8508 4770 8520
rect 4985 8517 4997 8520
rect 5031 8548 5043 8551
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 5031 8520 5089 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 5920 8548 5948 8588
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6135 8588 6193 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6181 8585 6193 8588
rect 6227 8616 6239 8619
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6227 8588 6561 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 8076 8588 8125 8616
rect 8076 8576 8082 8588
rect 8113 8585 8125 8588
rect 8159 8616 8171 8619
rect 10686 8616 10692 8628
rect 8159 8588 10692 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11514 8616 11520 8628
rect 10928 8588 11520 8616
rect 10928 8576 10934 8588
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13412 8588 13461 8616
rect 13412 8576 13418 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 13630 8576 13636 8628
rect 13688 8576 13694 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 15102 8616 15108 8628
rect 13872 8588 13917 8616
rect 15063 8588 15108 8616
rect 13872 8576 13878 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15470 8616 15476 8628
rect 15212 8588 15476 8616
rect 9858 8548 9864 8560
rect 5920 8520 9864 8548
rect 5077 8511 5135 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 11054 8548 11060 8560
rect 10967 8520 11060 8548
rect 11054 8508 11060 8520
rect 11112 8548 11118 8560
rect 11790 8548 11796 8560
rect 11112 8520 11796 8548
rect 11112 8508 11118 8520
rect 11790 8508 11796 8520
rect 11848 8548 11854 8560
rect 13372 8548 13400 8576
rect 11848 8520 13400 8548
rect 13648 8548 13676 8576
rect 13648 8520 13814 8548
rect 11848 8508 11854 8520
rect 569 8483 627 8489
rect 569 8449 581 8483
rect 615 8480 627 8483
rect 3142 8480 3148 8492
rect 615 8452 3148 8480
rect 615 8449 627 8452
rect 569 8443 627 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 4246 8480 4252 8492
rect 3319 8452 4252 8480
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 1708 8415 1766 8421
rect 1708 8412 1720 8415
rect 1550 8384 1720 8412
rect 14 8304 20 8356
rect 72 8344 78 8356
rect 1550 8344 1578 8384
rect 1708 8381 1720 8384
rect 1754 8381 1766 8415
rect 1708 8375 1766 8381
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3319 8412 3347 8452
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 5905 8483 5963 8489
rect 4488 8452 5120 8480
rect 4488 8440 4494 8452
rect 5092 8424 5120 8452
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7374 8480 7380 8492
rect 5951 8452 7380 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7374 8440 7380 8452
rect 7432 8480 7438 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 7432 8452 8677 8480
rect 7432 8440 7438 8452
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 8904 8452 9321 8480
rect 8904 8440 8910 8452
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 9309 8443 9367 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10134 8480 10140 8492
rect 10095 8452 10140 8480
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10502 8480 10508 8492
rect 10382 8452 10508 8480
rect 3016 8384 3347 8412
rect 3016 8372 3022 8384
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3568 8384 3709 8412
rect 3568 8372 3574 8384
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8412 3939 8415
rect 4338 8412 4344 8424
rect 3927 8384 4344 8412
rect 3927 8381 3939 8384
rect 3881 8375 3939 8381
rect 2225 8347 2283 8353
rect 2225 8344 2237 8347
rect 72 8316 1578 8344
rect 1733 8316 2237 8344
rect 72 8304 78 8316
rect 934 8236 940 8288
rect 992 8276 998 8288
rect 1733 8276 1761 8316
rect 2225 8313 2237 8316
rect 2271 8313 2283 8347
rect 2225 8307 2283 8313
rect 2317 8347 2375 8353
rect 2317 8313 2329 8347
rect 2363 8344 2375 8347
rect 2406 8344 2412 8356
rect 2363 8316 2412 8344
rect 2363 8313 2375 8316
rect 2317 8307 2375 8313
rect 2406 8304 2412 8316
rect 2464 8304 2470 8356
rect 2866 8344 2872 8356
rect 2827 8316 2872 8344
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 3234 8344 3240 8356
rect 3195 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3712 8344 3740 8375
rect 4338 8372 4344 8384
rect 4396 8412 4402 8424
rect 4396 8384 4660 8412
rect 4396 8372 4402 8384
rect 4154 8344 4160 8356
rect 3712 8316 4160 8344
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 4632 8344 4660 8384
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 6871 8384 7481 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7469 8381 7481 8384
rect 7515 8412 7527 8415
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7515 8384 7941 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 7929 8375 7987 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 5261 8347 5319 8353
rect 4304 8316 4936 8344
rect 4304 8304 4310 8316
rect 992 8248 1761 8276
rect 1811 8279 1869 8285
rect 992 8236 998 8248
rect 1811 8245 1823 8279
rect 1857 8276 1869 8279
rect 2958 8276 2964 8288
rect 1857 8248 2964 8276
rect 1857 8245 1869 8248
rect 1811 8239 1869 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 3605 8279 3663 8285
rect 3605 8276 3617 8279
rect 3467 8248 3617 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 3605 8245 3617 8248
rect 3651 8276 3663 8279
rect 3786 8276 3792 8288
rect 3651 8248 3792 8276
rect 3651 8245 3663 8248
rect 3605 8239 3663 8245
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4632 8285 4660 8316
rect 4617 8279 4675 8285
rect 4617 8245 4629 8279
rect 4663 8276 4675 8279
rect 4706 8276 4712 8288
rect 4663 8248 4712 8276
rect 4663 8245 4675 8248
rect 4617 8239 4675 8245
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 4908 8276 4936 8316
rect 5261 8313 5273 8347
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5626 8344 5632 8356
rect 5399 8316 5632 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5166 8276 5172 8288
rect 4908 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5276 8276 5304 8307
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 8202 8344 8208 8356
rect 6104 8316 8208 8344
rect 6104 8276 6132 8316
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8386 8344 8392 8356
rect 8347 8316 8392 8344
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 9858 8344 9864 8356
rect 8536 8316 8581 8344
rect 8909 8316 9864 8344
rect 8536 8304 8542 8316
rect 7006 8276 7012 8288
rect 5276 8248 6132 8276
rect 6967 8248 7012 8276
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7374 8276 7380 8288
rect 7156 8248 7380 8276
rect 7156 8236 7162 8248
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7929 8279 7987 8285
rect 7929 8245 7941 8279
rect 7975 8276 7987 8279
rect 8909 8276 8937 8316
rect 9858 8304 9864 8316
rect 9916 8344 9922 8356
rect 10382 8344 10410 8452
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11422 8440 11428 8492
rect 11480 8480 11486 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 11480 8452 12541 8480
rect 11480 8440 11486 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 13630 8480 13636 8492
rect 12768 8452 13636 8480
rect 12768 8440 12774 8452
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 12250 8412 12256 8424
rect 11572 8384 12256 8412
rect 11572 8372 11578 8384
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 10502 8353 10508 8356
rect 9916 8316 10410 8344
rect 9916 8304 9922 8316
rect 10499 8307 10508 8353
rect 10560 8344 10566 8356
rect 12621 8347 12679 8353
rect 10560 8316 11468 8344
rect 10502 8304 10508 8307
rect 10560 8304 10566 8316
rect 11440 8288 11468 8316
rect 12621 8313 12633 8347
rect 12667 8313 12679 8347
rect 13170 8344 13176 8356
rect 13131 8316 13176 8344
rect 12621 8307 12679 8313
rect 11422 8276 11428 8288
rect 7975 8248 8937 8276
rect 11383 8248 11428 8276
rect 7975 8245 7987 8248
rect 7929 8239 7987 8245
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 12158 8276 12164 8288
rect 12119 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8276 12222 8288
rect 12636 8276 12664 8307
rect 13170 8304 13176 8316
rect 13228 8344 13234 8356
rect 13786 8344 13814 8520
rect 14550 8508 14556 8560
rect 14608 8548 14614 8560
rect 15212 8548 15240 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16040 8588 16405 8616
rect 16040 8548 16068 8588
rect 16393 8585 16405 8588
rect 16439 8616 16451 8619
rect 16574 8616 16580 8628
rect 16439 8588 16580 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 16850 8616 16856 8628
rect 16811 8588 16856 8616
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 17083 8619 17141 8625
rect 17083 8585 17095 8619
rect 17129 8616 17141 8619
rect 18782 8616 18788 8628
rect 17129 8588 18788 8616
rect 17129 8585 17141 8588
rect 17083 8579 17141 8585
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 18932 8588 19533 8616
rect 18932 8576 18938 8588
rect 19521 8585 19533 8588
rect 19567 8616 19579 8619
rect 19794 8616 19800 8628
rect 19567 8588 19800 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20864 8588 20913 8616
rect 20864 8576 20870 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 21315 8619 21373 8625
rect 21315 8585 21327 8619
rect 21361 8616 21373 8619
rect 21910 8616 21916 8628
rect 21361 8588 21916 8616
rect 21361 8585 21373 8588
rect 21315 8579 21373 8585
rect 14608 8520 15240 8548
rect 15396 8520 16068 8548
rect 16117 8551 16175 8557
rect 14608 8508 14614 8520
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14332 8452 14749 8480
rect 14332 8440 14338 8452
rect 14737 8449 14749 8452
rect 14783 8480 14795 8483
rect 15396 8480 15424 8520
rect 16117 8517 16129 8551
rect 16163 8548 16175 8551
rect 19886 8548 19892 8560
rect 16163 8520 19892 8548
rect 16163 8517 16175 8520
rect 16117 8511 16175 8517
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 20990 8508 20996 8560
rect 21048 8548 21054 8560
rect 21330 8548 21358 8579
rect 21910 8576 21916 8588
rect 21968 8576 21974 8628
rect 21048 8520 21358 8548
rect 21048 8508 21054 8520
rect 21542 8508 21548 8560
rect 21600 8548 21606 8560
rect 22005 8551 22063 8557
rect 22005 8548 22017 8551
rect 21600 8520 22017 8548
rect 21600 8508 21606 8520
rect 22005 8517 22017 8520
rect 22051 8517 22063 8551
rect 22005 8511 22063 8517
rect 14783 8452 15424 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 14976 8384 15209 8412
rect 14976 8372 14982 8384
rect 15197 8381 15209 8384
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 15396 8344 15424 8452
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 17862 8480 17868 8492
rect 15528 8452 17868 8480
rect 15528 8440 15534 8452
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8480 18199 8483
rect 19242 8480 19248 8492
rect 18187 8452 19248 8480
rect 18187 8449 18199 8452
rect 18141 8443 18199 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 20438 8480 20444 8492
rect 19751 8452 20444 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 15930 8372 15936 8424
rect 15988 8412 15994 8424
rect 17012 8415 17070 8421
rect 17012 8412 17024 8415
rect 15988 8384 17024 8412
rect 15988 8372 15994 8384
rect 17012 8381 17024 8384
rect 17058 8412 17070 8415
rect 17218 8412 17224 8424
rect 17058 8384 17224 8412
rect 17058 8381 17070 8384
rect 17012 8375 17070 8381
rect 17218 8372 17224 8384
rect 17276 8412 17282 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 17276 8384 17417 8412
rect 17276 8372 17282 8384
rect 17405 8381 17417 8384
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8412 18843 8415
rect 19058 8412 19064 8424
rect 18831 8384 19064 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 21244 8415 21302 8421
rect 21244 8381 21256 8415
rect 21290 8412 21302 8415
rect 21726 8412 21732 8424
rect 21290 8384 21732 8412
rect 21290 8381 21302 8384
rect 21244 8375 21302 8381
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 15518 8347 15576 8353
rect 15518 8344 15530 8347
rect 13228 8316 14274 8344
rect 15396 8316 15530 8344
rect 13228 8304 13234 8316
rect 12216 8248 12664 8276
rect 12216 8236 12222 8248
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 12768 8248 14013 8276
rect 12768 8236 12774 8248
rect 14001 8245 14013 8248
rect 14047 8245 14059 8279
rect 14246 8276 14274 8316
rect 15518 8313 15530 8316
rect 15564 8313 15576 8347
rect 15518 8307 15576 8313
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 18233 8347 18291 8353
rect 18233 8344 18245 8347
rect 17368 8316 18245 8344
rect 17368 8304 17374 8316
rect 18233 8313 18245 8316
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 16022 8276 16028 8288
rect 14246 8248 16028 8276
rect 14001 8239 14059 8245
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 17770 8276 17776 8288
rect 17731 8248 17776 8276
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 18248 8276 18276 8307
rect 18414 8304 18420 8356
rect 18472 8344 18478 8356
rect 18472 8316 19702 8344
rect 18472 8304 18478 8316
rect 19061 8279 19119 8285
rect 19061 8276 19073 8279
rect 18248 8248 19073 8276
rect 19061 8245 19073 8248
rect 19107 8276 19119 8279
rect 19334 8276 19340 8288
rect 19107 8248 19340 8276
rect 19107 8245 19119 8248
rect 19061 8239 19119 8245
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 19674 8276 19702 8316
rect 19794 8304 19800 8356
rect 19852 8344 19858 8356
rect 20349 8347 20407 8353
rect 19852 8316 19897 8344
rect 19852 8304 19858 8316
rect 20349 8313 20361 8347
rect 20395 8313 20407 8347
rect 22094 8344 22100 8356
rect 20349 8307 20407 8313
rect 21284 8316 22100 8344
rect 20364 8276 20392 8307
rect 21284 8288 21312 8316
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 21266 8276 21272 8288
rect 19674 8248 21272 8276
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 22462 8276 22468 8288
rect 22423 8248 22468 8276
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 6914 8072 6920 8084
rect 1479 8044 6920 8072
rect 1479 7945 1507 8044
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 8159 8075 8217 8081
rect 8159 8072 8171 8075
rect 7340 8044 8171 8072
rect 7340 8032 7346 8044
rect 8159 8041 8171 8044
rect 8205 8041 8217 8075
rect 8159 8035 8217 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8352 8044 8953 8072
rect 8352 8032 8358 8044
rect 8941 8041 8953 8044
rect 8987 8072 8999 8075
rect 9398 8072 9404 8084
rect 8987 8044 9404 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10502 8072 10508 8084
rect 10275 8044 10508 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 11146 8072 11152 8084
rect 10933 8044 11152 8072
rect 2130 8004 2136 8016
rect 1964 7976 2136 8004
rect 1464 7939 1522 7945
rect 1464 7905 1476 7939
rect 1510 7905 1522 7939
rect 1464 7899 1522 7905
rect 1724 7939 1782 7945
rect 1724 7905 1736 7939
rect 1770 7936 1782 7939
rect 1964 7936 1992 7976
rect 2130 7964 2136 7976
rect 2188 7964 2194 8016
rect 2225 8007 2283 8013
rect 2225 7973 2237 8007
rect 2271 8004 2283 8007
rect 2406 8004 2412 8016
rect 2271 7976 2412 8004
rect 2271 7973 2283 7976
rect 2225 7967 2283 7973
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 3050 8004 3056 8016
rect 3011 7976 3056 8004
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 4890 7964 4896 8016
rect 4948 8004 4954 8016
rect 5071 8007 5129 8013
rect 5071 8004 5083 8007
rect 4948 7976 5083 8004
rect 4948 7964 4954 7976
rect 5071 7973 5083 7976
rect 5117 8004 5129 8007
rect 5905 8007 5963 8013
rect 5905 8004 5917 8007
rect 5117 7976 5917 8004
rect 5117 7973 5129 7976
rect 5071 7967 5129 7973
rect 5905 7973 5917 7976
rect 5951 8004 5963 8007
rect 6273 8007 6331 8013
rect 6273 8004 6285 8007
rect 5951 7976 6285 8004
rect 5951 7973 5963 7976
rect 5905 7967 5963 7973
rect 6273 7973 6285 7976
rect 6319 7973 6331 8007
rect 6546 8004 6552 8016
rect 6507 7976 6552 8004
rect 6273 7967 6331 7973
rect 1770 7908 1992 7936
rect 1770 7905 1782 7908
rect 1724 7899 1782 7905
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4709 7939 4767 7945
rect 4212 7908 4521 7936
rect 4212 7896 4218 7908
rect 1811 7871 1869 7877
rect 1811 7837 1823 7871
rect 1857 7868 1869 7871
rect 1946 7868 1952 7880
rect 1857 7840 1952 7868
rect 1857 7837 1869 7840
rect 1811 7831 1869 7837
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 2056 7840 2145 7868
rect 658 7760 664 7812
rect 716 7800 722 7812
rect 1394 7800 1400 7812
rect 716 7772 1400 7800
rect 716 7760 722 7772
rect 1394 7760 1400 7772
rect 1452 7800 1458 7812
rect 2056 7800 2084 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3142 7868 3148 7880
rect 3007 7840 3148 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 4493 7868 4521 7908
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 5350 7936 5356 7948
rect 4755 7908 5356 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 6288 7936 6316 7967
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 6641 8007 6699 8013
rect 6641 7973 6653 8007
rect 6687 8004 6699 8007
rect 7742 8004 7748 8016
rect 6687 7976 7748 8004
rect 6687 7973 6699 7976
rect 6641 7967 6699 7973
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8481 8007 8539 8013
rect 8481 8004 8493 8007
rect 7892 7976 8493 8004
rect 7892 7964 7898 7976
rect 8481 7973 8493 7976
rect 8527 7973 8539 8007
rect 10933 8004 10961 8044
rect 11146 8032 11152 8044
rect 11204 8072 11210 8084
rect 12437 8075 12495 8081
rect 11204 8044 11652 8072
rect 11204 8032 11210 8044
rect 11054 8004 11060 8016
rect 8481 7967 8539 7973
rect 8772 7976 10961 8004
rect 11015 7976 11060 8004
rect 6288 7908 6454 7936
rect 6270 7868 6276 7880
rect 3651 7840 6276 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 2682 7800 2688 7812
rect 1452 7772 2084 7800
rect 2643 7772 2688 7800
rect 1452 7760 1458 7772
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 4493 7800 4521 7840
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 5994 7800 6000 7812
rect 3292 7772 6000 7800
rect 3292 7760 3298 7772
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 1627 7735 1685 7741
rect 1627 7732 1639 7735
rect 1544 7704 1639 7732
rect 1544 7692 1550 7704
rect 1627 7701 1639 7704
rect 1673 7701 1685 7735
rect 1627 7695 1685 7701
rect 2958 7692 2964 7744
rect 3016 7732 3022 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 3016 7704 4261 7732
rect 3016 7692 3022 7704
rect 4249 7701 4261 7704
rect 4295 7732 4307 7735
rect 4430 7732 4436 7744
rect 4295 7704 4436 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4534 7732 4562 7772
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 5626 7732 5632 7744
rect 4534 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7732 5690 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5684 7704 6193 7732
rect 5684 7692 5690 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 6426 7732 6454 7908
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 8110 7945 8116 7948
rect 8056 7939 8116 7945
rect 8056 7936 8068 7939
rect 7616 7908 8068 7936
rect 7616 7896 7622 7908
rect 8056 7905 8068 7908
rect 8102 7905 8116 7939
rect 8056 7899 8116 7905
rect 8110 7896 8116 7899
rect 8168 7896 8174 7948
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8772 7936 8800 7976
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11624 8013 11652 8044
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12526 8072 12532 8084
rect 12483 8044 12532 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13446 8072 13452 8084
rect 13035 8044 13452 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 11609 8007 11667 8013
rect 11609 7973 11621 8007
rect 11655 7973 11667 8007
rect 11609 7967 11667 7973
rect 12342 7964 12348 8016
rect 12400 8004 12406 8016
rect 13004 8004 13032 8035
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 13998 8032 14004 8084
rect 14056 8072 14062 8084
rect 14734 8072 14740 8084
rect 14056 8044 14740 8072
rect 14056 8032 14062 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16945 8075 17003 8081
rect 15712 8044 16062 8072
rect 15712 8032 15718 8044
rect 13078 8004 13084 8016
rect 12400 7976 13032 8004
rect 13039 7976 13084 8004
rect 12400 7964 12406 7976
rect 13078 7964 13084 7976
rect 13136 7964 13142 8016
rect 13354 7964 13360 8016
rect 13412 8004 13418 8016
rect 13541 8007 13599 8013
rect 13541 8004 13553 8007
rect 13412 7976 13553 8004
rect 13412 7964 13418 7976
rect 13541 7973 13553 7976
rect 13587 7973 13599 8007
rect 13541 7967 13599 7973
rect 13630 7964 13636 8016
rect 13688 8004 13694 8016
rect 13688 7976 13733 8004
rect 13688 7964 13694 7976
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 14642 8004 14648 8016
rect 14516 7976 14648 8004
rect 14516 7964 14522 7976
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15930 8004 15936 8016
rect 15672 7976 15936 8004
rect 15672 7948 15700 7976
rect 15930 7964 15936 7976
rect 15988 7964 15994 8016
rect 16034 8004 16062 8044
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17770 8072 17776 8084
rect 16991 8044 17776 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 20806 8072 20812 8084
rect 19392 8044 20812 8072
rect 19392 8032 19398 8044
rect 20806 8032 20812 8044
rect 20864 8072 20870 8084
rect 20864 8044 21128 8072
rect 20864 8032 20870 8044
rect 16390 8013 16396 8016
rect 16034 7976 16344 8004
rect 8444 7908 8800 7936
rect 8444 7896 8450 7908
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9490 7936 9496 7948
rect 8904 7908 9496 7936
rect 8904 7896 8910 7908
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 13170 7936 13176 7948
rect 11756 7908 13176 7936
rect 11756 7896 11762 7908
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 15654 7896 15660 7948
rect 15712 7896 15718 7948
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 16025 7939 16083 7945
rect 16025 7936 16037 7939
rect 15896 7908 16037 7936
rect 15896 7896 15902 7908
rect 16025 7905 16037 7908
rect 16071 7905 16083 7939
rect 16316 7936 16344 7976
rect 16387 7967 16396 8013
rect 16448 8004 16454 8016
rect 16574 8004 16580 8016
rect 16448 7976 16580 8004
rect 16390 7964 16396 7967
rect 16448 7964 16454 7976
rect 16574 7964 16580 7976
rect 16632 7964 16638 8016
rect 17497 8007 17555 8013
rect 17497 8004 17509 8007
rect 17144 7976 17509 8004
rect 17144 7936 17172 7976
rect 17497 7973 17509 7976
rect 17543 7973 17555 8007
rect 17497 7967 17555 7973
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18094 8007 18152 8013
rect 18094 8004 18106 8007
rect 17920 7976 18106 8004
rect 17920 7964 17926 7976
rect 18094 7973 18106 7976
rect 18140 7973 18152 8007
rect 18094 7967 18152 7973
rect 19659 8007 19717 8013
rect 19659 7973 19671 8007
rect 19705 8004 19717 8007
rect 19978 8004 19984 8016
rect 19705 7976 19984 8004
rect 19705 7973 19717 7976
rect 19659 7967 19717 7973
rect 19978 7964 19984 7976
rect 20036 7964 20042 8016
rect 20990 8004 20996 8016
rect 20951 7976 20996 8004
rect 20990 7964 20996 7976
rect 21048 7964 21054 8016
rect 21100 8013 21128 8044
rect 21085 8007 21143 8013
rect 21085 7973 21097 8007
rect 21131 7973 21143 8007
rect 21085 7967 21143 7973
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 16316 7908 17172 7936
rect 17236 7908 18705 7936
rect 16025 7899 16083 7905
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 6788 7840 9689 7868
rect 6788 7828 6794 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 9677 7831 9735 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 14182 7868 14188 7880
rect 11204 7840 13400 7868
rect 14143 7840 14188 7868
rect 11204 7828 11210 7840
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 6972 7772 7113 7800
rect 6972 7760 6978 7772
rect 7101 7769 7113 7772
rect 7147 7800 7159 7803
rect 11054 7800 11060 7812
rect 7147 7772 11060 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 12253 7803 12311 7809
rect 12253 7800 12265 7803
rect 11388 7772 12265 7800
rect 11388 7760 11394 7772
rect 12253 7769 12265 7772
rect 12299 7769 12311 7803
rect 12253 7763 12311 7769
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 12584 7772 13277 7800
rect 12584 7760 12590 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 13372 7800 13400 7840
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 17236 7877 17264 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 17221 7871 17279 7877
rect 17221 7868 17233 7871
rect 16632 7840 17233 7868
rect 16632 7828 16638 7840
rect 17221 7837 17233 7840
rect 17267 7837 17279 7871
rect 17221 7831 17279 7837
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7868 17555 7871
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17543 7840 17785 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 17773 7837 17785 7840
rect 17819 7868 17831 7871
rect 18046 7868 18052 7880
rect 17819 7840 18052 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18708 7868 18736 7899
rect 19426 7896 19432 7948
rect 19484 7936 19490 7948
rect 19572 7939 19630 7945
rect 19572 7936 19584 7939
rect 19484 7908 19584 7936
rect 19484 7896 19490 7908
rect 19572 7905 19584 7908
rect 19618 7936 19630 7939
rect 20438 7936 20444 7948
rect 19618 7908 20444 7936
rect 19618 7905 19630 7908
rect 19572 7899 19630 7905
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 19794 7868 19800 7880
rect 18708 7840 19800 7868
rect 19794 7828 19800 7840
rect 19852 7868 19858 7880
rect 19981 7871 20039 7877
rect 19981 7868 19993 7871
rect 19852 7840 19993 7868
rect 19852 7828 19858 7840
rect 19981 7837 19993 7840
rect 20027 7837 20039 7871
rect 21266 7868 21272 7880
rect 21227 7840 21272 7868
rect 19981 7831 20039 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 13372 7772 13814 7800
rect 13265 7763 13323 7769
rect 7374 7732 7380 7744
rect 6426 7704 7380 7732
rect 6181 7695 6239 7701
rect 7374 7692 7380 7704
rect 7432 7732 7438 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 7432 7704 7481 7732
rect 7432 7692 7438 7704
rect 7469 7701 7481 7704
rect 7515 7732 7527 7735
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7515 7704 7849 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8754 7732 8760 7744
rect 8260 7704 8760 7732
rect 8260 7692 8266 7704
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9122 7732 9128 7744
rect 9035 7704 9128 7732
rect 9122 7692 9128 7704
rect 9180 7732 9186 7744
rect 10134 7732 10140 7744
rect 9180 7704 10140 7732
rect 9180 7692 9186 7704
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10502 7732 10508 7744
rect 10463 7704 10508 7732
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 11882 7732 11888 7744
rect 11843 7704 11888 7732
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 13081 7735 13139 7741
rect 13081 7701 13093 7735
rect 13127 7732 13139 7735
rect 13446 7732 13452 7744
rect 13127 7704 13452 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13786 7732 13814 7772
rect 14246 7772 17601 7800
rect 14246 7732 14274 7772
rect 17589 7769 17601 7772
rect 17635 7769 17647 7803
rect 17589 7763 17647 7769
rect 13786 7704 14274 7732
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 14642 7732 14648 7744
rect 14599 7704 14648 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 14826 7732 14832 7744
rect 14787 7704 14832 7732
rect 14826 7692 14832 7704
rect 14884 7692 14890 7744
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 14976 7704 15485 7732
rect 14976 7692 14982 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15930 7732 15936 7744
rect 15891 7704 15936 7732
rect 15473 7695 15531 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 18969 7735 19027 7741
rect 18969 7732 18981 7735
rect 18840 7704 18981 7732
rect 18840 7692 18846 7704
rect 18969 7701 18981 7704
rect 19015 7701 19027 7735
rect 19334 7732 19340 7744
rect 19295 7704 19340 7732
rect 18969 7695 19027 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 20717 7735 20775 7741
rect 20717 7701 20729 7735
rect 20763 7732 20775 7735
rect 21266 7732 21272 7744
rect 20763 7704 21272 7732
rect 20763 7701 20775 7704
rect 20717 7695 20775 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 21726 7692 21732 7744
rect 21784 7732 21790 7744
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 21784 7704 21925 7732
rect 21784 7692 21790 7704
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 22278 7732 22284 7744
rect 22239 7704 22284 7732
rect 21913 7695 21971 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 2406 7528 2412 7540
rect 2367 7500 2412 7528
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 2593 7531 2651 7537
rect 2593 7497 2605 7531
rect 2639 7528 2651 7531
rect 3234 7528 3240 7540
rect 2639 7500 3240 7528
rect 2639 7497 2651 7500
rect 2593 7491 2651 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 5350 7528 5356 7540
rect 4264 7500 5356 7528
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 4154 7460 4160 7472
rect 2087 7432 4160 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 4154 7420 4160 7432
rect 4212 7420 4218 7472
rect 1210 7352 1216 7404
rect 1268 7392 1274 7404
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 1268 7364 1501 7392
rect 1268 7352 1274 7364
rect 1489 7361 1501 7364
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 2958 7392 2964 7404
rect 1636 7364 2964 7392
rect 1636 7352 1642 7364
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3970 7392 3976 7404
rect 3931 7364 3976 7392
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4264 7392 4292 7500
rect 5350 7488 5356 7500
rect 5408 7528 5414 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5408 7500 5549 7528
rect 5408 7488 5414 7500
rect 5537 7497 5549 7500
rect 5583 7528 5595 7531
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5583 7500 6469 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7282 7528 7288 7540
rect 6972 7500 7288 7528
rect 6972 7488 6978 7500
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7742 7528 7748 7540
rect 7703 7500 7748 7528
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 8478 7528 8484 7540
rect 8343 7500 8484 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 8478 7488 8484 7500
rect 8536 7528 8542 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 8536 7500 9597 7528
rect 8536 7488 8542 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9585 7491 9643 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 10134 7488 10140 7500
rect 10192 7528 10198 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 10192 7500 10241 7528
rect 10192 7488 10198 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 10229 7491 10287 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 15749 7531 15807 7537
rect 13955 7500 15240 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 6638 7460 6644 7472
rect 4396 7432 6644 7460
rect 4396 7420 4402 7432
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 7558 7420 7564 7472
rect 7616 7460 7622 7472
rect 10042 7460 10048 7472
rect 7616 7432 10048 7460
rect 7616 7420 7622 7432
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 11517 7463 11575 7469
rect 10520 7432 11468 7460
rect 6730 7392 6736 7404
rect 4264 7364 4384 7392
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2314 7324 2320 7336
rect 2271 7296 2320 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 1670 7256 1676 7268
rect 1627 7228 1676 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 1596 7188 1624 7219
rect 1670 7216 1676 7228
rect 1728 7216 1734 7268
rect 2682 7216 2688 7268
rect 2740 7256 2746 7268
rect 2869 7259 2927 7265
rect 2869 7256 2881 7259
rect 2740 7228 2881 7256
rect 2740 7216 2746 7228
rect 2869 7225 2881 7228
rect 2915 7225 2927 7259
rect 2869 7219 2927 7225
rect 2961 7259 3019 7265
rect 2961 7225 2973 7259
rect 3007 7256 3019 7259
rect 3050 7256 3056 7268
rect 3007 7228 3056 7256
rect 3007 7225 3019 7228
rect 2961 7219 3019 7225
rect 992 7160 1624 7188
rect 992 7148 998 7160
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 2593 7191 2651 7197
rect 2593 7188 2605 7191
rect 2372 7160 2605 7188
rect 2372 7148 2378 7160
rect 2593 7157 2605 7160
rect 2639 7157 2651 7191
rect 2884 7188 2912 7219
rect 3050 7216 3056 7228
rect 3108 7216 3114 7268
rect 3697 7259 3755 7265
rect 3697 7225 3709 7259
rect 3743 7225 3755 7259
rect 3697 7219 3755 7225
rect 3789 7259 3847 7265
rect 3789 7225 3801 7259
rect 3835 7256 3847 7259
rect 4356 7256 4384 7364
rect 3835 7228 4384 7256
rect 4632 7364 6736 7392
rect 4632 7256 4660 7364
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7650 7392 7656 7404
rect 6871 7364 7656 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 10520 7392 10548 7432
rect 8803 7364 10548 7392
rect 10597 7395 10655 7401
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 10870 7392 10876 7404
rect 10643 7364 10876 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11440 7392 11468 7432
rect 11517 7429 11529 7463
rect 11563 7460 11575 7463
rect 14642 7460 14648 7472
rect 11563 7432 14648 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 13722 7392 13728 7404
rect 11440 7364 13728 7392
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15212 7401 15240 7500
rect 15749 7497 15761 7531
rect 15795 7528 15807 7531
rect 15838 7528 15844 7540
rect 15795 7500 15844 7528
rect 15795 7497 15807 7500
rect 15749 7491 15807 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16117 7531 16175 7537
rect 16117 7497 16129 7531
rect 16163 7528 16175 7531
rect 16390 7528 16396 7540
rect 16163 7500 16396 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17310 7528 17316 7540
rect 16500 7500 17316 7528
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15562 7392 15568 7404
rect 15243 7364 15568 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 16500 7401 16528 7500
rect 17310 7488 17316 7500
rect 17368 7528 17374 7540
rect 20070 7528 20076 7540
rect 17368 7500 20076 7528
rect 17368 7488 17374 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20864 7500 20913 7528
rect 20864 7488 20870 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 20901 7491 20959 7497
rect 17037 7463 17095 7469
rect 17037 7429 17049 7463
rect 17083 7460 17095 7463
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 17083 7432 18797 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 18785 7429 18797 7432
rect 18831 7460 18843 7463
rect 19058 7460 19064 7472
rect 18831 7432 19064 7460
rect 18831 7429 18843 7432
rect 18785 7423 18843 7429
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 20349 7463 20407 7469
rect 20349 7460 20361 7463
rect 19300 7432 20361 7460
rect 19300 7420 19306 7432
rect 20349 7429 20361 7432
rect 20395 7460 20407 7463
rect 20622 7460 20628 7472
rect 20395 7432 20628 7460
rect 20395 7429 20407 7432
rect 20349 7423 20407 7429
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 21453 7463 21511 7469
rect 21453 7429 21465 7463
rect 21499 7460 21511 7463
rect 23566 7460 23572 7472
rect 21499 7432 23572 7460
rect 21499 7429 21511 7432
rect 21453 7423 21511 7429
rect 23566 7420 23572 7432
rect 23624 7420 23630 7472
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 19978 7392 19984 7404
rect 18279 7364 19984 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 23198 7392 23204 7404
rect 20312 7364 23204 7392
rect 20312 7352 20318 7364
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 6178 7324 6184 7336
rect 5491 7296 6184 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 6840 7296 8309 7324
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4632 7228 4813 7256
rect 3835 7225 3847 7228
rect 3789 7219 3847 7225
rect 4801 7225 4813 7228
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5074 7256 5080 7268
rect 4939 7228 5080 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 3234 7188 3240 7200
rect 2884 7160 3240 7188
rect 2593 7151 2651 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 3602 7148 3608 7200
rect 3660 7188 3666 7200
rect 3712 7188 3740 7219
rect 5074 7216 5080 7228
rect 5132 7256 5138 7268
rect 5534 7256 5540 7268
rect 5132 7228 5540 7256
rect 5132 7216 5138 7228
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 5629 7259 5687 7265
rect 5629 7225 5641 7259
rect 5675 7256 5687 7259
rect 6840 7256 6868 7296
rect 8297 7293 8309 7296
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9585 7327 9643 7333
rect 9456 7296 9501 7324
rect 9456 7284 9462 7296
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 10980 7324 11008 7352
rect 9631 7296 11008 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12400 7296 12449 7324
rect 12400 7284 12406 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 12437 7287 12495 7293
rect 12544 7296 13921 7324
rect 5675 7228 6868 7256
rect 7187 7259 7245 7265
rect 5675 7225 5687 7228
rect 5629 7219 5687 7225
rect 7187 7225 7199 7259
rect 7233 7256 7245 7259
rect 7374 7256 7380 7268
rect 7233 7228 7380 7256
rect 7233 7225 7245 7228
rect 7187 7219 7245 7225
rect 7374 7216 7380 7228
rect 7432 7256 7438 7268
rect 8202 7256 8208 7268
rect 7432 7228 8208 7256
rect 7432 7216 7438 7228
rect 8202 7216 8208 7228
rect 8260 7256 8266 7268
rect 8389 7259 8447 7265
rect 8389 7256 8401 7259
rect 8260 7228 8401 7256
rect 8260 7216 8266 7228
rect 8389 7225 8401 7228
rect 8435 7225 8447 7259
rect 8389 7219 8447 7225
rect 8570 7216 8576 7268
rect 8628 7256 8634 7268
rect 8826 7259 8884 7265
rect 8826 7256 8838 7259
rect 8628 7228 8838 7256
rect 8628 7216 8634 7228
rect 8826 7225 8838 7228
rect 8872 7225 8884 7259
rect 8826 7219 8884 7225
rect 10413 7259 10471 7265
rect 10413 7225 10425 7259
rect 10459 7256 10471 7259
rect 10959 7259 11017 7265
rect 10959 7256 10971 7259
rect 10459 7228 10971 7256
rect 10459 7225 10471 7228
rect 10413 7219 10471 7225
rect 10959 7225 10971 7228
rect 11005 7225 11017 7259
rect 10959 7219 11017 7225
rect 3660 7160 3740 7188
rect 3660 7148 3666 7160
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 4488 7160 5733 7188
rect 4488 7148 4494 7160
rect 5721 7157 5733 7160
rect 5767 7157 5779 7191
rect 6086 7188 6092 7200
rect 6047 7160 6092 7188
rect 5721 7151 5779 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 8662 7188 8668 7200
rect 6319 7160 8668 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 10502 7188 10508 7200
rect 10275 7160 10508 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10980 7188 11008 7219
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 12544 7256 12572 7296
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 19426 7324 19432 7336
rect 18932 7296 19432 7324
rect 18932 7284 18938 7296
rect 19426 7284 19432 7296
rect 19484 7324 19490 7336
rect 19521 7327 19579 7333
rect 19521 7324 19533 7327
rect 19484 7296 19533 7324
rect 19484 7284 19490 7296
rect 19521 7293 19533 7296
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 20530 7284 20536 7336
rect 20588 7324 20594 7336
rect 21269 7327 21327 7333
rect 21269 7324 21281 7327
rect 20588 7296 21281 7324
rect 20588 7284 20594 7296
rect 21269 7293 21281 7296
rect 21315 7324 21327 7327
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21315 7296 21833 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 12799 7259 12857 7265
rect 12799 7256 12811 7259
rect 11112 7228 12572 7256
rect 11112 7216 11118 7228
rect 12774 7225 12811 7256
rect 12845 7256 12857 7259
rect 14274 7256 14280 7268
rect 12845 7228 14280 7256
rect 12845 7225 12857 7228
rect 12774 7219 12857 7225
rect 11422 7188 11428 7200
rect 10980 7160 11428 7188
rect 11422 7148 11428 7160
rect 11480 7188 11486 7200
rect 12158 7188 12164 7200
rect 11480 7160 12164 7188
rect 11480 7148 11486 7160
rect 12158 7148 12164 7160
rect 12216 7188 12222 7200
rect 12253 7191 12311 7197
rect 12253 7188 12265 7191
rect 12216 7160 12265 7188
rect 12216 7148 12222 7160
rect 12253 7157 12265 7160
rect 12299 7188 12311 7191
rect 12774 7188 12802 7219
rect 14274 7216 14280 7228
rect 14332 7216 14338 7268
rect 14642 7216 14648 7268
rect 14700 7256 14706 7268
rect 14700 7228 14745 7256
rect 14700 7216 14706 7228
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 18322 7256 18328 7268
rect 16632 7228 16677 7256
rect 17420 7228 18328 7256
rect 16632 7216 16638 7228
rect 13354 7188 13360 7200
rect 12299 7160 12802 7188
rect 13315 7160 13360 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14093 7191 14151 7197
rect 14093 7188 14105 7191
rect 13872 7160 14105 7188
rect 13872 7148 13878 7160
rect 14093 7157 14105 7160
rect 14139 7188 14151 7191
rect 15562 7188 15568 7200
rect 14139 7160 15568 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 17420 7197 17448 7228
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 19058 7216 19064 7268
rect 19116 7256 19122 7268
rect 19797 7259 19855 7265
rect 19797 7256 19809 7259
rect 19116 7228 19809 7256
rect 19116 7216 19122 7228
rect 19797 7225 19809 7228
rect 19843 7225 19855 7259
rect 19797 7219 19855 7225
rect 19886 7216 19892 7268
rect 19944 7256 19950 7268
rect 19944 7228 19989 7256
rect 19944 7216 19950 7228
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16908 7160 17417 7188
rect 16908 7148 16914 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17770 7188 17776 7200
rect 17731 7160 17776 7188
rect 17405 7151 17463 7157
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 18012 7160 19165 7188
rect 18012 7148 18018 7160
rect 19153 7157 19165 7160
rect 19199 7157 19211 7191
rect 19153 7151 19211 7157
rect 21910 7148 21916 7200
rect 21968 7188 21974 7200
rect 22189 7191 22247 7197
rect 22189 7188 22201 7191
rect 21968 7160 22201 7188
rect 21968 7148 21974 7160
rect 22189 7157 22201 7160
rect 22235 7157 22247 7191
rect 22189 7151 22247 7157
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 2409 6987 2467 6993
rect 2409 6953 2421 6987
rect 2455 6984 2467 6987
rect 2498 6984 2504 6996
rect 2455 6956 2504 6984
rect 2455 6953 2467 6956
rect 2409 6947 2467 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 3418 6984 3424 6996
rect 2976 6956 3424 6984
rect 2976 6928 3004 6956
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 3970 6984 3976 6996
rect 3671 6956 3976 6984
rect 1851 6919 1909 6925
rect 1851 6885 1863 6919
rect 1897 6916 1909 6919
rect 2038 6916 2044 6928
rect 1897 6888 2044 6916
rect 1897 6885 1909 6888
rect 1851 6879 1909 6885
rect 2038 6876 2044 6888
rect 2096 6876 2102 6928
rect 2685 6919 2743 6925
rect 2685 6885 2697 6919
rect 2731 6916 2743 6919
rect 2958 6916 2964 6928
rect 2731 6888 2964 6916
rect 2731 6885 2743 6888
rect 2685 6879 2743 6885
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 3234 6916 3240 6928
rect 3147 6888 3240 6916
rect 3234 6876 3240 6888
rect 3292 6916 3298 6928
rect 3671 6916 3699 6956
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 4065 6987 4123 6993
rect 4065 6953 4077 6987
rect 4111 6984 4123 6987
rect 4982 6984 4988 6996
rect 4111 6956 4521 6984
rect 4111 6953 4123 6956
rect 4065 6947 4123 6953
rect 4338 6916 4344 6928
rect 3292 6888 4344 6916
rect 3292 6876 3298 6888
rect 3671 6857 3699 6888
rect 4338 6876 4344 6888
rect 4396 6876 4402 6928
rect 4493 6925 4521 6956
rect 4908 6956 4988 6984
rect 4478 6919 4536 6925
rect 4478 6885 4490 6919
rect 4524 6885 4536 6919
rect 4908 6916 4936 6956
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6822 6984 6828 6996
rect 5592 6956 6828 6984
rect 5592 6944 5598 6956
rect 4478 6879 4536 6885
rect 4586 6888 5028 6916
rect 201 6851 259 6857
rect 201 6817 213 6851
rect 247 6848 259 6851
rect 1489 6851 1547 6857
rect 1489 6848 1501 6851
rect 247 6820 1501 6848
rect 247 6817 259 6820
rect 201 6811 259 6817
rect 1489 6817 1501 6820
rect 1535 6817 1547 6851
rect 1489 6811 1547 6817
rect 3380 6851 3438 6857
rect 3380 6817 3392 6851
rect 3426 6848 3438 6851
rect 3656 6851 3714 6857
rect 3426 6820 3602 6848
rect 3426 6817 3438 6820
rect 3380 6811 3438 6817
rect 1504 6780 1532 6811
rect 1854 6780 1860 6792
rect 1504 6752 1860 6780
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 2406 6740 2412 6792
rect 2464 6780 2470 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 2464 6752 2605 6780
rect 2464 6740 2470 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 3467 6783 3525 6789
rect 3467 6780 3479 6783
rect 2593 6743 2651 6749
rect 2745 6752 3479 6780
rect 661 6715 719 6721
rect 661 6681 673 6715
rect 707 6712 719 6715
rect 2745 6712 2773 6752
rect 3467 6749 3479 6752
rect 3513 6749 3525 6783
rect 3574 6780 3602 6820
rect 3656 6817 3668 6851
rect 3702 6817 3714 6851
rect 3878 6848 3884 6860
rect 3656 6811 3714 6817
rect 3747 6820 3884 6848
rect 3747 6780 3775 6820
rect 3878 6808 3884 6820
rect 3936 6848 3942 6860
rect 4586 6848 4614 6888
rect 3936 6820 4016 6848
rect 3936 6808 3942 6820
rect 3574 6752 3775 6780
rect 3988 6780 4016 6820
rect 4126 6820 4614 6848
rect 4126 6780 4154 6820
rect 3988 6752 4154 6780
rect 4157 6783 4215 6789
rect 3467 6743 3525 6749
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4203 6752 4292 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4264 6712 4292 6752
rect 4908 6712 4936 6888
rect 5000 6848 5028 6888
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 5994 6916 6000 6928
rect 5408 6888 6000 6916
rect 5408 6876 5414 6888
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 6104 6925 6132 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7282 6984 7288 6996
rect 7243 6956 7288 6984
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 8202 6984 8208 6996
rect 8163 6956 8208 6984
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 11057 6987 11115 6993
rect 11057 6984 11069 6987
rect 8720 6956 11069 6984
rect 8720 6944 8726 6956
rect 11057 6953 11069 6956
rect 11103 6953 11115 6987
rect 12158 6984 12164 6996
rect 12119 6956 12164 6984
rect 11057 6947 11115 6953
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 13538 6944 13544 6996
rect 13596 6984 13602 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 13596 6956 14657 6984
rect 13596 6944 13602 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 15010 6984 15016 6996
rect 14971 6956 15016 6984
rect 14645 6947 14703 6953
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 16301 6987 16359 6993
rect 16301 6953 16313 6987
rect 16347 6984 16359 6987
rect 16482 6984 16488 6996
rect 16347 6956 16488 6984
rect 16347 6953 16359 6956
rect 16301 6947 16359 6953
rect 16482 6944 16488 6956
rect 16540 6984 16546 6996
rect 17678 6984 17684 6996
rect 16540 6956 17684 6984
rect 16540 6944 16546 6956
rect 17678 6944 17684 6956
rect 17736 6944 17742 6996
rect 17865 6987 17923 6993
rect 17865 6953 17877 6987
rect 17911 6984 17923 6987
rect 18046 6984 18052 6996
rect 17911 6956 18052 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 19153 6987 19211 6993
rect 19153 6984 19165 6987
rect 18380 6956 19165 6984
rect 18380 6944 18386 6956
rect 19153 6953 19165 6956
rect 19199 6953 19211 6987
rect 19153 6947 19211 6953
rect 19797 6987 19855 6993
rect 19797 6953 19809 6987
rect 19843 6984 19855 6987
rect 19886 6984 19892 6996
rect 19843 6956 19892 6984
rect 19843 6953 19855 6956
rect 19797 6947 19855 6953
rect 19886 6944 19892 6956
rect 19944 6944 19950 6996
rect 6089 6919 6147 6925
rect 6089 6885 6101 6919
rect 6135 6885 6147 6919
rect 6638 6916 6644 6928
rect 6599 6888 6644 6916
rect 6089 6879 6147 6885
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 6733 6919 6791 6925
rect 6733 6885 6745 6919
rect 6779 6916 6791 6919
rect 7650 6916 7656 6928
rect 6779 6888 7656 6916
rect 6779 6885 6791 6888
rect 6733 6879 6791 6885
rect 7650 6876 7656 6888
rect 7708 6916 7714 6928
rect 8386 6916 8392 6928
rect 7708 6888 8392 6916
rect 7708 6876 7714 6888
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 8754 6876 8760 6928
rect 8812 6916 8818 6928
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 8812 6888 9873 6916
rect 8812 6876 8818 6888
rect 9861 6885 9873 6888
rect 9907 6916 9919 6919
rect 11146 6916 11152 6928
rect 9907 6888 11152 6916
rect 9907 6885 9919 6888
rect 9861 6879 9919 6885
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 13446 6876 13452 6928
rect 13504 6916 13510 6928
rect 13725 6919 13783 6925
rect 13725 6916 13737 6919
rect 13504 6888 13737 6916
rect 13504 6876 13510 6888
rect 13725 6885 13737 6888
rect 13771 6885 13783 6919
rect 13725 6879 13783 6885
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 13872 6888 13917 6916
rect 13872 6876 13878 6888
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15102 6916 15108 6928
rect 14424 6888 15108 6916
rect 14424 6876 14430 6888
rect 15102 6876 15108 6888
rect 15160 6916 15166 6928
rect 15749 6919 15807 6925
rect 15749 6916 15761 6919
rect 15160 6888 15761 6916
rect 15160 6876 15166 6888
rect 15749 6885 15761 6888
rect 15795 6885 15807 6919
rect 15749 6879 15807 6885
rect 16390 6876 16396 6928
rect 16448 6916 16454 6928
rect 16806 6919 16864 6925
rect 16806 6916 16818 6919
rect 16448 6888 16818 6916
rect 16448 6876 16454 6888
rect 16806 6885 16818 6888
rect 16852 6916 16864 6919
rect 17770 6916 17776 6928
rect 16852 6888 17776 6916
rect 16852 6885 16864 6888
rect 16806 6879 16864 6885
rect 17770 6876 17776 6888
rect 17828 6916 17834 6928
rect 18554 6919 18612 6925
rect 18554 6916 18566 6919
rect 17828 6888 18566 6916
rect 17828 6876 17834 6888
rect 18554 6885 18566 6888
rect 18600 6916 18612 6919
rect 19058 6916 19064 6928
rect 18600 6888 19064 6916
rect 18600 6885 18612 6888
rect 18554 6879 18612 6885
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 20806 6876 20812 6928
rect 20864 6916 20870 6928
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 20864 6888 21097 6916
rect 20864 6876 20870 6888
rect 21085 6885 21097 6888
rect 21131 6885 21143 6919
rect 21085 6879 21143 6885
rect 7837 6851 7895 6857
rect 5000 6820 5856 6848
rect 4982 6740 4988 6792
rect 5040 6780 5046 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5040 6752 5733 6780
rect 5040 6740 5046 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5828 6780 5856 6820
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 7926 6848 7932 6860
rect 7883 6820 7932 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8260 6820 9045 6848
rect 8260 6808 8266 6820
rect 9033 6817 9045 6820
rect 9079 6848 9091 6851
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9079 6820 9321 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9309 6817 9321 6820
rect 9355 6848 9367 6851
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 9355 6820 9413 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10560 6820 10793 6848
rect 10560 6808 10566 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 11793 6851 11851 6857
rect 11793 6817 11805 6851
rect 11839 6848 11851 6851
rect 11974 6848 11980 6860
rect 11839 6820 11980 6848
rect 11839 6817 11851 6820
rect 11793 6811 11851 6817
rect 11974 6808 11980 6820
rect 12032 6848 12038 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 12032 6820 13369 6848
rect 12032 6808 12038 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 15356 6851 15414 6857
rect 15356 6817 15368 6851
rect 15402 6817 15414 6851
rect 15356 6811 15414 6817
rect 8478 6780 8484 6792
rect 5828 6752 8484 6780
rect 5721 6743 5779 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9640 6752 9781 6780
rect 9640 6740 9646 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 10226 6780 10232 6792
rect 10187 6752 10232 6780
rect 9769 6743 9827 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 13538 6780 13544 6792
rect 10744 6752 13544 6780
rect 10744 6740 10750 6752
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 13998 6780 14004 6792
rect 13872 6752 14004 6780
rect 13872 6740 13878 6752
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 5074 6712 5080 6724
rect 707 6684 2773 6712
rect 4080 6684 4936 6712
rect 5035 6684 5080 6712
rect 707 6681 719 6684
rect 661 6675 719 6681
rect 293 6647 351 6653
rect 293 6613 305 6647
rect 339 6644 351 6647
rect 3234 6644 3240 6656
rect 339 6616 3240 6644
rect 339 6613 351 6616
rect 293 6607 351 6613
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3743 6647 3801 6653
rect 3743 6613 3755 6647
rect 3789 6644 3801 6647
rect 3878 6644 3884 6656
rect 3789 6616 3884 6644
rect 3789 6613 3801 6616
rect 3743 6607 3801 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4080 6653 4108 6684
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 4028 6616 4077 6644
rect 4028 6604 4034 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4264 6644 4292 6684
rect 5074 6672 5080 6684
rect 5132 6672 5138 6724
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 5684 6684 6745 6712
rect 5684 6672 5690 6684
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 6733 6675 6791 6681
rect 6822 6672 6828 6724
rect 6880 6712 6886 6724
rect 8294 6712 8300 6724
rect 6880 6684 8300 6712
rect 6880 6672 6886 6684
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 10134 6712 10140 6724
rect 8803 6684 10140 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 11020 6684 12725 6712
rect 11020 6672 11026 6684
rect 12713 6681 12725 6684
rect 12759 6712 12771 6715
rect 12989 6715 13047 6721
rect 12989 6712 13001 6715
rect 12759 6684 13001 6712
rect 12759 6681 12771 6684
rect 12713 6675 12771 6681
rect 12989 6681 13001 6684
rect 13035 6681 13047 6715
rect 12989 6675 13047 6681
rect 15010 6672 15016 6724
rect 15068 6712 15074 6724
rect 15371 6712 15399 6811
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 16080 6820 20453 6848
rect 16080 6808 16086 6820
rect 20441 6817 20453 6820
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 16482 6780 16488 6792
rect 16443 6752 16488 6780
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17828 6752 18245 6780
rect 17828 6740 17834 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20772 6752 21005 6780
rect 20772 6740 20778 6752
rect 20993 6749 21005 6752
rect 21039 6780 21051 6783
rect 21913 6783 21971 6789
rect 21913 6780 21925 6783
rect 21039 6752 21925 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21913 6749 21925 6752
rect 21959 6749 21971 6783
rect 21913 6743 21971 6749
rect 15068 6684 15399 6712
rect 17405 6715 17463 6721
rect 15068 6672 15074 6684
rect 17405 6681 17417 6715
rect 17451 6712 17463 6715
rect 17451 6684 18137 6712
rect 17451 6681 17463 6684
rect 17405 6675 17463 6681
rect 4212 6616 4292 6644
rect 4212 6604 4218 6616
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5353 6647 5411 6653
rect 5353 6644 5365 6647
rect 4764 6616 5365 6644
rect 4764 6604 4770 6616
rect 5353 6613 5365 6616
rect 5399 6613 5411 6647
rect 5353 6607 5411 6613
rect 6086 6604 6092 6656
rect 6144 6644 6150 6656
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 6144 6616 6929 6644
rect 6144 6604 6150 6616
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 7834 6644 7840 6656
rect 7791 6616 7840 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 9309 6647 9367 6653
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 10686 6644 10692 6656
rect 9355 6616 10692 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10928 6616 11437 6644
rect 10928 6604 10934 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11882 6644 11888 6656
rect 11572 6616 11888 6644
rect 11572 6604 11578 6616
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 15286 6644 15292 6656
rect 13780 6616 15292 6644
rect 13780 6604 13786 6616
rect 15286 6604 15292 6616
rect 15344 6644 15350 6656
rect 15427 6647 15485 6653
rect 15427 6644 15439 6647
rect 15344 6616 15439 6644
rect 15344 6604 15350 6616
rect 15427 6613 15439 6616
rect 15473 6613 15485 6647
rect 18109 6644 18137 6684
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 21545 6715 21603 6721
rect 21545 6712 21557 6715
rect 19668 6684 21557 6712
rect 19668 6672 19674 6684
rect 21545 6681 21557 6684
rect 21591 6712 21603 6715
rect 21634 6712 21640 6724
rect 21591 6684 21640 6712
rect 21591 6681 21603 6684
rect 21545 6675 21603 6681
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 18230 6644 18236 6656
rect 18109 6616 18236 6644
rect 15427 6607 15485 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 20070 6644 20076 6656
rect 20031 6616 20076 6644
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 22152 6616 22293 6644
rect 22152 6604 22158 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 750 6400 756 6452
rect 808 6440 814 6452
rect 1811 6443 1869 6449
rect 1811 6440 1823 6443
rect 808 6412 1823 6440
rect 808 6400 814 6412
rect 1811 6409 1823 6412
rect 1857 6440 1869 6443
rect 2406 6440 2412 6452
rect 1857 6412 2412 6440
rect 1857 6409 1869 6412
rect 1811 6403 1869 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 3050 6440 3056 6452
rect 3011 6412 3056 6440
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 4939 6443 4997 6449
rect 4939 6440 4951 6443
rect 3757 6412 4951 6440
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 1535 6375 1593 6381
rect 1535 6372 1547 6375
rect 1452 6344 1547 6372
rect 1452 6332 1458 6344
rect 1535 6341 1547 6344
rect 1581 6341 1593 6375
rect 2590 6372 2596 6384
rect 1535 6335 1593 6341
rect 1826 6344 2596 6372
rect 1826 6304 1854 6344
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 2682 6332 2688 6384
rect 2740 6372 2746 6384
rect 3757 6372 3785 6412
rect 4939 6409 4951 6412
rect 4985 6409 4997 6443
rect 5626 6440 5632 6452
rect 4939 6403 4997 6409
rect 5138 6412 5632 6440
rect 5138 6384 5166 6412
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6270 6440 6276 6452
rect 6052 6412 6276 6440
rect 6052 6400 6058 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6963 6443 7021 6449
rect 6963 6409 6975 6443
rect 7009 6440 7021 6443
rect 7098 6440 7104 6452
rect 7009 6412 7104 6440
rect 7009 6409 7021 6412
rect 6963 6403 7021 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 9306 6440 9312 6452
rect 8343 6412 9312 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 12250 6440 12256 6452
rect 12211 6412 12256 6440
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12618 6440 12624 6452
rect 12579 6412 12624 6440
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 13446 6440 13452 6452
rect 12851 6412 13452 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13538 6400 13544 6452
rect 13596 6440 13602 6452
rect 13998 6440 14004 6452
rect 13596 6412 14004 6440
rect 13596 6400 13602 6412
rect 13998 6400 14004 6412
rect 14056 6440 14062 6452
rect 14921 6443 14979 6449
rect 14921 6440 14933 6443
rect 14056 6412 14933 6440
rect 14056 6400 14062 6412
rect 14921 6409 14933 6412
rect 14967 6440 14979 6443
rect 15010 6440 15016 6452
rect 14967 6412 15016 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16485 6443 16543 6449
rect 16485 6440 16497 6443
rect 16448 6412 16497 6440
rect 16448 6400 16454 6412
rect 16485 6409 16497 6412
rect 16531 6409 16543 6443
rect 16485 6403 16543 6409
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17770 6440 17776 6452
rect 16632 6412 17776 6440
rect 16632 6400 16638 6412
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18506 6400 18512 6452
rect 18564 6440 18570 6452
rect 18690 6440 18696 6452
rect 18564 6412 18696 6440
rect 18564 6400 18570 6412
rect 18690 6400 18696 6412
rect 18748 6440 18754 6452
rect 18748 6412 20300 6440
rect 18748 6400 18754 6412
rect 2740 6344 3785 6372
rect 2740 6332 2746 6344
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 5074 6332 5080 6384
rect 5132 6344 5166 6384
rect 5810 6372 5816 6384
rect 5460 6344 5816 6372
rect 5132 6332 5138 6344
rect 1479 6276 1854 6304
rect 2133 6307 2191 6313
rect 1479 6245 1507 6276
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 2222 6304 2228 6316
rect 2179 6276 2228 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3513 6307 3571 6313
rect 3513 6304 3525 6307
rect 2924 6276 3525 6304
rect 2924 6264 2930 6276
rect 3513 6273 3525 6276
rect 3559 6304 3571 6307
rect 3559 6276 3924 6304
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 1464 6239 1522 6245
rect 1464 6205 1476 6239
rect 1510 6205 1522 6239
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1464 6199 1522 6205
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 2038 6168 2044 6180
rect 1912 6140 2044 6168
rect 1912 6128 1918 6140
rect 2038 6128 2044 6140
rect 2096 6168 2102 6180
rect 2454 6171 2512 6177
rect 2454 6168 2466 6171
rect 2096 6140 2466 6168
rect 2096 6128 2102 6140
rect 2454 6137 2466 6140
rect 2500 6137 2512 6171
rect 2454 6131 2512 6137
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 3329 6171 3387 6177
rect 3329 6168 3341 6171
rect 3292 6140 3341 6168
rect 3292 6128 3298 6140
rect 3329 6137 3341 6140
rect 3375 6168 3387 6171
rect 3418 6168 3424 6180
rect 3375 6140 3424 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 3896 6100 3924 6276
rect 3988 6168 4016 6332
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 4488 6276 4911 6304
rect 4488 6264 4494 6276
rect 4883 6245 4911 6276
rect 5460 6245 5488 6344
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 6411 6375 6469 6381
rect 6411 6341 6423 6375
rect 6457 6372 6469 6375
rect 7190 6372 7196 6384
rect 6457 6344 7196 6372
rect 6457 6341 6469 6344
rect 6411 6335 6469 6341
rect 7190 6332 7196 6344
rect 7248 6372 7254 6384
rect 7742 6372 7748 6384
rect 7248 6344 7748 6372
rect 7248 6332 7254 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 13630 6372 13636 6384
rect 7892 6344 13636 6372
rect 7892 6332 7898 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 14274 6332 14280 6384
rect 14332 6372 14338 6384
rect 14553 6375 14611 6381
rect 14553 6372 14565 6375
rect 14332 6344 14565 6372
rect 14332 6332 14338 6344
rect 14553 6341 14565 6344
rect 14599 6341 14611 6375
rect 14553 6335 14611 6341
rect 14642 6332 14648 6384
rect 14700 6372 14706 6384
rect 18874 6372 18880 6384
rect 14700 6344 18880 6372
rect 14700 6332 14706 6344
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 19058 6372 19064 6384
rect 19019 6344 19064 6372
rect 19058 6332 19064 6344
rect 19116 6332 19122 6384
rect 19245 6375 19303 6381
rect 19245 6341 19257 6375
rect 19291 6372 19303 6375
rect 20070 6372 20076 6384
rect 19291 6344 20076 6372
rect 19291 6341 19303 6344
rect 19245 6335 19303 6341
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 20272 6381 20300 6412
rect 20346 6400 20352 6452
rect 20404 6440 20410 6452
rect 21315 6443 21373 6449
rect 21315 6440 21327 6443
rect 20404 6412 21327 6440
rect 20404 6400 20410 6412
rect 21315 6409 21327 6412
rect 21361 6409 21373 6443
rect 21315 6403 21373 6409
rect 21450 6400 21456 6452
rect 21508 6440 21514 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 21508 6412 22385 6440
rect 21508 6400 21514 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 20257 6375 20315 6381
rect 20257 6341 20269 6375
rect 20303 6341 20315 6375
rect 20257 6335 20315 6341
rect 20806 6332 20812 6384
rect 20864 6372 20870 6384
rect 20901 6375 20959 6381
rect 20901 6372 20913 6375
rect 20864 6344 20913 6372
rect 20864 6332 20870 6344
rect 20901 6341 20913 6344
rect 20947 6341 20959 6375
rect 20901 6335 20959 6341
rect 21542 6332 21548 6384
rect 21600 6372 21606 6384
rect 21637 6375 21695 6381
rect 21637 6372 21649 6375
rect 21600 6344 21649 6372
rect 21600 6332 21606 6344
rect 21637 6341 21649 6344
rect 21683 6341 21695 6375
rect 22002 6372 22008 6384
rect 21963 6344 22008 6372
rect 21637 6335 21695 6341
rect 22002 6332 22008 6344
rect 22060 6332 22066 6384
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 5951 6276 7389 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 7377 6273 7389 6276
rect 7423 6304 7435 6307
rect 9398 6304 9404 6316
rect 7423 6276 9404 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 12158 6304 12164 6316
rect 11931 6276 12164 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 13906 6304 13912 6316
rect 12773 6276 13912 6304
rect 4868 6239 4926 6245
rect 4868 6205 4880 6239
rect 4914 6205 4926 6239
rect 4868 6199 4926 6205
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6205 5503 6239
rect 5626 6236 5632 6248
rect 5587 6208 5632 6236
rect 5445 6199 5503 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 6308 6239 6366 6245
rect 6308 6205 6320 6239
rect 6354 6205 6366 6239
rect 6308 6199 6366 6205
rect 6892 6239 6950 6245
rect 6892 6205 6904 6239
rect 6938 6236 6950 6239
rect 7834 6236 7840 6248
rect 6938 6208 7840 6236
rect 6938 6205 6950 6208
rect 6892 6199 6950 6205
rect 4065 6171 4123 6177
rect 4065 6168 4077 6171
rect 3988 6140 4077 6168
rect 4065 6137 4077 6140
rect 4111 6137 4123 6171
rect 4065 6131 4123 6137
rect 4157 6171 4215 6177
rect 4157 6137 4169 6171
rect 4203 6168 4215 6171
rect 4338 6168 4344 6180
rect 4203 6140 4344 6168
rect 4203 6137 4215 6140
rect 4157 6131 4215 6137
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4709 6171 4767 6177
rect 4709 6137 4721 6171
rect 4755 6137 4767 6171
rect 4709 6131 4767 6137
rect 4430 6100 4436 6112
rect 3896 6072 4436 6100
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4724 6100 4752 6131
rect 5626 6100 5632 6112
rect 4672 6072 5632 6100
rect 4672 6060 4678 6072
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6323 6100 6351 6199
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8260 6208 8585 6236
rect 8260 6196 8266 6208
rect 8573 6205 8585 6208
rect 8619 6236 8631 6239
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8619 6208 8953 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12773 6236 12801 6276
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 19334 6304 19340 6316
rect 14246 6276 19340 6304
rect 14246 6236 14274 6276
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 15102 6236 15108 6248
rect 11848 6208 12801 6236
rect 13648 6208 14274 6236
rect 15063 6208 15108 6236
rect 11848 6196 11854 6208
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 7739 6171 7797 6177
rect 7248 6140 7604 6168
rect 7248 6128 7254 6140
rect 6144 6072 6351 6100
rect 6144 6060 6150 6072
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7466 6100 7472 6112
rect 7340 6072 7472 6100
rect 7340 6060 7346 6072
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7576 6100 7604 6140
rect 7739 6137 7751 6171
rect 7785 6168 7797 6171
rect 8220 6168 8248 6196
rect 9030 6168 9036 6180
rect 7785 6140 8248 6168
rect 8588 6140 9036 6168
rect 7785 6137 7797 6140
rect 7739 6131 7797 6137
rect 8588 6100 8616 6140
rect 9030 6128 9036 6140
rect 9088 6128 9094 6180
rect 9217 6171 9275 6177
rect 9217 6137 9229 6171
rect 9263 6137 9275 6171
rect 9217 6131 9275 6137
rect 7576 6072 8616 6100
rect 9232 6100 9260 6131
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 9861 6171 9919 6177
rect 9364 6140 9409 6168
rect 9364 6128 9370 6140
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 10226 6168 10232 6180
rect 9907 6140 10232 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 10873 6171 10931 6177
rect 10873 6137 10885 6171
rect 10919 6137 10931 6171
rect 10873 6131 10931 6137
rect 9766 6100 9772 6112
rect 9232 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10183 6072 10609 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10597 6069 10609 6072
rect 10643 6100 10655 6103
rect 10686 6100 10692 6112
rect 10643 6072 10692 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10888 6100 10916 6131
rect 10962 6128 10968 6180
rect 11020 6168 11026 6180
rect 11020 6140 11065 6168
rect 11020 6128 11026 6140
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11204 6140 11529 6168
rect 11204 6128 11210 6140
rect 11517 6137 11529 6140
rect 11563 6168 11575 6171
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 11563 6140 12817 6168
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12986 6168 12992 6180
rect 12947 6140 12992 6168
rect 12805 6131 12863 6137
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 13081 6171 13139 6177
rect 13081 6137 13093 6171
rect 13127 6168 13139 6171
rect 13354 6168 13360 6180
rect 13127 6140 13360 6168
rect 13127 6137 13139 6140
rect 13081 6131 13139 6137
rect 13354 6128 13360 6140
rect 13412 6128 13418 6180
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 13648 6177 13676 6208
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 16920 6239 16978 6245
rect 16920 6205 16932 6239
rect 16966 6236 16978 6239
rect 18785 6239 18843 6245
rect 16966 6208 17448 6236
rect 16966 6205 16978 6208
rect 16920 6199 16978 6205
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 13504 6140 13645 6168
rect 13504 6128 13510 6140
rect 13633 6137 13645 6140
rect 13679 6137 13691 6171
rect 13633 6131 13691 6137
rect 14274 6128 14280 6180
rect 14332 6168 14338 6180
rect 14458 6168 14464 6180
rect 14332 6140 14464 6168
rect 14332 6128 14338 6140
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 15467 6171 15525 6177
rect 15467 6137 15479 6171
rect 15513 6168 15525 6171
rect 16390 6168 16396 6180
rect 15513 6140 16396 6168
rect 15513 6137 15525 6140
rect 15467 6131 15525 6137
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 17420 6177 17448 6208
rect 18785 6205 18797 6239
rect 18831 6236 18843 6239
rect 19242 6236 19248 6248
rect 18831 6208 19248 6236
rect 18831 6205 18843 6208
rect 18785 6199 18843 6205
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 20714 6196 20720 6248
rect 20772 6236 20778 6248
rect 21212 6239 21270 6245
rect 21212 6236 21224 6239
rect 20772 6208 21224 6236
rect 20772 6196 20778 6208
rect 21212 6205 21224 6208
rect 21258 6205 21270 6239
rect 21212 6199 21270 6205
rect 17405 6171 17463 6177
rect 17405 6137 17417 6171
rect 17451 6168 17463 6171
rect 18141 6171 18199 6177
rect 17451 6140 18000 6168
rect 17451 6137 17463 6140
rect 17405 6131 17463 6137
rect 11054 6100 11060 6112
rect 10888 6072 11060 6100
rect 11054 6060 11060 6072
rect 11112 6100 11118 6112
rect 11698 6100 11704 6112
rect 11112 6072 11704 6100
rect 11112 6060 11118 6072
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 13004 6100 13032 6128
rect 12032 6072 13032 6100
rect 13372 6100 13400 6128
rect 13909 6103 13967 6109
rect 13909 6100 13921 6103
rect 13372 6072 13921 6100
rect 12032 6060 12038 6072
rect 13909 6069 13921 6072
rect 13955 6069 13967 6103
rect 16022 6100 16028 6112
rect 15983 6072 16028 6100
rect 13909 6063 13967 6069
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16991 6103 17049 6109
rect 16991 6069 17003 6103
rect 17037 6100 17049 6103
rect 17310 6100 17316 6112
rect 17037 6072 17316 6100
rect 17037 6069 17049 6072
rect 16991 6063 17049 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17972 6100 18000 6140
rect 18141 6137 18153 6171
rect 18187 6137 18199 6171
rect 18141 6131 18199 6137
rect 18046 6100 18052 6112
rect 17972 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18156 6100 18184 6131
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 19518 6168 19524 6180
rect 18288 6140 18333 6168
rect 18937 6140 19524 6168
rect 18288 6128 18294 6140
rect 18414 6100 18420 6112
rect 18156 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 18506 6060 18512 6112
rect 18564 6100 18570 6112
rect 18937 6100 18965 6140
rect 19518 6128 19524 6140
rect 19576 6168 19582 6180
rect 19705 6171 19763 6177
rect 19705 6168 19717 6171
rect 19576 6140 19717 6168
rect 19576 6128 19582 6140
rect 19705 6137 19717 6140
rect 19751 6137 19763 6171
rect 19705 6131 19763 6137
rect 19797 6171 19855 6177
rect 19797 6137 19809 6171
rect 19843 6137 19855 6171
rect 19797 6131 19855 6137
rect 19242 6100 19248 6112
rect 18564 6072 18965 6100
rect 19203 6072 19248 6100
rect 18564 6060 18570 6072
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19426 6100 19432 6112
rect 19387 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6100 19490 6112
rect 19812 6100 19840 6131
rect 19484 6072 19840 6100
rect 19484 6060 19490 6072
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5865 2375 5899
rect 4062 5896 4068 5908
rect 2317 5859 2375 5865
rect 2976 5868 4068 5896
rect 1759 5831 1817 5837
rect 1759 5797 1771 5831
rect 1805 5828 1817 5831
rect 1854 5828 1860 5840
rect 1805 5800 1860 5828
rect 1805 5797 1817 5800
rect 1759 5791 1817 5797
rect 1854 5788 1860 5800
rect 1912 5788 1918 5840
rect 2222 5788 2228 5840
rect 2280 5828 2286 5840
rect 2332 5828 2360 5859
rect 2280 5800 2360 5828
rect 2280 5788 2286 5800
rect 2682 5760 2688 5772
rect 2643 5732 2688 5760
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 2976 5769 3004 5868
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 5067 5868 8125 5896
rect 3142 5788 3148 5840
rect 3200 5828 3206 5840
rect 4338 5828 4344 5840
rect 3200 5800 3786 5828
rect 4299 5800 4344 5828
rect 3200 5788 3206 5800
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5729 3019 5763
rect 3234 5760 3240 5772
rect 3195 5732 3240 5760
rect 2961 5723 3019 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3758 5769 3786 5800
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 4430 5788 4436 5840
rect 4488 5828 4494 5840
rect 4488 5800 4936 5828
rect 4488 5788 4494 5800
rect 3743 5763 3801 5769
rect 3743 5729 3755 5763
rect 3789 5760 3801 5763
rect 4062 5760 4068 5772
rect 3789 5732 4068 5760
rect 3789 5729 3801 5732
rect 3743 5723 3801 5729
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 2866 5692 2872 5704
rect 1443 5664 2872 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3142 5692 3148 5704
rect 3103 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 3896 5664 4261 5692
rect 1762 5584 1768 5636
rect 1820 5624 1826 5636
rect 3375 5627 3433 5633
rect 3375 5624 3387 5627
rect 1820 5596 3387 5624
rect 1820 5584 1826 5596
rect 3375 5593 3387 5596
rect 3421 5593 3433 5627
rect 3375 5587 3433 5593
rect 3694 5584 3700 5636
rect 3752 5624 3758 5636
rect 3896 5624 3924 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 3752 5596 3924 5624
rect 3752 5584 3758 5596
rect 3970 5584 3976 5636
rect 4028 5624 4034 5636
rect 4724 5624 4752 5652
rect 4028 5596 4752 5624
rect 4801 5627 4859 5633
rect 4028 5584 4034 5596
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 4908 5624 4936 5800
rect 5067 5769 5095 5868
rect 8113 5865 8125 5868
rect 8159 5896 8171 5899
rect 8202 5896 8208 5908
rect 8159 5868 8208 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8444 5868 9045 5896
rect 8444 5856 8450 5868
rect 9033 5865 9045 5868
rect 9079 5896 9091 5899
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 9079 5868 9229 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9217 5865 9229 5868
rect 9263 5865 9275 5899
rect 9217 5859 9275 5865
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 13538 5896 13544 5908
rect 10284 5868 13544 5896
rect 10284 5856 10290 5868
rect 5445 5831 5503 5837
rect 5445 5797 5457 5831
rect 5491 5828 5503 5831
rect 5534 5828 5540 5840
rect 5491 5800 5540 5828
rect 5491 5797 5503 5800
rect 5445 5791 5503 5797
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 5994 5828 6000 5840
rect 5955 5800 6000 5828
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 6270 5828 6276 5840
rect 6231 5800 6276 5828
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 6546 5788 6552 5840
rect 6604 5828 6610 5840
rect 9309 5831 9367 5837
rect 9309 5828 9321 5831
rect 6604 5800 9321 5828
rect 6604 5788 6610 5800
rect 9309 5797 9321 5800
rect 9355 5828 9367 5831
rect 9401 5831 9459 5837
rect 9401 5828 9413 5831
rect 9355 5800 9413 5828
rect 9355 5797 9367 5800
rect 9309 5791 9367 5797
rect 9401 5797 9413 5800
rect 9447 5797 9459 5831
rect 9401 5791 9459 5797
rect 9490 5788 9496 5840
rect 9548 5828 9554 5840
rect 9769 5831 9827 5837
rect 9769 5828 9781 5831
rect 9548 5800 9781 5828
rect 9548 5788 9554 5800
rect 9769 5797 9781 5800
rect 9815 5797 9827 5831
rect 9769 5791 9827 5797
rect 9861 5831 9919 5837
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 10152 5828 10180 5856
rect 10428 5837 10456 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 14553 5899 14611 5905
rect 14553 5896 14565 5899
rect 13780 5868 14565 5896
rect 13780 5856 13786 5868
rect 14553 5865 14565 5868
rect 14599 5865 14611 5899
rect 14553 5859 14611 5865
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14792 5868 14933 5896
rect 14792 5856 14798 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 16574 5896 16580 5908
rect 16535 5868 16580 5896
rect 14921 5859 14979 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18230 5896 18236 5908
rect 18187 5868 18236 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 18322 5856 18328 5908
rect 18380 5896 18386 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 18380 5868 19809 5896
rect 18380 5856 18386 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 19797 5859 19855 5865
rect 21358 5856 21364 5908
rect 21416 5896 21422 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21416 5868 21925 5896
rect 21416 5856 21422 5868
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 21913 5859 21971 5865
rect 9907 5800 10180 5828
rect 10413 5831 10471 5837
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10413 5797 10425 5831
rect 10459 5797 10471 5831
rect 10413 5791 10471 5797
rect 10686 5788 10692 5840
rect 10744 5828 10750 5840
rect 10781 5831 10839 5837
rect 10781 5828 10793 5831
rect 10744 5800 10793 5828
rect 10744 5788 10750 5800
rect 10781 5797 10793 5800
rect 10827 5828 10839 5831
rect 11149 5831 11207 5837
rect 11149 5828 11161 5831
rect 10827 5800 11161 5828
rect 10827 5797 10839 5800
rect 10781 5791 10839 5797
rect 11149 5797 11161 5800
rect 11195 5828 11207 5831
rect 11787 5831 11845 5837
rect 11787 5828 11799 5831
rect 11195 5800 11799 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 11787 5797 11799 5800
rect 11833 5828 11845 5831
rect 12158 5828 12164 5840
rect 11833 5800 12164 5828
rect 11833 5797 11845 5800
rect 11787 5791 11845 5797
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12710 5828 12716 5840
rect 12671 5800 12716 5828
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 13357 5831 13415 5837
rect 13357 5797 13369 5831
rect 13403 5828 13415 5831
rect 14182 5828 14188 5840
rect 13403 5800 14188 5828
rect 13403 5797 13415 5800
rect 13357 5791 13415 5797
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 15654 5828 15660 5840
rect 15615 5800 15660 5828
rect 15654 5788 15660 5800
rect 15712 5788 15718 5840
rect 16022 5788 16028 5840
rect 16080 5828 16086 5840
rect 17221 5831 17279 5837
rect 17221 5828 17233 5831
rect 16080 5800 17233 5828
rect 16080 5788 16086 5800
rect 17221 5797 17233 5800
rect 17267 5828 17279 5831
rect 17770 5828 17776 5840
rect 17267 5800 17776 5828
rect 17267 5797 17279 5800
rect 17221 5791 17279 5797
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 18963 5831 19021 5837
rect 18963 5797 18975 5831
rect 19009 5828 19021 5831
rect 19058 5828 19064 5840
rect 19009 5800 19064 5828
rect 19009 5797 19021 5800
rect 18963 5791 19021 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 20496 5800 21097 5828
rect 20496 5788 20502 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21634 5828 21640 5840
rect 21595 5800 21640 5828
rect 21085 5791 21143 5797
rect 21634 5788 21640 5800
rect 21692 5788 21698 5840
rect 5052 5763 5110 5769
rect 5052 5729 5064 5763
rect 5098 5729 5110 5763
rect 5052 5723 5110 5729
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 6914 5760 6920 5772
rect 6871 5732 6920 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7282 5760 7288 5772
rect 7243 5732 7288 5760
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 7650 5760 7656 5772
rect 7607 5732 7656 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 7926 5760 7932 5772
rect 7791 5732 7932 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 10594 5720 10600 5772
rect 10652 5760 10658 5772
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 10652 5732 12357 5760
rect 10652 5720 10658 5732
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 13078 5760 13084 5772
rect 12345 5723 12403 5729
rect 12728 5732 13084 5760
rect 5166 5652 5172 5704
rect 5224 5692 5230 5704
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 5224 5664 5365 5692
rect 5224 5652 5230 5664
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 8846 5692 8852 5704
rect 6227 5664 8852 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9263 5664 9904 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 5994 5624 6000 5636
rect 4847 5596 6000 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 5994 5584 6000 5596
rect 6052 5624 6058 5636
rect 6270 5624 6276 5636
rect 6052 5596 6276 5624
rect 6052 5584 6058 5596
rect 6270 5584 6276 5596
rect 6328 5584 6334 5636
rect 8711 5627 8769 5633
rect 8711 5593 8723 5627
rect 8757 5624 8769 5627
rect 9674 5624 9680 5636
rect 8757 5596 9680 5624
rect 8757 5593 8769 5596
rect 8711 5587 8769 5593
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 9876 5624 9904 5664
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 10008 5664 11437 5692
rect 10008 5652 10014 5664
rect 11425 5661 11437 5664
rect 11471 5692 11483 5695
rect 12728 5692 12756 5732
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13909 5763 13967 5769
rect 13909 5729 13921 5763
rect 13955 5760 13967 5763
rect 15010 5760 15016 5772
rect 13955 5732 15016 5760
rect 13955 5729 13967 5732
rect 13909 5723 13967 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5760 16267 5763
rect 16298 5760 16304 5772
rect 16255 5732 16304 5760
rect 16255 5729 16267 5732
rect 16209 5723 16267 5729
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16540 5732 16896 5760
rect 16540 5720 16546 5732
rect 11471 5664 12756 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12860 5664 13277 5692
rect 12860 5652 12866 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 13504 5664 15577 5692
rect 13504 5652 13510 5664
rect 15565 5661 15577 5664
rect 15611 5692 15623 5695
rect 16758 5692 16764 5704
rect 15611 5664 16764 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 11790 5624 11796 5636
rect 9876 5596 11796 5624
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 12342 5584 12348 5636
rect 12400 5624 12406 5636
rect 12989 5627 13047 5633
rect 12989 5624 13001 5627
rect 12400 5596 13001 5624
rect 12400 5584 12406 5596
rect 12989 5593 13001 5596
rect 13035 5593 13047 5627
rect 12989 5587 13047 5593
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13722 5624 13728 5636
rect 13136 5596 13728 5624
rect 13136 5584 13142 5596
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 14826 5624 14832 5636
rect 14016 5596 14832 5624
rect 753 5559 811 5565
rect 753 5525 765 5559
rect 799 5556 811 5559
rect 3835 5559 3893 5565
rect 3835 5556 3847 5559
rect 799 5528 3847 5556
rect 799 5525 811 5528
rect 753 5519 811 5525
rect 3835 5525 3847 5528
rect 3881 5525 3893 5559
rect 3835 5519 3893 5525
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 5123 5559 5181 5565
rect 5123 5556 5135 5559
rect 4672 5528 5135 5556
rect 4672 5516 4678 5528
rect 5123 5525 5135 5528
rect 5169 5556 5181 5559
rect 6362 5556 6368 5568
rect 5169 5528 6368 5556
rect 5169 5525 5181 5528
rect 5123 5519 5181 5525
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 8386 5556 8392 5568
rect 8347 5528 8392 5556
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9309 5559 9367 5565
rect 9309 5525 9321 5559
rect 9355 5556 9367 5559
rect 10594 5556 10600 5568
rect 9355 5528 10600 5556
rect 9355 5525 9367 5528
rect 9309 5519 9367 5525
rect 10594 5516 10600 5528
rect 10652 5516 10658 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 14016 5556 14044 5596
rect 14826 5584 14832 5596
rect 14884 5624 14890 5636
rect 16868 5624 16896 5732
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 17920 5732 20177 5760
rect 17920 5720 17926 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 17402 5692 17408 5704
rect 17175 5664 17408 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 17494 5652 17500 5704
rect 17552 5692 17558 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 17552 5664 18613 5692
rect 17552 5652 17558 5664
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 19610 5652 19616 5704
rect 19668 5692 19674 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 19668 5664 21005 5692
rect 19668 5652 19674 5664
rect 20993 5661 21005 5664
rect 21039 5692 21051 5695
rect 22094 5692 22100 5704
rect 21039 5664 22100 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 22094 5652 22100 5664
rect 22152 5652 22158 5704
rect 17310 5624 17316 5636
rect 14884 5596 16804 5624
rect 16868 5596 17316 5624
rect 14884 5584 14890 5596
rect 14182 5556 14188 5568
rect 11204 5528 14044 5556
rect 14143 5528 14188 5556
rect 11204 5516 11210 5528
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 16574 5556 16580 5568
rect 15436 5528 16580 5556
rect 15436 5516 15442 5528
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 16776 5556 16804 5596
rect 17310 5584 17316 5596
rect 17368 5624 17374 5636
rect 17678 5624 17684 5636
rect 17368 5596 17684 5624
rect 17368 5584 17374 5596
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 18322 5584 18328 5636
rect 18380 5624 18386 5636
rect 18380 5596 19702 5624
rect 18380 5584 18386 5596
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 16776 5528 18429 5556
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 18966 5516 18972 5568
rect 19024 5556 19030 5568
rect 19150 5556 19156 5568
rect 19024 5528 19156 5556
rect 19024 5516 19030 5528
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 19518 5556 19524 5568
rect 19479 5528 19524 5556
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 19674 5556 19702 5596
rect 20254 5584 20260 5636
rect 20312 5624 20318 5636
rect 22281 5627 22339 5633
rect 22281 5624 22293 5627
rect 20312 5596 22293 5624
rect 20312 5584 20318 5596
rect 22281 5593 22293 5596
rect 22327 5593 22339 5627
rect 22281 5587 22339 5593
rect 20533 5559 20591 5565
rect 20533 5556 20545 5559
rect 19674 5528 20545 5556
rect 20533 5525 20545 5528
rect 20579 5525 20591 5559
rect 20533 5519 20591 5525
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 290 5312 296 5364
rect 348 5352 354 5364
rect 2317 5355 2375 5361
rect 2317 5352 2329 5355
rect 348 5324 2329 5352
rect 348 5312 354 5324
rect 2317 5321 2329 5324
rect 2363 5321 2375 5355
rect 2317 5315 2375 5321
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 9122 5352 9128 5364
rect 3108 5324 9128 5352
rect 3108 5312 3114 5324
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 11471 5355 11529 5361
rect 11471 5321 11483 5355
rect 11517 5352 11529 5355
rect 12802 5352 12808 5364
rect 11517 5324 12808 5352
rect 11517 5321 11529 5324
rect 11471 5315 11529 5321
rect 12802 5312 12808 5324
rect 12860 5312 12866 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 12912 5324 13461 5352
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 3513 5287 3571 5293
rect 3513 5284 3525 5287
rect 2832 5256 3525 5284
rect 2832 5244 2838 5256
rect 3513 5253 3525 5256
rect 3559 5253 3571 5287
rect 5074 5284 5080 5296
rect 3513 5247 3571 5253
rect 4908 5256 5080 5284
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 3142 5216 3148 5228
rect 1443 5188 3148 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 1946 5108 1952 5160
rect 2004 5148 2010 5160
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 2004 5120 2421 5148
rect 2004 5108 2010 5120
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 2498 5108 2504 5160
rect 2556 5148 2562 5160
rect 3234 5148 3240 5160
rect 2556 5120 3240 5148
rect 2556 5108 2562 5120
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3510 5148 3516 5160
rect 3471 5120 3516 5148
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 3970 5148 3976 5160
rect 3883 5120 3976 5148
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 4430 5148 4436 5160
rect 4391 5120 4436 5148
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 4908 5148 4936 5256
rect 5074 5244 5080 5256
rect 5132 5284 5138 5296
rect 5132 5256 5488 5284
rect 5132 5244 5138 5256
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5460 5216 5488 5256
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 5684 5256 6561 5284
rect 5684 5244 5690 5256
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 8570 5284 8576 5296
rect 7524 5256 8576 5284
rect 7524 5244 7530 5256
rect 8570 5244 8576 5256
rect 8628 5284 8634 5296
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8628 5256 9045 5284
rect 8628 5244 8634 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 9033 5247 9091 5253
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 9364 5256 9812 5284
rect 9364 5244 9370 5256
rect 9784 5228 9812 5256
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 10502 5284 10508 5296
rect 9916 5256 10508 5284
rect 9916 5244 9922 5256
rect 10502 5244 10508 5256
rect 10560 5284 10566 5296
rect 11793 5287 11851 5293
rect 11793 5284 11805 5287
rect 10560 5256 11805 5284
rect 10560 5244 10566 5256
rect 7834 5216 7840 5228
rect 5031 5188 7840 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 4847 5120 4936 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 2130 5040 2136 5092
rect 2188 5080 2194 5092
rect 2516 5080 2544 5108
rect 2188 5052 2544 5080
rect 2188 5040 2194 5052
rect 3602 5040 3608 5092
rect 3660 5080 3666 5092
rect 3988 5080 4016 5108
rect 3660 5052 4016 5080
rect 3660 5040 3666 5052
rect 4614 5040 4620 5092
rect 4672 5080 4678 5092
rect 5169 5083 5227 5089
rect 5169 5080 5181 5083
rect 4672 5052 5181 5080
rect 4672 5040 4678 5052
rect 5169 5049 5181 5052
rect 5215 5049 5227 5083
rect 5169 5043 5227 5049
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 5460 5080 5488 5188
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 9490 5216 9496 5228
rect 8174 5188 9496 5216
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5148 7619 5151
rect 8174 5148 8202 5188
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9674 5216 9680 5228
rect 9635 5188 9680 5216
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 10318 5216 10324 5228
rect 9824 5188 10324 5216
rect 9824 5176 9830 5188
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 8754 5148 8760 5160
rect 7607 5120 8202 5148
rect 8715 5120 8760 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 11383 5157 11411 5256
rect 11793 5253 11805 5256
rect 11839 5253 11851 5287
rect 11793 5247 11851 5253
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12912 5284 12940 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 14185 5355 14243 5361
rect 14185 5352 14197 5355
rect 14047 5324 14197 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 14185 5321 14197 5324
rect 14231 5352 14243 5355
rect 14231 5324 15470 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 12124 5256 12940 5284
rect 13771 5287 13829 5293
rect 12124 5244 12130 5256
rect 13771 5253 13783 5287
rect 13817 5284 13829 5287
rect 15442 5284 15470 5324
rect 15654 5312 15660 5364
rect 15712 5352 15718 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 15712 5324 16497 5352
rect 15712 5312 15718 5324
rect 16485 5321 16497 5324
rect 16531 5352 16543 5355
rect 19981 5355 20039 5361
rect 19981 5352 19993 5355
rect 16531 5324 19993 5352
rect 16531 5321 16543 5324
rect 16485 5315 16543 5321
rect 19981 5321 19993 5324
rect 20027 5352 20039 5355
rect 20806 5352 20812 5364
rect 20027 5324 20812 5352
rect 20027 5321 20039 5324
rect 19981 5315 20039 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 15746 5284 15752 5296
rect 13817 5256 14780 5284
rect 15442 5256 15752 5284
rect 13817 5253 13829 5256
rect 13771 5247 13829 5253
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12703 5188 13185 5216
rect 12703 5157 12731 5188
rect 13173 5185 13185 5188
rect 13219 5216 13231 5219
rect 14366 5216 14372 5228
rect 13219 5188 14372 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 14752 5225 14780 5256
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 16114 5244 16120 5296
rect 16172 5284 16178 5296
rect 17402 5284 17408 5296
rect 16172 5256 17408 5284
rect 16172 5244 16178 5256
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 17494 5244 17500 5296
rect 17552 5284 17558 5296
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 17552 5256 17785 5284
rect 17552 5244 17558 5256
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 17862 5244 17868 5296
rect 17920 5284 17926 5296
rect 18187 5287 18245 5293
rect 18187 5284 18199 5287
rect 17920 5256 18199 5284
rect 17920 5244 17926 5256
rect 18187 5253 18199 5256
rect 18233 5253 18245 5287
rect 18187 5247 18245 5253
rect 18969 5287 19027 5293
rect 18969 5253 18981 5287
rect 19015 5284 19027 5287
rect 19058 5284 19064 5296
rect 19015 5256 19064 5284
rect 19015 5253 19027 5256
rect 18969 5247 19027 5253
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 19794 5244 19800 5296
rect 19852 5284 19858 5296
rect 20257 5287 20315 5293
rect 20257 5284 20269 5287
rect 19852 5256 20269 5284
rect 19852 5244 19858 5256
rect 20257 5253 20269 5256
rect 20303 5253 20315 5287
rect 20257 5247 20315 5253
rect 20622 5244 20628 5296
rect 20680 5284 20686 5296
rect 21315 5287 21373 5293
rect 21315 5284 21327 5287
rect 20680 5256 21327 5284
rect 20680 5244 20686 5256
rect 21315 5253 21327 5256
rect 21361 5253 21373 5287
rect 21315 5247 21373 5253
rect 14737 5219 14795 5225
rect 14737 5185 14749 5219
rect 14783 5216 14795 5219
rect 18322 5216 18328 5228
rect 14783 5188 18328 5216
rect 14783 5185 14795 5188
rect 14737 5179 14795 5185
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 19076 5216 19104 5244
rect 19076 5188 19196 5216
rect 11368 5151 11426 5157
rect 11368 5117 11380 5151
rect 11414 5117 11426 5151
rect 11368 5111 11426 5117
rect 12688 5151 12746 5157
rect 12688 5117 12700 5151
rect 12734 5117 12746 5151
rect 12688 5111 12746 5117
rect 13700 5151 13758 5157
rect 13700 5117 13712 5151
rect 13746 5148 13758 5151
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13746 5120 14013 5148
rect 13746 5117 13758 5120
rect 13700 5111 13758 5117
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14001 5111 14059 5117
rect 15381 5151 15439 5157
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 15427 5120 15485 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 15654 5148 15660 5160
rect 15615 5120 15660 5148
rect 15473 5111 15531 5117
rect 5626 5080 5632 5092
rect 5316 5052 5361 5080
rect 5460 5052 5632 5080
rect 5316 5040 5322 5052
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 5813 5083 5871 5089
rect 5813 5049 5825 5083
rect 5859 5049 5871 5083
rect 5994 5080 6000 5092
rect 5955 5052 6000 5080
rect 5813 5043 5871 5049
rect 845 5015 903 5021
rect 845 4981 857 5015
rect 891 5012 903 5015
rect 1946 5012 1952 5024
rect 891 4984 1952 5012
rect 891 4981 903 4984
rect 845 4975 903 4981
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 2774 5012 2780 5024
rect 2735 4984 2780 5012
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 3329 5015 3387 5021
rect 3329 4981 3341 5015
rect 3375 5012 3387 5015
rect 4338 5012 4344 5024
rect 3375 4984 4344 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 4338 4972 4344 4984
rect 4396 5012 4402 5024
rect 5276 5012 5304 5040
rect 4396 4984 5304 5012
rect 5828 5012 5856 5043
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 6089 5083 6147 5089
rect 6089 5049 6101 5083
rect 6135 5080 6147 5083
rect 6362 5080 6368 5092
rect 6135 5052 6368 5080
rect 6135 5049 6147 5052
rect 6089 5043 6147 5049
rect 6362 5040 6368 5052
rect 6420 5040 6426 5092
rect 6638 5040 6644 5092
rect 6696 5080 6702 5092
rect 6917 5083 6975 5089
rect 6917 5080 6929 5083
rect 6696 5052 6929 5080
rect 6696 5040 6702 5052
rect 6917 5049 6929 5052
rect 6963 5049 6975 5083
rect 6917 5043 6975 5049
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 7064 5052 7109 5080
rect 7064 5040 7070 5052
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 8352 5052 9781 5080
rect 8352 5040 8358 5052
rect 9769 5049 9781 5052
rect 9815 5080 9827 5083
rect 12066 5080 12072 5092
rect 9815 5052 12072 5080
rect 9815 5049 9827 5052
rect 9769 5043 9827 5049
rect 12066 5040 12072 5052
rect 12124 5040 12130 5092
rect 13078 5040 13084 5092
rect 13136 5080 13142 5092
rect 14461 5083 14519 5089
rect 14461 5080 14473 5083
rect 13136 5052 14473 5080
rect 13136 5040 13142 5052
rect 14461 5049 14473 5052
rect 14507 5080 14519 5083
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 14507 5052 14841 5080
rect 14507 5049 14519 5052
rect 14461 5043 14519 5049
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 14829 5043 14887 5049
rect 6730 5012 6736 5024
rect 5828 4984 6736 5012
rect 4396 4972 4402 4984
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 8168 4984 8217 5012
rect 8168 4972 8174 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 8444 4984 9413 5012
rect 8444 4972 8450 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 10686 5012 10692 5024
rect 10599 4984 10692 5012
rect 9401 4975 9459 4981
rect 10686 4972 10692 4984
rect 10744 5012 10750 5024
rect 11057 5015 11115 5021
rect 11057 5012 11069 5015
rect 10744 4984 11069 5012
rect 10744 4972 10750 4984
rect 11057 4981 11069 4984
rect 11103 5012 11115 5015
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11103 4984 12265 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 12253 4981 12265 4984
rect 12299 5012 12311 5015
rect 12618 5012 12624 5024
rect 12299 4984 12624 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 12759 5015 12817 5021
rect 12759 4981 12771 5015
rect 12805 5012 12817 5015
rect 12894 5012 12900 5024
rect 12805 4984 12900 5012
rect 12805 4981 12817 4984
rect 12759 4975 12817 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 14001 5015 14059 5021
rect 14001 5012 14013 5015
rect 13688 4984 14013 5012
rect 13688 4972 13694 4984
rect 14001 4981 14013 4984
rect 14047 4981 14059 5015
rect 14844 5012 14872 5043
rect 15010 5040 15016 5092
rect 15068 5080 15074 5092
rect 15396 5080 15424 5111
rect 15654 5108 15660 5120
rect 15712 5148 15718 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15712 5120 16037 5148
rect 15712 5108 15718 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16025 5111 16083 5117
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 18084 5151 18142 5157
rect 18084 5148 18096 5151
rect 17736 5120 18096 5148
rect 17736 5108 17742 5120
rect 18084 5117 18096 5120
rect 18130 5148 18142 5151
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 18130 5120 18521 5148
rect 18130 5117 18142 5120
rect 18084 5111 18142 5117
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 18966 5108 18972 5160
rect 19024 5148 19030 5160
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 19024 5120 19073 5148
rect 19024 5108 19030 5120
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 16482 5080 16488 5092
rect 15068 5052 15424 5080
rect 15488 5052 16488 5080
rect 15068 5040 15074 5052
rect 15488 5012 15516 5052
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 16991 5083 17049 5089
rect 16991 5049 17003 5083
rect 17037 5080 17049 5083
rect 17494 5080 17500 5092
rect 17037 5052 17500 5080
rect 17037 5049 17049 5052
rect 16991 5043 17049 5049
rect 17494 5040 17500 5052
rect 17552 5040 17558 5092
rect 18325 5083 18383 5089
rect 18325 5049 18337 5083
rect 18371 5080 18383 5083
rect 19168 5080 19196 5188
rect 21244 5151 21302 5157
rect 21244 5117 21256 5151
rect 21290 5148 21302 5151
rect 21637 5151 21695 5157
rect 21637 5148 21649 5151
rect 21290 5120 21649 5148
rect 21290 5117 21302 5120
rect 21244 5111 21302 5117
rect 21637 5117 21649 5120
rect 21683 5148 21695 5151
rect 22738 5148 22744 5160
rect 21683 5120 22744 5148
rect 21683 5117 21695 5120
rect 21637 5111 21695 5117
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 19382 5083 19440 5089
rect 19382 5080 19394 5083
rect 18371 5052 19394 5080
rect 18371 5049 18383 5052
rect 18325 5043 18383 5049
rect 19382 5049 19394 5052
rect 19428 5049 19440 5083
rect 19382 5043 19440 5049
rect 14844 4984 15516 5012
rect 15565 5015 15623 5021
rect 14001 4975 14059 4981
rect 15565 4981 15577 5015
rect 15611 5012 15623 5015
rect 16114 5012 16120 5024
rect 15611 4984 16120 5012
rect 15611 4981 15623 4984
rect 15565 4975 15623 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 16908 4984 17417 5012
rect 16908 4972 16914 4984
rect 17405 4981 17417 4984
rect 17451 5012 17463 5015
rect 17586 5012 17592 5024
rect 17451 4984 17592 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 20438 4972 20444 5024
rect 20496 5012 20502 5024
rect 20901 5015 20959 5021
rect 20901 5012 20913 5015
rect 20496 4984 20913 5012
rect 20496 4972 20502 4984
rect 20901 4981 20913 4984
rect 20947 4981 20959 5015
rect 22002 5012 22008 5024
rect 21963 4984 22008 5012
rect 20901 4975 20959 4981
rect 22002 4972 22008 4984
rect 22060 4972 22066 5024
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 22373 5015 22431 5021
rect 22373 5012 22385 5015
rect 22244 4984 22385 5012
rect 22244 4972 22250 4984
rect 22373 4981 22385 4984
rect 22419 4981 22431 5015
rect 22373 4975 22431 4981
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 1762 4808 1768 4820
rect 1723 4780 1768 4808
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 3418 4808 3424 4820
rect 2363 4780 3424 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 4338 4768 4344 4820
rect 4396 4808 4402 4820
rect 5350 4808 5356 4820
rect 4396 4780 5356 4808
rect 4396 4768 4402 4780
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 5626 4808 5632 4820
rect 5583 4780 5632 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 6420 4780 6776 4808
rect 6420 4768 6426 4780
rect 1780 4740 1808 4768
rect 2774 4749 2780 4752
rect 2730 4743 2780 4749
rect 2730 4740 2742 4743
rect 1780 4712 2742 4740
rect 2730 4709 2742 4712
rect 2776 4709 2780 4743
rect 2730 4703 2780 4709
rect 2774 4700 2780 4703
rect 2832 4700 2838 4752
rect 3640 4743 3698 4749
rect 3640 4709 3652 4743
rect 3686 4740 3698 4743
rect 3878 4740 3884 4752
rect 3686 4712 3884 4740
rect 3686 4709 3698 4712
rect 3640 4703 3698 4709
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4614 4700 4620 4752
rect 4672 4700 4678 4752
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 5905 4743 5963 4749
rect 5905 4740 5917 4743
rect 4856 4712 5917 4740
rect 4856 4700 4862 4712
rect 5905 4709 5917 4712
rect 5951 4740 5963 4743
rect 6638 4740 6644 4752
rect 5951 4712 6500 4740
rect 6599 4712 6644 4740
rect 5951 4709 5963 4712
rect 5905 4703 5963 4709
rect 382 4632 388 4684
rect 440 4672 446 4684
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 440 4644 2421 4672
rect 440 4632 446 4644
rect 2409 4641 2421 4644
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4672 3479 4675
rect 3510 4672 3516 4684
rect 3467 4644 3516 4672
rect 3467 4641 3479 4644
rect 3421 4635 3479 4641
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 3764 4675 3822 4681
rect 3764 4641 3776 4675
rect 3810 4641 3822 4675
rect 3764 4635 3822 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4522 4672 4528 4684
rect 4483 4644 4528 4672
rect 4341 4635 4399 4641
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1486 4604 1492 4616
rect 1443 4576 1492 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1486 4564 1492 4576
rect 1544 4564 1550 4616
rect 3779 4604 3807 4635
rect 3970 4604 3976 4616
rect 3779 4576 3976 4604
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4356 4604 4384 4635
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 4632 4672 4660 4700
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4632 4644 4905 4672
rect 4893 4641 4905 4644
rect 4939 4641 4951 4675
rect 4893 4635 4951 4641
rect 5040 4675 5098 4681
rect 5040 4641 5052 4675
rect 5086 4672 5098 4675
rect 5166 4672 5172 4684
rect 5086 4644 5172 4672
rect 5086 4641 5098 4644
rect 5040 4635 5098 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 5534 4672 5540 4684
rect 5408 4644 5540 4672
rect 5408 4632 5414 4644
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 4430 4604 4436 4616
rect 4356 4576 4436 4604
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4614 4604 4620 4616
rect 4575 4576 4620 4604
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5626 4604 5632 4616
rect 5307 4576 5632 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 5813 4567 5871 4573
rect 3329 4539 3387 4545
rect 3329 4505 3341 4539
rect 3375 4536 3387 4539
rect 3375 4508 4154 4536
rect 3375 4505 3387 4508
rect 3329 4499 3387 4505
rect 477 4471 535 4477
rect 477 4437 489 4471
rect 523 4468 535 4471
rect 3835 4471 3893 4477
rect 3835 4468 3847 4471
rect 523 4440 3847 4468
rect 523 4437 535 4440
rect 477 4431 535 4437
rect 3835 4437 3847 4440
rect 3881 4437 3893 4471
rect 4126 4468 4154 4508
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 5828 4536 5856 4567
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 6472 4604 6500 4712
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 6748 4749 6776 4780
rect 7374 4768 7380 4820
rect 7432 4808 7438 4820
rect 8478 4808 8484 4820
rect 7432 4780 8484 4808
rect 7432 4768 7438 4780
rect 8478 4768 8484 4780
rect 8536 4808 8542 4820
rect 11054 4808 11060 4820
rect 8536 4780 11060 4808
rect 8536 4768 8542 4780
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 14148 4780 14289 4808
rect 14148 4768 14154 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 14277 4771 14335 4777
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 16850 4808 16856 4820
rect 14424 4780 16856 4808
rect 14424 4768 14430 4780
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 17770 4808 17776 4820
rect 17731 4780 17776 4808
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 17920 4780 21925 4808
rect 17920 4768 17926 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 21913 4771 21971 4777
rect 6733 4743 6791 4749
rect 6733 4709 6745 4743
rect 6779 4740 6791 4743
rect 7098 4740 7104 4752
rect 6779 4712 7104 4740
rect 6779 4709 6791 4712
rect 6733 4703 6791 4709
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 7558 4740 7564 4752
rect 7340 4712 7564 4740
rect 7340 4700 7346 4712
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 8110 4740 8116 4752
rect 8071 4712 8116 4740
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 8352 4712 8401 4740
rect 8352 4700 8358 4712
rect 8389 4709 8401 4712
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 7469 4607 7527 4613
rect 6472 4576 6868 4604
rect 6288 4536 6316 4564
rect 4304 4508 5165 4536
rect 4304 4496 4310 4508
rect 4430 4468 4436 4480
rect 4126 4440 4436 4468
rect 3835 4431 3893 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 4522 4428 4528 4480
rect 4580 4468 4586 4480
rect 4706 4468 4712 4480
rect 4580 4440 4712 4468
rect 4580 4428 4586 4440
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 5137 4468 5165 4508
rect 5276 4508 5672 4536
rect 5828 4508 6316 4536
rect 5169 4471 5227 4477
rect 5169 4468 5181 4471
rect 5137 4440 5181 4468
rect 5169 4437 5181 4440
rect 5215 4468 5227 4471
rect 5276 4468 5304 4508
rect 5644 4480 5672 4508
rect 5215 4440 5304 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5626 4428 5632 4480
rect 5684 4428 5690 4480
rect 6840 4468 6868 4576
rect 7469 4573 7481 4607
rect 7515 4604 7527 4607
rect 7650 4604 7656 4616
rect 7515 4576 7656 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 7190 4536 7196 4548
rect 7151 4508 7196 4536
rect 7190 4496 7196 4508
rect 7248 4536 7254 4548
rect 7248 4508 7696 4536
rect 7248 4496 7254 4508
rect 7668 4468 7696 4508
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8312 4536 8340 4567
rect 7800 4508 8340 4536
rect 8496 4536 8524 4768
rect 8662 4700 8668 4752
rect 8720 4740 8726 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 8720 4712 9873 4740
rect 8720 4700 8726 4712
rect 9861 4709 9873 4712
rect 9907 4740 9919 4743
rect 11146 4740 11152 4752
rect 9907 4712 11152 4740
rect 9907 4709 9919 4712
rect 9861 4703 9919 4709
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 11787 4743 11845 4749
rect 11787 4709 11799 4743
rect 11833 4740 11845 4743
rect 12618 4740 12624 4752
rect 11833 4712 12624 4740
rect 11833 4709 11845 4712
rect 11787 4703 11845 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 13262 4740 13268 4752
rect 13223 4712 13268 4740
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 13357 4743 13415 4749
rect 13357 4709 13369 4743
rect 13403 4740 13415 4743
rect 14182 4740 14188 4752
rect 13403 4712 14188 4740
rect 13403 4709 13415 4712
rect 13357 4703 13415 4709
rect 14182 4700 14188 4712
rect 14240 4740 14246 4752
rect 14240 4712 15608 4740
rect 14240 4700 14246 4712
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9490 4672 9496 4684
rect 8987 4644 9496 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 12250 4672 12256 4684
rect 11471 4644 12256 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 13078 4672 13084 4684
rect 12391 4644 13084 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14458 4672 14464 4684
rect 13955 4644 14464 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14458 4632 14464 4644
rect 14516 4672 14522 4684
rect 14516 4644 15470 4672
rect 14516 4632 14522 4644
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 8628 4576 9229 4604
rect 8628 4564 8634 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 9766 4604 9772 4616
rect 9727 4576 9772 4604
rect 9217 4567 9275 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 9916 4576 11161 4604
rect 9916 4564 9922 4576
rect 11149 4573 11161 4576
rect 11195 4604 11207 4607
rect 12802 4604 12808 4616
rect 11195 4576 12808 4604
rect 11195 4573 11207 4576
rect 11149 4567 11207 4573
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 15286 4604 15292 4616
rect 13688 4576 15292 4604
rect 13688 4564 13694 4576
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 8496 4508 8708 4536
rect 7800 4496 7806 4508
rect 8570 4468 8576 4480
rect 6840 4440 8576 4468
rect 7668 4400 7696 4440
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8680 4468 8708 4508
rect 9582 4496 9588 4548
rect 9640 4536 9646 4548
rect 10321 4539 10379 4545
rect 10321 4536 10333 4539
rect 9640 4508 10333 4536
rect 9640 4496 9646 4508
rect 10321 4505 10333 4508
rect 10367 4505 10379 4539
rect 10321 4499 10379 4505
rect 13538 4496 13544 4548
rect 13596 4536 13602 4548
rect 14553 4539 14611 4545
rect 14553 4536 14565 4539
rect 13596 4508 14565 4536
rect 13596 4496 13602 4508
rect 14553 4505 14565 4508
rect 14599 4536 14611 4539
rect 14921 4539 14979 4545
rect 14921 4536 14933 4539
rect 14599 4508 14933 4536
rect 14599 4505 14611 4508
rect 14553 4499 14611 4505
rect 14921 4505 14933 4508
rect 14967 4505 14979 4539
rect 15442 4536 15470 4644
rect 15580 4613 15608 4712
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 16530 4743 16588 4749
rect 16530 4740 16542 4743
rect 16356 4712 16542 4740
rect 16356 4700 16362 4712
rect 16530 4709 16542 4712
rect 16576 4709 16588 4743
rect 19426 4740 19432 4752
rect 16530 4703 16588 4709
rect 18937 4712 19432 4740
rect 16206 4672 16212 4684
rect 16167 4644 16212 4672
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4672 17187 4675
rect 18937 4672 18965 4712
rect 19426 4700 19432 4712
rect 19484 4740 19490 4752
rect 20806 4740 20812 4752
rect 19484 4712 20812 4740
rect 19484 4700 19490 4712
rect 20806 4700 20812 4712
rect 20864 4740 20870 4752
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 20864 4712 21097 4740
rect 20864 4700 20870 4712
rect 21085 4709 21097 4712
rect 21131 4709 21143 4743
rect 21634 4740 21640 4752
rect 21595 4712 21640 4740
rect 21085 4703 21143 4709
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 17175 4644 18965 4672
rect 19751 4675 19809 4681
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 19751 4641 19763 4675
rect 19797 4641 19809 4675
rect 19751 4635 19809 4641
rect 19843 4675 19901 4681
rect 19843 4641 19855 4675
rect 19889 4672 19901 4675
rect 19978 4672 19984 4684
rect 19889 4644 19984 4672
rect 19889 4641 19901 4644
rect 19843 4635 19901 4641
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4604 15623 4607
rect 16025 4607 16083 4613
rect 16025 4604 16037 4607
rect 15611 4576 16037 4604
rect 15611 4573 15623 4576
rect 15565 4567 15623 4573
rect 16025 4573 16037 4576
rect 16071 4573 16083 4607
rect 16224 4604 16252 4632
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 16224 4576 17417 4604
rect 16025 4567 16083 4573
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17586 4564 17592 4616
rect 17644 4604 17650 4616
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17644 4576 17969 4604
rect 17644 4564 17650 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 19058 4564 19064 4616
rect 19116 4604 19122 4616
rect 19153 4607 19211 4613
rect 19153 4604 19165 4607
rect 19116 4576 19165 4604
rect 19116 4564 19122 4576
rect 19153 4573 19165 4576
rect 19199 4573 19211 4607
rect 19766 4604 19794 4635
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 20162 4672 20168 4684
rect 20123 4644 20168 4672
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 20346 4632 20352 4684
rect 20404 4672 20410 4684
rect 20533 4675 20591 4681
rect 20533 4672 20545 4675
rect 20404 4644 20545 4672
rect 20404 4632 20410 4644
rect 20533 4641 20545 4644
rect 20579 4672 20591 4675
rect 20622 4672 20628 4684
rect 20579 4644 20628 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 21729 4675 21787 4681
rect 21729 4641 21741 4675
rect 21775 4672 21787 4675
rect 22281 4675 22339 4681
rect 22281 4672 22293 4675
rect 21775 4644 22293 4672
rect 21775 4641 21787 4644
rect 21729 4635 21787 4641
rect 22281 4641 22293 4644
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 20070 4604 20076 4616
rect 19766 4576 20076 4604
rect 19153 4567 19211 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20990 4604 20996 4616
rect 20903 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4604 21054 4616
rect 21910 4604 21916 4616
rect 21048 4576 21916 4604
rect 21048 4564 21054 4576
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 16206 4536 16212 4548
rect 15442 4508 16212 4536
rect 14921 4499 14979 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 18877 4539 18935 4545
rect 18877 4536 18889 4539
rect 16586 4508 18889 4536
rect 10689 4471 10747 4477
rect 10689 4468 10701 4471
rect 8680 4440 10701 4468
rect 10689 4437 10701 4440
rect 10735 4468 10747 4471
rect 12158 4468 12164 4480
rect 10735 4440 12164 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 12713 4471 12771 4477
rect 12713 4468 12725 4471
rect 12676 4440 12725 4468
rect 12676 4428 12682 4440
rect 12713 4437 12725 4440
rect 12759 4468 12771 4471
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 12759 4440 13093 4468
rect 12759 4437 12771 4440
rect 12713 4431 12771 4437
rect 13081 4437 13093 4440
rect 13127 4468 13139 4471
rect 13354 4468 13360 4480
rect 13127 4440 13360 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14090 4468 14096 4480
rect 13780 4440 14096 4468
rect 13780 4428 13786 4440
rect 14090 4428 14096 4440
rect 14148 4468 14154 4480
rect 14826 4468 14832 4480
rect 14148 4440 14832 4468
rect 14148 4428 14154 4440
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15562 4428 15568 4480
rect 15620 4468 15626 4480
rect 15841 4471 15899 4477
rect 15841 4468 15853 4471
rect 15620 4440 15853 4468
rect 15620 4428 15626 4440
rect 15841 4437 15853 4440
rect 15887 4437 15899 4471
rect 15841 4431 15899 4437
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4468 16083 4471
rect 16586 4468 16614 4508
rect 18877 4505 18889 4508
rect 18923 4505 18935 4539
rect 18877 4499 18935 4505
rect 18966 4496 18972 4548
rect 19024 4536 19030 4548
rect 19521 4539 19579 4545
rect 19521 4536 19533 4539
rect 19024 4508 19533 4536
rect 19024 4496 19030 4508
rect 19521 4505 19533 4508
rect 19567 4505 19579 4539
rect 19521 4499 19579 4505
rect 16071 4440 16614 4468
rect 16071 4437 16083 4440
rect 16025 4431 16083 4437
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 18138 4468 18144 4480
rect 17736 4440 18144 4468
rect 17736 4428 17742 4440
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 21729 4471 21787 4477
rect 21729 4468 21741 4471
rect 19668 4440 21741 4468
rect 19668 4428 19674 4440
rect 21729 4437 21741 4440
rect 21775 4437 21787 4471
rect 21729 4431 21787 4437
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 2409 4267 2467 4273
rect 2409 4233 2421 4267
rect 2455 4264 2467 4267
rect 4893 4267 4951 4273
rect 2455 4236 4660 4264
rect 2455 4233 2467 4236
rect 2409 4227 2467 4233
rect 2682 4196 2688 4208
rect 2643 4168 2688 4196
rect 2682 4156 2688 4168
rect 2740 4156 2746 4208
rect 4338 4156 4344 4208
rect 4396 4205 4402 4208
rect 4396 4199 4445 4205
rect 4396 4165 4399 4199
rect 4433 4165 4445 4199
rect 4396 4159 4445 4165
rect 4396 4156 4402 4159
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 3050 4128 3056 4140
rect 1535 4100 3056 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 4632 4128 4660 4236
rect 4893 4233 4905 4267
rect 4939 4264 4951 4267
rect 6089 4267 6147 4273
rect 6089 4264 6101 4267
rect 4939 4236 6101 4264
rect 4939 4233 4951 4236
rect 4893 4227 4951 4233
rect 6089 4233 6101 4236
rect 6135 4233 6147 4267
rect 6089 4227 6147 4233
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7668 4264 7696 4304
rect 7156 4236 8064 4264
rect 7156 4224 7162 4236
rect 4709 4199 4767 4205
rect 4709 4165 4721 4199
rect 4755 4196 4767 4199
rect 7374 4196 7380 4208
rect 4755 4168 7380 4196
rect 4755 4165 4767 4168
rect 4709 4159 4767 4165
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 7668 4196 7696 4236
rect 8036 4196 8064 4236
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8168 4236 8340 4264
rect 8168 4224 8174 4236
rect 8312 4205 8340 4236
rect 9306 4224 9312 4276
rect 9364 4224 9370 4276
rect 11471 4267 11529 4273
rect 9646 4236 10916 4264
rect 8297 4199 8355 4205
rect 8297 4196 8309 4199
rect 7668 4168 7788 4196
rect 8036 4168 8309 4196
rect 7760 4137 7788 4168
rect 8297 4165 8309 4168
rect 8343 4196 8355 4199
rect 8846 4196 8852 4208
rect 8343 4168 8852 4196
rect 8343 4165 8355 4168
rect 8297 4159 8355 4165
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 7745 4131 7803 4137
rect 4632 4100 7604 4128
rect 7576 4072 7604 4100
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9324 4128 9352 4224
rect 9646 4208 9674 4236
rect 9582 4156 9588 4208
rect 9640 4168 9674 4208
rect 9640 4156 9646 4168
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9263 4100 10057 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10226 4128 10232 4140
rect 10187 4100 10232 4128
rect 10045 4091 10103 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 2498 4060 2504 4072
rect 2459 4032 2504 4060
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 3237 4063 3295 4069
rect 2915 4032 3188 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 3160 3992 3188 4032
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3326 4060 3332 4072
rect 3283 4032 3332 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 4284 4063 4342 4069
rect 4284 4060 4296 4063
rect 3936 4032 4296 4060
rect 3936 4020 3942 4032
rect 4284 4029 4296 4032
rect 4330 4029 4342 4063
rect 4522 4060 4528 4072
rect 4483 4032 4528 4060
rect 4284 4023 4342 4029
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4060 5043 4063
rect 5902 4060 5908 4072
rect 5031 4032 5908 4060
rect 5031 4029 5043 4032
rect 4985 4023 5043 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6064 4063 6122 4069
rect 6064 4029 6076 4063
rect 6110 4060 6122 4063
rect 6178 4060 6184 4072
rect 6110 4032 6184 4060
rect 6110 4029 6122 4032
rect 6064 4023 6122 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6324 4063 6382 4069
rect 6324 4029 6336 4063
rect 6370 4060 6382 4063
rect 6546 4060 6552 4072
rect 6370 4032 6552 4060
rect 6370 4029 6382 4032
rect 6324 4023 6382 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6822 4060 6828 4072
rect 6783 4032 6828 4060
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7248 4032 7297 4060
rect 7248 4020 7254 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7558 4020 7564 4072
rect 7616 4020 7622 4072
rect 3559 3995 3617 4001
rect 3160 3964 3280 3992
rect 3252 3936 3280 3964
rect 3559 3961 3571 3995
rect 3605 3961 3617 3995
rect 3559 3955 3617 3961
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1820 3896 1869 3924
rect 1820 3884 1826 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 3234 3884 3240 3936
rect 3292 3884 3298 3936
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3574 3924 3602 3955
rect 3694 3952 3700 4004
rect 3752 3992 3758 4004
rect 4893 3995 4951 4001
rect 4893 3992 4905 3995
rect 3752 3964 4905 3992
rect 3752 3952 3758 3964
rect 4893 3961 4905 3964
rect 4939 3961 4951 3995
rect 4893 3955 4951 3961
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7837 3995 7895 4001
rect 7837 3992 7849 3995
rect 6788 3964 7849 3992
rect 6788 3952 6794 3964
rect 7837 3961 7849 3964
rect 7883 3961 7895 3995
rect 7837 3955 7895 3961
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 8573 3995 8631 4001
rect 8573 3992 8585 3995
rect 8168 3964 8585 3992
rect 8168 3952 8174 3964
rect 8573 3961 8585 3964
rect 8619 3961 8631 3995
rect 8573 3955 8631 3961
rect 8662 3952 8668 4004
rect 8720 3992 8726 4004
rect 8720 3964 8765 3992
rect 8720 3952 8726 3964
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9401 3995 9459 4001
rect 9401 3992 9413 3995
rect 9272 3964 9413 3992
rect 9272 3952 9278 3964
rect 9401 3961 9413 3964
rect 9447 3961 9459 3995
rect 9401 3955 9459 3961
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3961 9551 3995
rect 9493 3955 9551 3961
rect 3384 3896 3602 3924
rect 4157 3927 4215 3933
rect 3384 3884 3390 3896
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4798 3924 4804 3936
rect 4203 3896 4804 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 5316 3896 5365 3924
rect 5316 3884 5322 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5353 3887 5411 3893
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 6411 3927 6469 3933
rect 6411 3893 6423 3927
rect 6457 3924 6469 3927
rect 6638 3924 6644 3936
rect 6457 3896 6644 3924
rect 6457 3893 6469 3896
rect 6411 3887 6469 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 6917 3927 6975 3933
rect 6917 3924 6929 3927
rect 6880 3896 6929 3924
rect 6880 3884 6886 3896
rect 6917 3893 6929 3896
rect 6963 3893 6975 3927
rect 6917 3887 6975 3893
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 7742 3924 7748 3936
rect 7248 3896 7748 3924
rect 7248 3884 7254 3896
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9508 3924 9536 3955
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 10888 4001 10916 4236
rect 11471 4233 11483 4267
rect 11517 4264 11529 4267
rect 13630 4264 13636 4276
rect 11517 4236 13636 4264
rect 11517 4233 11529 4236
rect 11471 4227 11529 4233
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 13906 4224 13912 4276
rect 13964 4264 13970 4276
rect 14642 4264 14648 4276
rect 13964 4236 14648 4264
rect 13964 4224 13970 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 15243 4267 15301 4273
rect 15243 4264 15255 4267
rect 15160 4236 15255 4264
rect 15160 4224 15166 4236
rect 15243 4233 15255 4236
rect 15289 4233 15301 4267
rect 15243 4227 15301 4233
rect 16025 4267 16083 4273
rect 16025 4233 16037 4267
rect 16071 4264 16083 4267
rect 16298 4264 16304 4276
rect 16071 4236 16304 4264
rect 16071 4233 16083 4236
rect 16025 4227 16083 4233
rect 11790 4196 11796 4208
rect 11751 4168 11796 4196
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12575 4199 12633 4205
rect 12575 4165 12587 4199
rect 12621 4196 12633 4199
rect 13262 4196 13268 4208
rect 12621 4168 13268 4196
rect 12621 4165 12633 4168
rect 12575 4159 12633 4165
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 14826 4196 14832 4208
rect 14787 4168 14832 4196
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 16040 4196 16068 4227
rect 16298 4224 16304 4236
rect 16356 4264 16362 4276
rect 16850 4264 16856 4276
rect 16356 4236 16856 4264
rect 16356 4224 16362 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 19058 4264 19064 4276
rect 17911 4236 19064 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 19518 4224 19524 4276
rect 19576 4264 19582 4276
rect 19576 4236 20024 4264
rect 19576 4224 19582 4236
rect 19245 4199 19303 4205
rect 19245 4196 19257 4199
rect 15371 4168 16068 4196
rect 17880 4168 18920 4196
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11974 4128 11980 4140
rect 11204 4100 11980 4128
rect 11204 4088 11210 4100
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 13354 4128 13360 4140
rect 13267 4100 13360 4128
rect 13354 4088 13360 4100
rect 13412 4128 13418 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 13412 4100 14565 4128
rect 13412 4088 13418 4100
rect 14553 4097 14565 4100
rect 14599 4128 14611 4131
rect 14734 4128 14740 4140
rect 14599 4100 14740 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 14734 4088 14740 4100
rect 14792 4128 14798 4140
rect 15371 4128 15399 4168
rect 14792 4100 15399 4128
rect 14792 4088 14798 4100
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 17402 4128 17408 4140
rect 16264 4100 16896 4128
rect 17363 4100 17408 4128
rect 16264 4088 16270 4100
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11368 4063 11426 4069
rect 11368 4060 11380 4063
rect 11296 4032 11380 4060
rect 11296 4020 11302 4032
rect 11368 4029 11380 4032
rect 11414 4029 11426 4063
rect 11368 4023 11426 4029
rect 10873 3995 10931 4001
rect 10376 3964 10469 3992
rect 10376 3952 10382 3964
rect 10873 3961 10885 3995
rect 10919 3992 10931 3995
rect 10919 3964 11284 3992
rect 10919 3961 10931 3964
rect 10873 3955 10931 3961
rect 10336 3924 10364 3952
rect 11256 3936 11284 3964
rect 8352 3896 10364 3924
rect 8352 3884 8358 3896
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11112 3896 11161 3924
rect 11112 3884 11118 3896
rect 11149 3893 11161 3896
rect 11195 3893 11207 3927
rect 11149 3887 11207 3893
rect 11238 3884 11244 3936
rect 11296 3884 11302 3936
rect 11383 3924 11411 4023
rect 11606 4020 11612 4072
rect 11664 4060 11670 4072
rect 12250 4060 12256 4072
rect 11664 4032 12256 4060
rect 11664 4020 11670 4032
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12504 4063 12562 4069
rect 12504 4029 12516 4063
rect 12550 4060 12562 4063
rect 12710 4060 12716 4072
rect 12550 4032 12716 4060
rect 12550 4029 12562 4032
rect 12504 4023 12562 4029
rect 12710 4020 12716 4032
rect 12768 4060 12774 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12768 4032 12909 4060
rect 12768 4020 12774 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 16868 4069 16896 4100
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 15140 4063 15198 4069
rect 15140 4060 15152 4063
rect 14332 4032 15152 4060
rect 14332 4020 14338 4032
rect 15140 4029 15152 4032
rect 15186 4060 15198 4063
rect 15565 4063 15623 4069
rect 15565 4060 15577 4063
rect 15186 4032 15577 4060
rect 15186 4029 15198 4032
rect 15140 4023 15198 4029
rect 15565 4029 15577 4032
rect 15611 4029 15623 4063
rect 15565 4023 15623 4029
rect 16853 4063 16911 4069
rect 16853 4029 16865 4063
rect 16899 4060 16911 4063
rect 17880 4060 17908 4168
rect 18414 4128 18420 4140
rect 18375 4100 18420 4128
rect 18414 4088 18420 4100
rect 18472 4128 18478 4140
rect 18782 4128 18788 4140
rect 18472 4100 18788 4128
rect 18472 4088 18478 4100
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 16899 4032 17908 4060
rect 16899 4029 16911 4032
rect 16853 4023 16911 4029
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3961 13599 3995
rect 13541 3955 13599 3961
rect 12250 3924 12256 3936
rect 11383 3896 12256 3924
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 13556 3924 13584 3955
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 14185 3995 14243 4001
rect 13688 3964 13733 3992
rect 13688 3952 13694 3964
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 15010 3992 15016 4004
rect 14231 3964 15016 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 16209 3995 16267 4001
rect 16209 3992 16221 3995
rect 15344 3964 16221 3992
rect 15344 3952 15350 3964
rect 16209 3961 16221 3964
rect 16255 3961 16267 3995
rect 16209 3955 16267 3961
rect 14366 3924 14372 3936
rect 13556 3896 14372 3924
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 16224 3924 16252 3955
rect 16298 3952 16304 4004
rect 16356 3992 16362 4004
rect 17954 3992 17960 4004
rect 16356 3964 16401 3992
rect 16408 3964 17960 3992
rect 16356 3952 16362 3964
rect 16408 3924 16436 3964
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 18138 3992 18144 4004
rect 18099 3964 18144 3992
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18288 3964 18333 3992
rect 18288 3952 18294 3964
rect 18782 3952 18788 4004
rect 18840 3992 18846 4004
rect 18892 3992 18920 4168
rect 18984 4168 19257 4196
rect 18984 4072 19012 4168
rect 19245 4165 19257 4168
rect 19291 4165 19303 4199
rect 19794 4196 19800 4208
rect 19245 4159 19303 4165
rect 19397 4168 19800 4196
rect 19397 4154 19425 4168
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 19352 4128 19425 4154
rect 19996 4137 20024 4236
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 21634 4224 21640 4276
rect 21692 4264 21698 4276
rect 21910 4264 21916 4276
rect 21692 4236 21916 4264
rect 21692 4224 21698 4236
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 22428 4236 22473 4264
rect 22428 4224 22434 4236
rect 19076 4126 19425 4128
rect 19981 4131 20039 4137
rect 19076 4100 19380 4126
rect 18966 4020 18972 4072
rect 19024 4020 19030 4072
rect 18840 3964 18920 3992
rect 18840 3952 18846 3964
rect 16224 3896 16436 3924
rect 16482 3884 16488 3936
rect 16540 3924 16546 3936
rect 19076 3933 19104 4100
rect 19981 4097 19993 4131
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 21212 4063 21270 4069
rect 21212 4060 21224 4063
rect 20404 4032 21224 4060
rect 20404 4020 20410 4032
rect 21212 4029 21224 4032
rect 21258 4060 21270 4063
rect 21637 4063 21695 4069
rect 21637 4060 21649 4063
rect 21258 4032 21649 4060
rect 21258 4029 21270 4032
rect 21212 4023 21270 4029
rect 21637 4029 21649 4032
rect 21683 4029 21695 4063
rect 21637 4023 21695 4029
rect 19245 3995 19303 4001
rect 19245 3961 19257 3995
rect 19291 3992 19303 3995
rect 19705 3995 19763 4001
rect 19705 3992 19717 3995
rect 19291 3964 19717 3992
rect 19291 3961 19303 3964
rect 19245 3955 19303 3961
rect 19705 3961 19717 3964
rect 19751 3961 19763 3995
rect 19705 3955 19763 3961
rect 19061 3927 19119 3933
rect 19061 3924 19073 3927
rect 16540 3896 19073 3924
rect 16540 3884 16546 3896
rect 19061 3893 19073 3896
rect 19107 3893 19119 3927
rect 19518 3924 19524 3936
rect 19479 3896 19524 3924
rect 19061 3887 19119 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 19720 3924 19748 3955
rect 19794 3952 19800 4004
rect 19852 3992 19858 4004
rect 19852 3964 19897 3992
rect 19852 3952 19858 3964
rect 19668 3896 19748 3924
rect 19668 3884 19674 3896
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 21315 3927 21373 3933
rect 21315 3924 21327 3927
rect 19944 3896 21327 3924
rect 19944 3884 19950 3896
rect 21315 3893 21327 3896
rect 21361 3893 21373 3927
rect 21315 3887 21373 3893
rect 21726 3884 21732 3936
rect 21784 3924 21790 3936
rect 22005 3927 22063 3933
rect 22005 3924 22017 3927
rect 21784 3896 22017 3924
rect 21784 3884 21790 3896
rect 22005 3893 22017 3896
rect 22051 3893 22063 3927
rect 22005 3887 22063 3893
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 1762 3720 1768 3732
rect 1723 3692 1768 3720
rect 1762 3680 1768 3692
rect 1820 3720 1826 3732
rect 3234 3720 3240 3732
rect 1820 3692 3240 3720
rect 1820 3680 1826 3692
rect 2745 3661 2773 3692
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4522 3720 4528 3732
rect 4483 3692 4528 3720
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5077 3723 5135 3729
rect 5077 3689 5089 3723
rect 5123 3720 5135 3723
rect 5350 3720 5356 3732
rect 5123 3692 5356 3720
rect 5123 3689 5135 3692
rect 5077 3683 5135 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 6089 3723 6147 3729
rect 6089 3689 6101 3723
rect 6135 3720 6147 3723
rect 7006 3720 7012 3732
rect 6135 3692 7012 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 8294 3720 8300 3732
rect 8251 3692 8300 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10183 3723 10241 3729
rect 10183 3720 10195 3723
rect 10008 3692 10195 3720
rect 10008 3680 10014 3692
rect 10183 3689 10195 3692
rect 10229 3689 10241 3723
rect 10183 3683 10241 3689
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 10744 3692 10793 3720
rect 10744 3680 10750 3692
rect 10781 3689 10793 3692
rect 10827 3689 10839 3723
rect 10781 3683 10839 3689
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 11379 3692 12801 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 2730 3655 2788 3661
rect 2730 3621 2742 3655
rect 2776 3621 2788 3655
rect 2730 3615 2788 3621
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 4540 3652 4568 3680
rect 5258 3652 5264 3664
rect 2924 3624 4430 3652
rect 4540 3624 5264 3652
rect 2924 3612 2930 3624
rect 1026 3544 1032 3596
rect 1084 3584 1090 3596
rect 1397 3587 1455 3593
rect 1397 3584 1409 3587
rect 1084 3556 1409 3584
rect 1084 3544 1090 3556
rect 1397 3553 1409 3556
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 2004 3556 3341 3584
rect 2004 3544 2010 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3329 3547 3387 3553
rect 3764 3587 3822 3593
rect 3764 3553 3776 3587
rect 3810 3584 3822 3587
rect 4062 3584 4068 3596
rect 3810 3556 4068 3584
rect 3810 3553 3822 3556
rect 3764 3547 3822 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 2682 3516 2688 3528
rect 2455 3488 2688 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 4065 3451 4123 3457
rect 4065 3417 4077 3451
rect 4111 3448 4123 3451
rect 4154 3448 4160 3460
rect 4111 3420 4160 3448
rect 4111 3417 4123 3420
rect 4065 3411 4123 3417
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4402 3448 4430 3624
rect 5258 3612 5264 3624
rect 5316 3652 5322 3664
rect 5490 3655 5548 3661
rect 5490 3652 5502 3655
rect 5316 3624 5502 3652
rect 5316 3612 5322 3624
rect 5490 3621 5502 3624
rect 5536 3621 5548 3655
rect 6362 3652 6368 3664
rect 6323 3624 6368 3652
rect 5490 3615 5548 3621
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 7647 3655 7705 3661
rect 7647 3621 7659 3655
rect 7693 3652 7705 3655
rect 7742 3652 7748 3664
rect 7693 3624 7748 3652
rect 7693 3621 7705 3624
rect 7647 3615 7705 3621
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 7926 3612 7932 3664
rect 7984 3652 7990 3664
rect 8389 3655 8447 3661
rect 8389 3652 8401 3655
rect 7984 3624 8401 3652
rect 7984 3612 7990 3624
rect 8389 3621 8401 3624
rect 8435 3621 8447 3655
rect 8389 3615 8447 3621
rect 8490 3655 8548 3661
rect 8490 3621 8502 3655
rect 8536 3652 8548 3655
rect 9030 3652 9036 3664
rect 8536 3624 9036 3652
rect 8536 3621 8548 3624
rect 8490 3615 8548 3621
rect 9030 3612 9036 3624
rect 9088 3612 9094 3664
rect 9263 3655 9321 3661
rect 9263 3652 9275 3655
rect 9173 3624 9275 3652
rect 9263 3621 9275 3624
rect 9309 3652 9321 3655
rect 9858 3652 9864 3664
rect 9309 3624 9864 3652
rect 9309 3621 9321 3624
rect 9263 3615 9321 3621
rect 9858 3612 9864 3624
rect 9916 3652 9922 3664
rect 9916 3624 10272 3652
rect 9916 3612 9922 3624
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5810 3584 5816 3596
rect 5215 3556 5816 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 9122 3584 9128 3596
rect 6963 3556 7649 3584
rect 9083 3556 9128 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 5776 3488 6285 3516
rect 5776 3476 5782 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 7006 3516 7012 3528
rect 6967 3488 7012 3516
rect 6273 3479 6331 3485
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 7466 3516 7472 3528
rect 7331 3488 7472 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7621 3516 7649 3556
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9674 3584 9680 3596
rect 9732 3593 9738 3596
rect 9732 3587 9770 3593
rect 9548 3556 9680 3584
rect 9548 3544 9554 3556
rect 9674 3544 9680 3556
rect 9758 3584 9770 3587
rect 10080 3587 10138 3593
rect 10080 3584 10092 3587
rect 9758 3556 10092 3584
rect 9758 3553 9770 3556
rect 9732 3547 9770 3553
rect 10080 3553 10092 3556
rect 10126 3553 10138 3587
rect 10244 3584 10272 3624
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 12299 3655 12357 3661
rect 12299 3652 12311 3655
rect 11756 3624 12311 3652
rect 11756 3612 11762 3624
rect 12299 3621 12311 3624
rect 12345 3621 12357 3655
rect 12773 3652 12801 3692
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12952 3692 13001 3720
rect 12952 3680 12958 3692
rect 12989 3689 13001 3692
rect 13035 3720 13047 3723
rect 13262 3720 13268 3732
rect 13035 3692 13268 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13630 3720 13636 3732
rect 13407 3692 13636 3720
rect 13407 3652 13435 3692
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 14461 3723 14519 3729
rect 14461 3689 14473 3723
rect 14507 3720 14519 3723
rect 14734 3720 14740 3732
rect 14507 3692 14740 3720
rect 14507 3689 14519 3692
rect 14461 3683 14519 3689
rect 12773 3624 13435 3652
rect 13535 3655 13593 3661
rect 12299 3615 12357 3621
rect 13535 3621 13547 3655
rect 13581 3652 13593 3655
rect 14476 3652 14504 3683
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 15470 3720 15476 3732
rect 15431 3692 15476 3720
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15979 3723 16037 3729
rect 15979 3689 15991 3723
rect 16025 3720 16037 3723
rect 16114 3720 16120 3732
rect 16025 3692 16120 3720
rect 16025 3689 16037 3692
rect 15979 3683 16037 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 17402 3720 17408 3732
rect 16776 3692 17408 3720
rect 13581 3624 14504 3652
rect 13581 3621 13593 3624
rect 13535 3615 13593 3621
rect 15746 3612 15752 3664
rect 15804 3652 15810 3664
rect 16393 3655 16451 3661
rect 16393 3652 16405 3655
rect 15804 3624 16405 3652
rect 15804 3612 15810 3624
rect 16393 3621 16405 3624
rect 16439 3621 16451 3655
rect 16393 3615 16451 3621
rect 16485 3655 16543 3661
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 16776 3652 16804 3692
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 17773 3723 17831 3729
rect 17773 3689 17785 3723
rect 17819 3689 17831 3723
rect 17773 3683 17831 3689
rect 17865 3723 17923 3729
rect 17865 3689 17877 3723
rect 17911 3720 17923 3723
rect 18046 3720 18052 3732
rect 17911 3692 18052 3720
rect 17911 3689 17923 3692
rect 17865 3683 17923 3689
rect 16531 3624 16804 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 16850 3612 16856 3664
rect 16908 3652 16914 3664
rect 17174 3655 17232 3661
rect 17174 3652 17186 3655
rect 16908 3624 17186 3652
rect 16908 3612 16914 3624
rect 17174 3621 17186 3624
rect 17220 3621 17232 3655
rect 17788 3652 17816 3683
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 19150 3720 19156 3732
rect 19111 3692 19156 3720
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 19702 3720 19708 3732
rect 19663 3692 19708 3720
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 20530 3720 20536 3732
rect 20491 3692 20536 3720
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 21913 3723 21971 3729
rect 21913 3720 21925 3723
rect 20680 3692 21925 3720
rect 20680 3680 20686 3692
rect 21913 3689 21925 3692
rect 21959 3689 21971 3723
rect 21913 3683 21971 3689
rect 18230 3652 18236 3664
rect 17788 3624 18236 3652
rect 17174 3615 17232 3621
rect 18230 3612 18236 3624
rect 18288 3652 18294 3664
rect 18509 3655 18567 3661
rect 18509 3652 18521 3655
rect 18288 3624 18521 3652
rect 18288 3612 18294 3624
rect 18509 3621 18521 3624
rect 18555 3652 18567 3655
rect 20438 3652 20444 3664
rect 18555 3624 20444 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 20438 3612 20444 3624
rect 20496 3612 20502 3664
rect 20806 3612 20812 3664
rect 20864 3652 20870 3664
rect 21085 3655 21143 3661
rect 21085 3652 21097 3655
rect 20864 3624 21097 3652
rect 20864 3612 20870 3624
rect 21085 3621 21097 3624
rect 21131 3621 21143 3655
rect 21085 3615 21143 3621
rect 10244 3556 10640 3584
rect 10080 3547 10138 3553
rect 9732 3544 9738 3547
rect 10226 3516 10232 3528
rect 7621 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10409 3519 10467 3525
rect 10409 3516 10421 3519
rect 10382 3485 10421 3516
rect 10455 3485 10467 3519
rect 10612 3516 10640 3556
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11146 3584 11152 3596
rect 10744 3556 11152 3584
rect 10744 3544 10750 3556
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 12212 3587 12270 3593
rect 12212 3553 12224 3587
rect 12258 3584 12270 3587
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12258 3556 12725 3584
rect 12258 3553 12270 3556
rect 12212 3547 12270 3553
rect 12713 3553 12725 3556
rect 12759 3584 12771 3587
rect 13906 3584 13912 3596
rect 12759 3556 13912 3584
rect 12759 3553 12771 3556
rect 12713 3547 12771 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14093 3587 14151 3593
rect 14093 3553 14105 3587
rect 14139 3584 14151 3587
rect 15562 3584 15568 3596
rect 14139 3556 15568 3584
rect 14139 3553 14151 3556
rect 14093 3547 14151 3553
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 15908 3587 15966 3593
rect 15908 3553 15920 3587
rect 15954 3584 15966 3587
rect 16114 3584 16120 3596
rect 15954 3556 16120 3584
rect 15954 3553 15966 3556
rect 15908 3547 15966 3553
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16206 3544 16212 3596
rect 16264 3584 16270 3596
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 16264 3556 16681 3584
rect 16264 3544 16270 3556
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 18322 3584 18328 3596
rect 18104 3556 18328 3584
rect 18104 3544 18110 3556
rect 18322 3544 18328 3556
rect 18380 3584 18386 3596
rect 18601 3587 18659 3593
rect 18601 3584 18613 3587
rect 18380 3556 18613 3584
rect 18380 3544 18386 3556
rect 18601 3553 18613 3556
rect 18647 3553 18659 3587
rect 18601 3547 18659 3553
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 20257 3587 20315 3593
rect 20257 3584 20269 3587
rect 18748 3556 20269 3584
rect 18748 3544 18754 3556
rect 20257 3553 20269 3556
rect 20303 3553 20315 3587
rect 20257 3547 20315 3553
rect 10778 3516 10784 3528
rect 10612 3488 10784 3516
rect 10382 3479 10467 3485
rect 6730 3448 6736 3460
rect 4402 3420 6736 3448
rect 6730 3408 6736 3420
rect 6788 3408 6794 3460
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 7708 3420 8953 3448
rect 7708 3408 7714 3420
rect 8941 3417 8953 3420
rect 8987 3448 8999 3451
rect 9582 3448 9588 3460
rect 8987 3420 9588 3448
rect 8987 3417 8999 3420
rect 8941 3411 8999 3417
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 10382 3448 10410 3479
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 13780 3488 16497 3516
rect 13780 3476 13786 3488
rect 16485 3485 16497 3488
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16632 3488 16865 3516
rect 16632 3476 16638 3488
rect 16853 3485 16865 3488
rect 16899 3516 16911 3519
rect 19426 3516 19432 3528
rect 16899 3488 19432 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 20772 3488 21005 3516
rect 20772 3476 20778 3488
rect 20993 3485 21005 3488
rect 21039 3516 21051 3519
rect 21174 3516 21180 3528
rect 21039 3488 21180 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3516 21327 3519
rect 21910 3516 21916 3528
rect 21315 3488 21916 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 10962 3448 10968 3460
rect 10382 3420 10968 3448
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 11112 3420 11989 3448
rect 11112 3408 11118 3420
rect 11977 3417 11989 3420
rect 12023 3417 12035 3451
rect 11977 3411 12035 3417
rect 2314 3380 2320 3392
rect 2275 3352 2320 3380
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 3835 3383 3893 3389
rect 3835 3349 3847 3383
rect 3881 3380 3893 3383
rect 8754 3380 8760 3392
rect 3881 3352 8760 3380
rect 3881 3349 3893 3352
rect 3835 3343 3893 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9815 3383 9873 3389
rect 9815 3349 9827 3383
rect 9861 3380 9873 3383
rect 11422 3380 11428 3392
rect 9861 3352 11428 3380
rect 9861 3349 9873 3352
rect 9815 3343 9873 3349
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 11698 3380 11704 3392
rect 11659 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 13188 3380 13216 3476
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 18785 3451 18843 3457
rect 18785 3448 18797 3451
rect 13688 3420 18797 3448
rect 13688 3408 13694 3420
rect 18785 3417 18797 3420
rect 18831 3417 18843 3451
rect 21284 3448 21312 3479
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 18785 3411 18843 3417
rect 19352 3420 21312 3448
rect 14274 3380 14280 3392
rect 13188 3352 14280 3380
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 15804 3352 17877 3380
rect 15804 3340 15810 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 17865 3343 17923 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 19352 3380 19380 3420
rect 19518 3380 19524 3392
rect 18196 3352 19380 3380
rect 19479 3352 19524 3380
rect 18196 3340 18202 3352
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 22278 3380 22284 3392
rect 22239 3352 22284 3380
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 937 3179 995 3185
rect 937 3145 949 3179
rect 983 3176 995 3179
rect 4341 3179 4399 3185
rect 983 3148 4154 3176
rect 983 3145 995 3148
rect 937 3139 995 3145
rect 1118 3068 1124 3120
rect 1176 3108 1182 3120
rect 4126 3108 4154 3148
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 7282 3176 7288 3188
rect 4387 3148 7288 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 8202 3176 8208 3188
rect 7616 3148 8208 3176
rect 7616 3136 7622 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10686 3176 10692 3188
rect 9548 3148 10692 3176
rect 9548 3136 9554 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 11931 3179 11989 3185
rect 11931 3176 11943 3179
rect 10933 3148 11943 3176
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 1176 3080 3464 3108
rect 4126 3080 6377 3108
rect 1176 3068 1182 3080
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 3436 3049 3464 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6365 3071 6423 3077
rect 6546 3068 6552 3120
rect 6604 3108 6610 3120
rect 8220 3108 8248 3136
rect 9766 3108 9772 3120
rect 6604 3080 7281 3108
rect 8220 3080 9772 3108
rect 6604 3068 6610 3080
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 7098 3040 7104 3052
rect 4479 3012 7104 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7253 3040 7281 3080
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 9950 3108 9956 3120
rect 9911 3080 9956 3108
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 10933 3108 10961 3148
rect 11931 3145 11943 3148
rect 11977 3145 11989 3179
rect 11931 3139 11989 3145
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12207 3179 12265 3185
rect 12207 3176 12219 3179
rect 12124 3148 12219 3176
rect 12124 3136 12130 3148
rect 12207 3145 12219 3148
rect 12253 3145 12265 3179
rect 12207 3139 12265 3145
rect 12575 3179 12633 3185
rect 12575 3145 12587 3179
rect 12621 3176 12633 3179
rect 12621 3148 13814 3176
rect 12621 3145 12633 3148
rect 12575 3139 12633 3145
rect 11790 3108 11796 3120
rect 10100 3080 10961 3108
rect 11716 3080 11796 3108
rect 10100 3068 10106 3080
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7253 3012 7757 3040
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 8386 3040 8392 3052
rect 8347 3012 8392 3040
rect 7745 3003 7803 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 8570 3040 8576 3052
rect 8531 3012 8576 3040
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3040 9275 3043
rect 9398 3040 9404 3052
rect 9263 3012 9404 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 10410 3040 10416 3052
rect 10275 3012 10416 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3040 11115 3043
rect 11330 3040 11336 3052
rect 11103 3012 11336 3040
rect 11103 3009 11115 3012
rect 11057 3003 11115 3009
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 2406 2972 2412 2984
rect 2367 2944 2412 2972
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 5445 2975 5503 2981
rect 2556 2944 4911 2972
rect 2556 2932 2562 2944
rect 3742 2907 3800 2913
rect 3742 2904 3754 2907
rect 2792 2876 3754 2904
rect 2792 2848 2820 2876
rect 3742 2873 3754 2876
rect 3788 2904 3800 2907
rect 3970 2904 3976 2916
rect 3788 2876 3976 2904
rect 3788 2873 3800 2876
rect 3742 2867 3800 2873
rect 3970 2864 3976 2876
rect 4028 2904 4034 2916
rect 4522 2904 4528 2916
rect 4028 2876 4528 2904
rect 4028 2864 4034 2876
rect 4522 2864 4528 2876
rect 4580 2904 4586 2916
rect 4754 2907 4812 2913
rect 4754 2904 4766 2907
rect 4580 2876 4766 2904
rect 4580 2864 4586 2876
rect 4754 2873 4766 2876
rect 4800 2873 4812 2907
rect 4883 2904 4911 2944
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 6362 2972 6368 2984
rect 5491 2944 6368 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 6917 2975 6975 2981
rect 6512 2944 6557 2972
rect 6512 2932 6518 2944
rect 6917 2941 6929 2975
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 5718 2904 5724 2916
rect 4883 2876 5482 2904
rect 5679 2876 5724 2904
rect 4754 2867 4812 2873
rect 1762 2836 1768 2848
rect 1723 2808 1768 2836
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 2314 2836 2320 2848
rect 2275 2808 2320 2836
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 2774 2836 2780 2848
rect 2735 2808 2780 2836
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3326 2836 3332 2848
rect 3287 2808 3332 2836
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 5350 2836 5356 2848
rect 5311 2808 5356 2836
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 5454 2836 5482 2876
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 6932 2904 6960 2935
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7248 2944 7297 2972
rect 7248 2932 7254 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7524 2944 7573 2972
rect 7524 2932 7530 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 11716 2972 11744 3080
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 13262 3108 13268 3120
rect 13223 3080 13268 3108
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 13786 3108 13814 3148
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 14424 3148 17785 3176
rect 14424 3136 14430 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 21729 3179 21787 3185
rect 21729 3176 21741 3179
rect 17920 3148 21741 3176
rect 17920 3136 17926 3148
rect 15286 3108 15292 3120
rect 13786 3080 15292 3108
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 15654 3108 15660 3120
rect 15615 3080 15660 3108
rect 15654 3068 15660 3080
rect 15712 3068 15718 3120
rect 15746 3068 15752 3120
rect 15804 3108 15810 3120
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 15804 3080 17049 3108
rect 15804 3068 15810 3080
rect 17037 3077 17049 3080
rect 17083 3077 17095 3111
rect 17037 3071 17095 3077
rect 17310 3068 17316 3120
rect 17368 3108 17374 3120
rect 17368 3080 18460 3108
rect 17368 3068 17374 3080
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13722 3040 13728 3052
rect 13596 3012 13728 3040
rect 13596 3000 13602 3012
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14734 3040 14740 3052
rect 14599 3012 14740 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 14734 3000 14740 3012
rect 14792 3040 14798 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14792 3012 14933 3040
rect 14792 3000 14798 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 14921 3003 14979 3009
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 18432 3049 18460 3080
rect 18506 3068 18512 3120
rect 18564 3108 18570 3120
rect 18564 3080 20024 3108
rect 18564 3068 18570 3080
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19058 3040 19064 3052
rect 18463 3012 19064 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 19886 3040 19892 3052
rect 19751 3012 19892 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 19996 3049 20024 3080
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 11828 2975 11886 2981
rect 11828 2972 11840 2975
rect 11716 2944 11840 2972
rect 7561 2935 7619 2941
rect 11828 2941 11840 2944
rect 11874 2941 11886 2975
rect 12066 2972 12072 2984
rect 12027 2944 12072 2972
rect 11828 2935 11886 2941
rect 6052 2876 6960 2904
rect 7576 2904 7604 2935
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 12472 2975 12530 2981
rect 12472 2972 12484 2975
rect 12452 2941 12484 2972
rect 12518 2941 12530 2975
rect 12452 2935 12530 2941
rect 7742 2904 7748 2916
rect 7576 2876 7748 2904
rect 6052 2864 6058 2876
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2873 7895 2907
rect 7837 2867 7895 2873
rect 6454 2836 6460 2848
rect 5454 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 6595 2839 6653 2845
rect 6595 2805 6607 2839
rect 6641 2836 6653 2839
rect 6822 2836 6828 2848
rect 6641 2808 6828 2836
rect 6641 2805 6653 2808
rect 6595 2799 6653 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 7852 2836 7880 2867
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 8642 2907 8700 2913
rect 8642 2904 8654 2907
rect 8260 2876 8654 2904
rect 8260 2864 8266 2876
rect 8642 2873 8654 2876
rect 8688 2873 8700 2907
rect 8642 2867 8700 2873
rect 8938 2864 8944 2916
rect 8996 2864 9002 2916
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 9390 2907 9448 2913
rect 9390 2904 9402 2907
rect 9272 2876 9402 2904
rect 9272 2864 9278 2876
rect 9390 2873 9402 2876
rect 9436 2873 9448 2907
rect 9390 2867 9448 2873
rect 9493 2907 9551 2913
rect 9493 2873 9505 2907
rect 9539 2873 9551 2907
rect 10318 2904 10324 2916
rect 10279 2876 10324 2904
rect 9493 2867 9551 2873
rect 7064 2808 7880 2836
rect 8956 2836 8984 2864
rect 9508 2836 9536 2867
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 11146 2904 11152 2916
rect 11107 2876 11152 2904
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 11701 2907 11759 2913
rect 11701 2873 11713 2907
rect 11747 2904 11759 2907
rect 12342 2904 12348 2916
rect 11747 2876 12348 2904
rect 11747 2873 11759 2876
rect 11701 2867 11759 2873
rect 12342 2864 12348 2876
rect 12400 2864 12406 2916
rect 12452 2904 12480 2935
rect 12618 2932 12624 2984
rect 12676 2972 12682 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12676 2944 12909 2972
rect 12676 2932 12682 2944
rect 12897 2941 12909 2944
rect 12943 2972 12955 2975
rect 13354 2972 13360 2984
rect 12943 2944 13360 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 14458 2972 14464 2984
rect 14231 2944 14464 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2972 16911 2975
rect 17512 2972 17540 3000
rect 21192 2981 21220 3148
rect 21729 3145 21741 3148
rect 21775 3145 21787 3179
rect 21729 3139 21787 3145
rect 16899 2944 17540 2972
rect 21177 2975 21235 2981
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 21177 2941 21189 2975
rect 21223 2941 21235 2975
rect 21177 2935 21235 2941
rect 12636 2904 12664 2932
rect 13538 2904 13544 2916
rect 12452 2876 12664 2904
rect 12820 2876 13032 2904
rect 13499 2876 13544 2904
rect 8956 2808 9536 2836
rect 7064 2796 7070 2808
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 11054 2836 11060 2848
rect 9732 2808 11060 2836
rect 9732 2796 9738 2808
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11790 2836 11796 2848
rect 11296 2808 11796 2836
rect 11296 2796 11302 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12158 2796 12164 2848
rect 12216 2836 12222 2848
rect 12820 2836 12848 2876
rect 12216 2808 12848 2836
rect 13004 2836 13032 2876
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 13722 2904 13728 2916
rect 13679 2876 13728 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 15102 2904 15108 2916
rect 15063 2876 15108 2904
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 15197 2907 15255 2913
rect 15197 2873 15209 2907
rect 15243 2904 15255 2907
rect 15562 2904 15568 2916
rect 15243 2876 15568 2904
rect 15243 2873 15255 2876
rect 15197 2867 15255 2873
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 15838 2864 15844 2916
rect 15896 2904 15902 2916
rect 17862 2904 17868 2916
rect 15896 2876 17868 2904
rect 15896 2864 15902 2876
rect 17862 2864 17868 2876
rect 17920 2864 17926 2916
rect 18138 2904 18144 2916
rect 18099 2876 18144 2904
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 19518 2904 19524 2916
rect 18288 2876 19524 2904
rect 18288 2864 18294 2876
rect 19518 2864 19524 2876
rect 19576 2864 19582 2916
rect 19797 2907 19855 2913
rect 19797 2873 19809 2907
rect 19843 2873 19855 2907
rect 22094 2904 22100 2916
rect 22055 2876 22100 2904
rect 19797 2867 19855 2873
rect 13814 2836 13820 2848
rect 13004 2808 13820 2836
rect 12216 2796 12222 2808
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16761 2839 16819 2845
rect 16761 2836 16773 2839
rect 16172 2808 16773 2836
rect 16172 2796 16178 2808
rect 16761 2805 16773 2808
rect 16807 2836 16819 2839
rect 16850 2836 16856 2848
rect 16807 2808 16856 2836
rect 16807 2805 16819 2808
rect 16761 2799 16819 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 18322 2796 18328 2848
rect 18380 2836 18386 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 18380 2808 19073 2836
rect 18380 2796 18386 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 19061 2799 19119 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19812 2836 19840 2867
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 20625 2839 20683 2845
rect 20625 2836 20637 2839
rect 19392 2808 20637 2836
rect 19392 2796 19398 2808
rect 20625 2805 20637 2808
rect 20671 2836 20683 2839
rect 20806 2836 20812 2848
rect 20671 2808 20812 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 20806 2796 20812 2808
rect 20864 2836 20870 2848
rect 20993 2839 21051 2845
rect 20993 2836 21005 2839
rect 20864 2808 21005 2836
rect 20864 2796 20870 2808
rect 20993 2805 21005 2808
rect 21039 2805 21051 2839
rect 21358 2836 21364 2848
rect 21319 2808 21364 2836
rect 20993 2799 21051 2805
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 569 2635 627 2641
rect 569 2601 581 2635
rect 615 2632 627 2635
rect 2317 2635 2375 2641
rect 2317 2632 2329 2635
rect 615 2604 2329 2632
rect 615 2601 627 2604
rect 569 2595 627 2601
rect 2317 2601 2329 2604
rect 2363 2632 2375 2635
rect 2590 2632 2596 2644
rect 2363 2604 2596 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 6178 2632 6184 2644
rect 3651 2604 6184 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 7837 2635 7895 2641
rect 6564 2604 7144 2632
rect 1762 2573 1768 2576
rect 1759 2564 1768 2573
rect 1675 2536 1768 2564
rect 1759 2527 1768 2536
rect 1820 2564 1826 2576
rect 2774 2573 2780 2576
rect 2730 2567 2780 2573
rect 2730 2564 2742 2567
rect 1820 2536 2742 2564
rect 1762 2524 1768 2527
rect 1820 2524 1826 2536
rect 2730 2533 2742 2536
rect 2776 2533 2780 2567
rect 2730 2527 2780 2533
rect 2774 2524 2780 2527
rect 2832 2524 2838 2576
rect 3970 2524 3976 2576
rect 4028 2564 4034 2576
rect 4386 2567 4444 2573
rect 4386 2564 4398 2567
rect 4028 2536 4398 2564
rect 4028 2524 4034 2536
rect 4386 2533 4398 2536
rect 4432 2564 4444 2567
rect 5398 2567 5456 2573
rect 5398 2564 5410 2567
rect 4432 2536 5410 2564
rect 4432 2533 4444 2536
rect 4386 2527 4444 2533
rect 5398 2533 5410 2536
rect 5444 2564 5456 2567
rect 5718 2564 5724 2576
rect 5444 2536 5724 2564
rect 5444 2533 5456 2536
rect 5398 2527 5456 2533
rect 5718 2524 5724 2536
rect 5776 2564 5782 2576
rect 6564 2564 6592 2604
rect 7006 2564 7012 2576
rect 5776 2536 6592 2564
rect 6656 2536 7012 2564
rect 5776 2524 5782 2536
rect 198 2456 204 2508
rect 256 2496 262 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 256 2468 1409 2496
rect 256 2456 262 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3510 2496 3516 2508
rect 3467 2468 3516 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 6086 2496 6092 2508
rect 6047 2468 6092 2496
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6482 2499 6540 2505
rect 6482 2465 6494 2499
rect 6528 2496 6540 2499
rect 6656 2496 6684 2536
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 7116 2564 7144 2604
rect 7837 2601 7849 2635
rect 7883 2632 7895 2635
rect 8018 2632 8024 2644
rect 7883 2604 8024 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 10594 2592 10600 2644
rect 10652 2592 10658 2644
rect 12158 2632 12164 2644
rect 11532 2604 12164 2632
rect 7238 2567 7296 2573
rect 7238 2564 7250 2567
rect 7116 2536 7250 2564
rect 7238 2533 7250 2536
rect 7284 2564 7296 2567
rect 7650 2564 7656 2576
rect 7284 2536 7656 2564
rect 7284 2533 7296 2536
rect 7238 2527 7296 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 8110 2564 8116 2576
rect 8071 2536 8116 2564
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8846 2564 8852 2576
rect 8807 2536 8852 2564
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 8938 2524 8944 2576
rect 8996 2564 9002 2576
rect 9490 2564 9496 2576
rect 8996 2536 9041 2564
rect 9451 2536 9496 2564
rect 8996 2524 9002 2536
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 9858 2564 9864 2576
rect 9819 2536 9864 2564
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2564 10011 2567
rect 10134 2564 10140 2576
rect 9999 2536 10140 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 10612 2564 10640 2592
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 10612 2536 10793 2564
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 11532 2564 11560 2604
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 13998 2632 14004 2644
rect 12314 2604 14004 2632
rect 11379 2536 11560 2564
rect 11609 2567 11667 2573
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 11609 2533 11621 2567
rect 11655 2564 11667 2567
rect 11974 2564 11980 2576
rect 11655 2536 11980 2564
rect 11655 2533 11667 2536
rect 11609 2527 11667 2533
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 6528 2468 6684 2496
rect 6917 2499 6975 2505
rect 6528 2465 6540 2468
rect 6482 2459 6540 2465
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7834 2496 7840 2508
rect 6963 2468 7840 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 12314 2505 12342 2604
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14792 2604 15025 2632
rect 14792 2592 14798 2604
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 17310 2632 17316 2644
rect 15013 2595 15071 2601
rect 15442 2604 17316 2632
rect 12802 2564 12808 2576
rect 12715 2536 12808 2564
rect 12802 2524 12808 2536
rect 12860 2564 12866 2576
rect 15442 2564 15470 2604
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 18690 2592 18696 2644
rect 18748 2632 18754 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 18748 2604 21373 2632
rect 18748 2592 18754 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 22097 2635 22155 2641
rect 22097 2632 22109 2635
rect 21876 2604 22109 2632
rect 21876 2592 21882 2604
rect 22097 2601 22109 2604
rect 22143 2601 22155 2635
rect 22097 2595 22155 2601
rect 12860 2536 15470 2564
rect 16019 2567 16077 2573
rect 12860 2524 12866 2536
rect 16019 2533 16031 2567
rect 16065 2564 16077 2567
rect 16114 2564 16120 2576
rect 16065 2536 16120 2564
rect 16065 2533 16077 2536
rect 16019 2527 16077 2533
rect 16114 2524 16120 2536
rect 16172 2524 16178 2576
rect 16666 2524 16672 2576
rect 16724 2564 16730 2576
rect 17957 2567 18015 2573
rect 17957 2564 17969 2567
rect 16724 2536 17969 2564
rect 16724 2524 16730 2536
rect 17957 2533 17969 2536
rect 18003 2533 18015 2567
rect 18414 2564 18420 2576
rect 18375 2536 18420 2564
rect 17957 2527 18015 2533
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18506 2524 18512 2576
rect 18564 2564 18570 2576
rect 18564 2536 18609 2564
rect 18564 2524 18570 2536
rect 18874 2524 18880 2576
rect 18932 2564 18938 2576
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 18932 2536 19349 2564
rect 18932 2524 18938 2536
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19337 2527 19395 2533
rect 12299 2499 12357 2505
rect 12299 2465 12311 2499
rect 12345 2465 12357 2499
rect 12299 2459 12357 2465
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13412 2468 13645 2496
rect 13412 2456 13418 2468
rect 13633 2465 13645 2468
rect 13679 2496 13691 2499
rect 14252 2499 14310 2505
rect 13679 2468 13814 2496
rect 13679 2465 13691 2468
rect 13633 2459 13691 2465
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 900 2400 2421 2428
rect 900 2388 906 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5123 2400 6592 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 3329 2363 3387 2369
rect 3329 2329 3341 2363
rect 3375 2360 3387 2363
rect 4246 2360 4252 2372
rect 3375 2332 4252 2360
rect 3375 2329 3387 2332
rect 3329 2323 3387 2329
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 5997 2363 6055 2369
rect 5997 2360 6009 2363
rect 4402 2332 6009 2360
rect 474 2252 480 2304
rect 532 2292 538 2304
rect 4402 2292 4430 2332
rect 5997 2329 6009 2332
rect 6043 2329 6055 2363
rect 5997 2323 6055 2329
rect 532 2264 4430 2292
rect 4985 2295 5043 2301
rect 532 2252 538 2264
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 5442 2292 5448 2304
rect 5031 2264 5448 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 6273 2295 6331 2301
rect 6273 2292 6285 2295
rect 5592 2264 6285 2292
rect 5592 2252 5598 2264
rect 6273 2261 6285 2264
rect 6319 2261 6331 2295
rect 6564 2292 6592 2400
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7616 2400 8033 2428
rect 7616 2388 7622 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 10137 2431 10195 2437
rect 8711 2400 9812 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 8386 2360 8392 2372
rect 6687 2332 8392 2360
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 9784 2360 9812 2400
rect 10137 2397 10149 2431
rect 10183 2397 10195 2431
rect 10686 2428 10692 2440
rect 10647 2400 10692 2428
rect 10137 2391 10195 2397
rect 10152 2360 10180 2391
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2428 11575 2431
rect 11606 2428 11612 2440
rect 11563 2400 11612 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11790 2428 11796 2440
rect 11751 2400 11796 2428
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12894 2428 12900 2440
rect 12759 2400 12900 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13786 2428 13814 2468
rect 14252 2465 14264 2499
rect 14298 2496 14310 2499
rect 14734 2496 14740 2508
rect 14298 2468 14740 2496
rect 14298 2465 14310 2468
rect 14252 2459 14310 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 15838 2496 15844 2508
rect 15580 2468 15844 2496
rect 15580 2428 15608 2468
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 18230 2496 18236 2508
rect 16623 2468 18236 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19889 2499 19947 2505
rect 19116 2468 19161 2496
rect 19116 2456 19122 2468
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 20254 2496 20260 2508
rect 19935 2468 20260 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 21177 2499 21235 2505
rect 21177 2465 21189 2499
rect 21223 2496 21235 2499
rect 21266 2496 21272 2508
rect 21223 2468 21272 2496
rect 21223 2465 21235 2468
rect 21177 2459 21235 2465
rect 21266 2456 21272 2468
rect 21324 2456 21330 2508
rect 13786 2400 15608 2428
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 15703 2400 17049 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17218 2428 17224 2440
rect 17179 2400 17224 2428
rect 17037 2391 17095 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 20441 2431 20499 2437
rect 20441 2428 20453 2431
rect 19567 2400 20453 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 20441 2397 20453 2400
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 9784 2332 10180 2360
rect 10042 2292 10048 2304
rect 6564 2264 10048 2292
rect 6273 2255 6331 2261
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10152 2292 10180 2332
rect 11532 2332 13277 2360
rect 11532 2292 11560 2332
rect 13265 2329 13277 2332
rect 13311 2360 13323 2363
rect 15562 2360 15568 2372
rect 13311 2332 15568 2360
rect 13311 2329 13323 2332
rect 13265 2323 13323 2329
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 16850 2360 16856 2372
rect 16811 2332 16856 2360
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 19242 2360 19248 2372
rect 18564 2332 19248 2360
rect 18564 2320 18570 2332
rect 19242 2320 19248 2332
rect 19300 2360 19306 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 19300 2332 20821 2360
rect 19300 2320 19306 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 10152 2264 11560 2292
rect 12391 2295 12449 2301
rect 12391 2261 12403 2295
rect 12437 2292 12449 2295
rect 13446 2292 13452 2304
rect 12437 2264 13452 2292
rect 12437 2261 12449 2264
rect 12391 2255 12449 2261
rect 13446 2252 13452 2264
rect 13504 2252 13510 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14458 2292 14464 2304
rect 13596 2264 14464 2292
rect 13596 2252 13602 2264
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14734 2292 14740 2304
rect 14695 2264 14740 2292
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 17037 2295 17095 2301
rect 17037 2261 17049 2295
rect 17083 2292 17095 2295
rect 18782 2292 18788 2304
rect 17083 2264 18788 2292
rect 17083 2261 17095 2264
rect 17037 2255 17095 2261
rect 18782 2252 18788 2264
rect 18840 2292 18846 2304
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 18840 2264 19533 2292
rect 18840 2252 18846 2264
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19702 2292 19708 2304
rect 19663 2264 19708 2292
rect 19521 2255 19579 2261
rect 19702 2252 19708 2264
rect 19760 2252 19766 2304
rect 19794 2252 19800 2304
rect 19852 2292 19858 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 19852 2264 20085 2292
rect 19852 2252 19858 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 21726 2292 21732 2304
rect 21687 2264 21732 2292
rect 20073 2255 20131 2261
rect 21726 2252 21732 2264
rect 21784 2252 21790 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
rect 6270 2048 6276 2100
rect 6328 2088 6334 2100
rect 11514 2088 11520 2100
rect 6328 2060 11520 2088
rect 6328 2048 6334 2060
rect 11514 2048 11520 2060
rect 11572 2048 11578 2100
rect 12066 2048 12072 2100
rect 12124 2088 12130 2100
rect 16206 2088 16212 2100
rect 12124 2060 16212 2088
rect 12124 2048 12130 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 106 1980 112 2032
rect 164 2020 170 2032
rect 4798 2020 4804 2032
rect 164 1992 4804 2020
rect 164 1980 170 1992
rect 4798 1980 4804 1992
rect 4856 1980 4862 2032
rect 6730 2020 6736 2032
rect 5276 1992 6736 2020
rect 934 1912 940 1964
rect 992 1952 998 1964
rect 5276 1952 5304 1992
rect 6730 1980 6736 1992
rect 6788 2020 6794 2032
rect 8938 2020 8944 2032
rect 6788 1992 8944 2020
rect 6788 1980 6794 1992
rect 8938 1980 8944 1992
rect 8996 1980 9002 2032
rect 14458 1980 14464 2032
rect 14516 2020 14522 2032
rect 22186 2020 22192 2032
rect 14516 1992 22192 2020
rect 14516 1980 14522 1992
rect 22186 1980 22192 1992
rect 22244 1980 22250 2032
rect 992 1924 5304 1952
rect 992 1912 998 1924
rect 5350 1912 5356 1964
rect 5408 1952 5414 1964
rect 15378 1952 15384 1964
rect 5408 1924 15384 1952
rect 5408 1912 5414 1924
rect 15378 1912 15384 1924
rect 15436 1912 15442 1964
rect 4706 1844 4712 1896
rect 4764 1884 4770 1896
rect 9306 1884 9312 1896
rect 4764 1856 9312 1884
rect 4764 1844 4770 1856
rect 9306 1844 9312 1856
rect 9364 1884 9370 1896
rect 11698 1884 11704 1896
rect 9364 1856 11704 1884
rect 9364 1844 9370 1856
rect 11698 1844 11704 1856
rect 11756 1844 11762 1896
rect 4246 1776 4252 1828
rect 4304 1816 4310 1828
rect 10134 1816 10140 1828
rect 4304 1788 10140 1816
rect 4304 1776 4310 1788
rect 10134 1776 10140 1788
rect 10192 1776 10198 1828
rect 109 119 167 125
rect 109 85 121 119
rect 155 116 167 119
rect 2406 116 2412 128
rect 155 88 2412 116
rect 155 85 167 88
rect 109 79 167 85
rect 2406 76 2412 88
rect 2464 76 2470 128
rect 16758 76 16764 128
rect 16816 116 16822 128
rect 17402 116 17408 128
rect 16816 88 17408 116
rect 16816 76 16822 88
rect 17402 76 17408 88
rect 17460 76 17466 128
rect 14458 8 14464 60
rect 14516 48 14522 60
rect 21358 48 21364 60
rect 14516 20 21364 48
rect 14516 8 14522 20
rect 21358 8 21364 20
rect 21416 8 21422 60
<< via1 >>
rect 2872 23536 2924 23588
rect 15108 23536 15160 23588
rect 19340 23536 19392 23588
rect 3700 23128 3752 23180
rect 9588 23128 9640 23180
rect 2228 22992 2280 23044
rect 7196 22992 7248 23044
rect 14740 22992 14792 23044
rect 572 22924 624 22976
rect 1124 22856 1176 22908
rect 19156 22856 19208 22908
rect 940 22788 992 22840
rect 7564 22788 7616 22840
rect 7656 22788 7708 22840
rect 19248 22788 19300 22840
rect 2044 22720 2096 22772
rect 8668 22720 8720 22772
rect 9956 22720 10008 22772
rect 19340 22720 19392 22772
rect 1860 22652 1912 22704
rect 17960 22652 18012 22704
rect 1952 22584 2004 22636
rect 16212 22584 16264 22636
rect 1492 22516 1544 22568
rect 13636 22516 13688 22568
rect 14280 22448 14332 22500
rect 9220 22380 9272 22432
rect 3700 22312 3752 22364
rect 7840 22312 7892 22364
rect 8024 22312 8076 22364
rect 3240 22244 3292 22296
rect 9772 22244 9824 22296
rect 10600 22244 10652 22296
rect 15660 22244 15712 22296
rect 1032 22176 1084 22228
rect 4068 22108 4120 22160
rect 20904 22176 20956 22228
rect 10968 22108 11020 22160
rect 16948 22108 17000 22160
rect 19064 22040 19116 22092
rect 20444 21972 20496 22024
rect 3884 21904 3936 21956
rect 5540 21904 5592 21956
rect 18328 21904 18380 21956
rect 2596 21836 2648 21888
rect 4712 21836 4764 21888
rect 15476 21836 15528 21888
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 2228 21675 2280 21684
rect 2228 21641 2237 21675
rect 2237 21641 2271 21675
rect 2271 21641 2280 21675
rect 2228 21632 2280 21641
rect 4436 21632 4488 21684
rect 5908 21632 5960 21684
rect 6644 21632 6696 21684
rect 3424 21564 3476 21616
rect 4252 21607 4304 21616
rect 4252 21573 4276 21607
rect 4276 21573 4304 21607
rect 4252 21564 4304 21573
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 1216 21360 1268 21412
rect 2596 21360 2648 21412
rect 3148 21403 3200 21412
rect 3148 21369 3157 21403
rect 3157 21369 3191 21403
rect 3191 21369 3200 21403
rect 3148 21360 3200 21369
rect 2136 21292 2188 21344
rect 3424 21335 3476 21344
rect 3424 21301 3433 21335
rect 3433 21301 3467 21335
rect 3467 21301 3476 21335
rect 3424 21292 3476 21301
rect 4712 21564 4764 21616
rect 7288 21564 7340 21616
rect 10048 21632 10100 21684
rect 15384 21632 15436 21684
rect 15568 21632 15620 21684
rect 10232 21564 10284 21616
rect 12532 21564 12584 21616
rect 12900 21564 12952 21616
rect 18052 21564 18104 21616
rect 18144 21564 18196 21616
rect 18604 21607 18656 21616
rect 4804 21496 4856 21548
rect 3976 21428 4028 21480
rect 7012 21539 7064 21548
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 9588 21496 9640 21548
rect 18604 21573 18613 21607
rect 18613 21573 18647 21607
rect 18647 21573 18656 21607
rect 18604 21564 18656 21573
rect 7288 21428 7340 21480
rect 7840 21428 7892 21480
rect 8576 21428 8628 21480
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 7104 21360 7156 21412
rect 9312 21360 9364 21412
rect 9404 21360 9456 21412
rect 10416 21428 10468 21480
rect 12164 21428 12216 21480
rect 4712 21335 4764 21344
rect 4712 21301 4721 21335
rect 4721 21301 4755 21335
rect 4755 21301 4764 21335
rect 4712 21292 4764 21301
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 6000 21292 6052 21344
rect 6828 21292 6880 21344
rect 8116 21292 8168 21344
rect 11244 21360 11296 21412
rect 12532 21360 12584 21412
rect 12716 21403 12768 21412
rect 12716 21369 12725 21403
rect 12725 21369 12759 21403
rect 12759 21369 12768 21403
rect 12716 21360 12768 21369
rect 12900 21360 12952 21412
rect 11060 21292 11112 21344
rect 11336 21335 11388 21344
rect 11336 21301 11345 21335
rect 11345 21301 11379 21335
rect 11379 21301 11388 21335
rect 15016 21360 15068 21412
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 15752 21360 15804 21412
rect 11336 21292 11388 21301
rect 15108 21292 15160 21344
rect 16028 21292 16080 21344
rect 16764 21292 16816 21344
rect 17776 21471 17828 21480
rect 17776 21437 17785 21471
rect 17785 21437 17819 21471
rect 17819 21437 17828 21471
rect 17776 21428 17828 21437
rect 18144 21428 18196 21480
rect 18788 21496 18840 21548
rect 20720 21428 20772 21480
rect 16948 21360 17000 21412
rect 18328 21403 18380 21412
rect 18328 21369 18337 21403
rect 18337 21369 18371 21403
rect 18371 21369 18380 21403
rect 18328 21360 18380 21369
rect 17500 21292 17552 21344
rect 18604 21292 18656 21344
rect 18696 21292 18748 21344
rect 19432 21292 19484 21344
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 1400 21088 1452 21140
rect 4252 21088 4304 21140
rect 2596 21063 2648 21072
rect 2596 21029 2605 21063
rect 2605 21029 2639 21063
rect 2639 21029 2648 21063
rect 2596 21020 2648 21029
rect 3148 21020 3200 21072
rect 4344 21020 4396 21072
rect 4620 21020 4672 21072
rect 1768 20995 1820 21004
rect 1768 20961 1777 20995
rect 1777 20961 1811 20995
rect 1811 20961 1820 20995
rect 1768 20952 1820 20961
rect 2780 20952 2832 21004
rect 3424 20952 3476 21004
rect 3516 20884 3568 20936
rect 2412 20816 2464 20868
rect 3976 20816 4028 20868
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 5080 21088 5132 21140
rect 5908 21131 5960 21140
rect 5908 21097 5917 21131
rect 5917 21097 5951 21131
rect 5951 21097 5960 21131
rect 5908 21088 5960 21097
rect 7840 21088 7892 21140
rect 8760 21088 8812 21140
rect 14004 21131 14056 21140
rect 5816 21020 5868 21072
rect 7196 21020 7248 21072
rect 9588 21020 9640 21072
rect 6184 20952 6236 21004
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 5724 20884 5776 20936
rect 5908 20884 5960 20936
rect 7472 20952 7524 21004
rect 7932 20995 7984 21004
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 7564 20884 7616 20936
rect 9220 20952 9272 21004
rect 9956 20995 10008 21004
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 11888 21020 11940 21072
rect 11428 20952 11480 21004
rect 4344 20816 4396 20868
rect 4712 20816 4764 20868
rect 5356 20816 5408 20868
rect 5632 20816 5684 20868
rect 7656 20816 7708 20868
rect 11336 20927 11388 20936
rect 8484 20816 8536 20868
rect 9680 20816 9732 20868
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11980 20927 12032 20936
rect 11336 20884 11388 20893
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 14004 21097 14013 21131
rect 14013 21097 14047 21131
rect 14047 21097 14056 21131
rect 14004 21088 14056 21097
rect 14556 21088 14608 21140
rect 15016 21131 15068 21140
rect 15016 21097 15025 21131
rect 15025 21097 15059 21131
rect 15059 21097 15068 21131
rect 15016 21088 15068 21097
rect 15292 21088 15344 21140
rect 15568 21088 15620 21140
rect 15476 21063 15528 21072
rect 15476 21029 15485 21063
rect 15485 21029 15519 21063
rect 15519 21029 15528 21063
rect 15476 21020 15528 21029
rect 16764 21020 16816 21072
rect 18052 21020 18104 21072
rect 18512 21063 18564 21072
rect 18512 21029 18521 21063
rect 18521 21029 18555 21063
rect 18555 21029 18564 21063
rect 18512 21020 18564 21029
rect 18972 21020 19024 21072
rect 20812 21020 20864 21072
rect 21364 21020 21416 21072
rect 12808 20952 12860 21004
rect 12992 20952 13044 21004
rect 14832 20952 14884 21004
rect 4528 20748 4580 20800
rect 5448 20748 5500 20800
rect 7196 20748 7248 20800
rect 8944 20748 8996 20800
rect 12992 20816 13044 20868
rect 14924 20884 14976 20936
rect 15752 20884 15804 20936
rect 16672 20884 16724 20936
rect 21272 20884 21324 20936
rect 21548 20859 21600 20868
rect 21548 20825 21557 20859
rect 21557 20825 21591 20859
rect 21591 20825 21600 20859
rect 21548 20816 21600 20825
rect 10692 20791 10744 20800
rect 10692 20757 10701 20791
rect 10701 20757 10735 20791
rect 10735 20757 10744 20791
rect 10692 20748 10744 20757
rect 11428 20748 11480 20800
rect 12624 20791 12676 20800
rect 12624 20757 12633 20791
rect 12633 20757 12667 20791
rect 12667 20757 12676 20791
rect 12624 20748 12676 20757
rect 14740 20748 14792 20800
rect 16120 20748 16172 20800
rect 17684 20748 17736 20800
rect 18696 20748 18748 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 3424 20544 3476 20596
rect 4620 20587 4672 20596
rect 4620 20553 4629 20587
rect 4629 20553 4663 20587
rect 4663 20553 4672 20587
rect 4620 20544 4672 20553
rect 5448 20544 5500 20596
rect 5724 20587 5776 20596
rect 5724 20553 5733 20587
rect 5733 20553 5767 20587
rect 5767 20553 5776 20587
rect 5724 20544 5776 20553
rect 7288 20544 7340 20596
rect 9956 20544 10008 20596
rect 13728 20544 13780 20596
rect 18512 20544 18564 20596
rect 20812 20587 20864 20596
rect 20812 20553 20821 20587
rect 20821 20553 20855 20587
rect 20855 20553 20864 20587
rect 20812 20544 20864 20553
rect 21456 20587 21508 20596
rect 21456 20553 21465 20587
rect 21465 20553 21499 20587
rect 21499 20553 21508 20587
rect 21456 20544 21508 20553
rect 3332 20476 3384 20528
rect 4160 20476 4212 20528
rect 5908 20476 5960 20528
rect 6828 20476 6880 20528
rect 8300 20476 8352 20528
rect 9588 20519 9640 20528
rect 4620 20408 4672 20460
rect 4896 20408 4948 20460
rect 9588 20485 9597 20519
rect 9597 20485 9631 20519
rect 9631 20485 9640 20519
rect 9588 20476 9640 20485
rect 9680 20476 9732 20528
rect 11060 20476 11112 20528
rect 12348 20476 12400 20528
rect 112 20204 164 20256
rect 3424 20340 3476 20392
rect 3608 20340 3660 20392
rect 6828 20340 6880 20392
rect 4160 20272 4212 20324
rect 4988 20272 5040 20324
rect 5724 20272 5776 20324
rect 6368 20272 6420 20324
rect 7840 20340 7892 20392
rect 8300 20340 8352 20392
rect 9036 20340 9088 20392
rect 7288 20272 7340 20324
rect 7932 20272 7984 20324
rect 2688 20204 2740 20256
rect 3700 20204 3752 20256
rect 3884 20204 3936 20256
rect 4896 20204 4948 20256
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 6920 20204 6972 20256
rect 9772 20272 9824 20324
rect 10784 20340 10836 20392
rect 11888 20383 11940 20392
rect 11888 20349 11897 20383
rect 11897 20349 11931 20383
rect 11931 20349 11940 20383
rect 11888 20340 11940 20349
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 12716 20340 12768 20392
rect 14004 20408 14056 20460
rect 16856 20476 16908 20528
rect 16948 20476 17000 20528
rect 20076 20476 20128 20528
rect 10416 20315 10468 20324
rect 10048 20204 10100 20256
rect 10416 20281 10425 20315
rect 10425 20281 10459 20315
rect 10459 20281 10468 20315
rect 10416 20272 10468 20281
rect 11704 20272 11756 20324
rect 14556 20383 14608 20392
rect 14556 20349 14565 20383
rect 14565 20349 14599 20383
rect 14599 20349 14608 20383
rect 14556 20340 14608 20349
rect 14740 20340 14792 20392
rect 15200 20340 15252 20392
rect 18880 20408 18932 20460
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 15384 20272 15436 20324
rect 16764 20272 16816 20324
rect 18420 20340 18472 20392
rect 22652 20476 22704 20528
rect 21456 20340 21508 20392
rect 19524 20272 19576 20324
rect 20536 20272 20588 20324
rect 21364 20272 21416 20324
rect 12808 20204 12860 20256
rect 13544 20204 13596 20256
rect 14188 20204 14240 20256
rect 15660 20247 15712 20256
rect 15660 20213 15669 20247
rect 15669 20213 15703 20247
rect 15703 20213 15712 20247
rect 15660 20204 15712 20213
rect 16672 20204 16724 20256
rect 18144 20247 18196 20256
rect 18144 20213 18153 20247
rect 18153 20213 18187 20247
rect 18187 20213 18196 20247
rect 18144 20204 18196 20213
rect 18972 20204 19024 20256
rect 19616 20204 19668 20256
rect 19892 20204 19944 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 1676 20000 1728 20052
rect 1768 20000 1820 20052
rect 3792 20000 3844 20052
rect 2320 19864 2372 19916
rect 3700 19932 3752 19984
rect 3976 19932 4028 19984
rect 4160 19932 4212 19984
rect 2596 19864 2648 19916
rect 1768 19796 1820 19848
rect 3056 19796 3108 19848
rect 3976 19796 4028 19848
rect 4528 19864 4580 19916
rect 4988 20000 5040 20052
rect 5540 20000 5592 20052
rect 5908 20043 5960 20052
rect 5908 20009 5917 20043
rect 5917 20009 5951 20043
rect 5951 20009 5960 20043
rect 5908 20000 5960 20009
rect 6092 20043 6144 20052
rect 6092 20009 6101 20043
rect 6101 20009 6135 20043
rect 6135 20009 6144 20043
rect 6092 20000 6144 20009
rect 6460 20000 6512 20052
rect 6828 20000 6880 20052
rect 15384 20043 15436 20052
rect 5816 19932 5868 19984
rect 7288 19932 7340 19984
rect 7564 19932 7616 19984
rect 7748 19932 7800 19984
rect 11152 19932 11204 19984
rect 6368 19864 6420 19916
rect 8300 19907 8352 19916
rect 8300 19873 8309 19907
rect 8309 19873 8343 19907
rect 8343 19873 8352 19907
rect 8300 19864 8352 19873
rect 8392 19864 8444 19916
rect 8944 19907 8996 19916
rect 8944 19873 8953 19907
rect 8953 19873 8987 19907
rect 8987 19873 8996 19907
rect 8944 19864 8996 19873
rect 9588 19864 9640 19916
rect 9864 19864 9916 19916
rect 11060 19864 11112 19916
rect 12072 19932 12124 19984
rect 12256 19932 12308 19984
rect 15384 20009 15393 20043
rect 15393 20009 15427 20043
rect 15427 20009 15436 20043
rect 15384 20000 15436 20009
rect 16120 20000 16172 20052
rect 12808 19907 12860 19916
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 7656 19796 7708 19848
rect 8116 19796 8168 19848
rect 12808 19873 12817 19907
rect 12817 19873 12851 19907
rect 12851 19873 12860 19907
rect 12808 19864 12860 19873
rect 12900 19907 12952 19916
rect 12900 19873 12909 19907
rect 12909 19873 12943 19907
rect 12943 19873 12952 19907
rect 15660 19932 15712 19984
rect 16580 19932 16632 19984
rect 21640 20000 21692 20052
rect 12900 19864 12952 19873
rect 13360 19864 13412 19916
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 12348 19796 12400 19848
rect 13452 19796 13504 19848
rect 15016 19864 15068 19916
rect 15568 19907 15620 19916
rect 15568 19873 15577 19907
rect 15577 19873 15611 19907
rect 15611 19873 15620 19907
rect 15568 19864 15620 19873
rect 14004 19796 14056 19848
rect 15476 19796 15528 19848
rect 2504 19771 2556 19780
rect 2504 19737 2513 19771
rect 2513 19737 2547 19771
rect 2547 19737 2556 19771
rect 2504 19728 2556 19737
rect 3608 19728 3660 19780
rect 9496 19728 9548 19780
rect 10048 19728 10100 19780
rect 1216 19660 1268 19712
rect 2228 19703 2280 19712
rect 2228 19669 2237 19703
rect 2237 19669 2271 19703
rect 2271 19669 2280 19703
rect 2228 19660 2280 19669
rect 2320 19660 2372 19712
rect 2872 19660 2924 19712
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 4252 19660 4304 19712
rect 4620 19660 4672 19712
rect 5724 19660 5776 19712
rect 6368 19660 6420 19712
rect 7288 19660 7340 19712
rect 8760 19660 8812 19712
rect 9956 19660 10008 19712
rect 10784 19703 10836 19712
rect 10784 19669 10793 19703
rect 10793 19669 10827 19703
rect 10827 19669 10836 19703
rect 10784 19660 10836 19669
rect 11428 19660 11480 19712
rect 12256 19660 12308 19712
rect 13636 19728 13688 19780
rect 14188 19728 14240 19780
rect 14556 19728 14608 19780
rect 16856 19907 16908 19916
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 17408 19907 17460 19916
rect 17408 19873 17417 19907
rect 17417 19873 17451 19907
rect 17451 19873 17460 19907
rect 17408 19864 17460 19873
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19984 19864 20036 19916
rect 20812 19864 20864 19916
rect 15844 19728 15896 19780
rect 18328 19728 18380 19780
rect 12716 19660 12768 19712
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 16028 19660 16080 19712
rect 16672 19660 16724 19712
rect 21364 19660 21416 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 2228 19456 2280 19508
rect 2136 19388 2188 19440
rect 2596 19388 2648 19440
rect 2780 19431 2832 19440
rect 2780 19397 2789 19431
rect 2789 19397 2823 19431
rect 2823 19397 2832 19431
rect 2780 19388 2832 19397
rect 3056 19456 3108 19508
rect 3884 19456 3936 19508
rect 4804 19456 4856 19508
rect 5448 19456 5500 19508
rect 6368 19456 6420 19508
rect 4712 19388 4764 19440
rect 5264 19388 5316 19440
rect 6460 19388 6512 19440
rect 7012 19431 7064 19440
rect 7012 19397 7021 19431
rect 7021 19397 7055 19431
rect 7055 19397 7064 19431
rect 7012 19388 7064 19397
rect 7472 19456 7524 19508
rect 9588 19456 9640 19508
rect 11152 19456 11204 19508
rect 11612 19456 11664 19508
rect 13544 19499 13596 19508
rect 13544 19465 13553 19499
rect 13553 19465 13587 19499
rect 13587 19465 13596 19499
rect 13544 19456 13596 19465
rect 13912 19456 13964 19508
rect 14096 19456 14148 19508
rect 15384 19456 15436 19508
rect 16672 19456 16724 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 20628 19456 20680 19508
rect 1216 19252 1268 19304
rect 2136 19252 2188 19304
rect 2780 19294 2832 19346
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 4160 19252 4212 19304
rect 4620 19320 4672 19372
rect 5816 19320 5868 19372
rect 6184 19320 6236 19372
rect 8576 19388 8628 19440
rect 4436 19295 4488 19304
rect 4436 19261 4445 19295
rect 4445 19261 4479 19295
rect 4479 19261 4488 19295
rect 4436 19252 4488 19261
rect 4528 19252 4580 19304
rect 6644 19252 6696 19304
rect 6920 19252 6972 19304
rect 7196 19252 7248 19304
rect 7932 19295 7984 19304
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 9036 19320 9088 19372
rect 11244 19320 11296 19372
rect 12072 19320 12124 19372
rect 3700 19184 3752 19236
rect 5908 19184 5960 19236
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 2872 19116 2924 19168
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 6644 19116 6696 19168
rect 7196 19116 7248 19168
rect 8024 19159 8076 19168
rect 8024 19125 8033 19159
rect 8033 19125 8067 19159
rect 8067 19125 8076 19159
rect 8024 19116 8076 19125
rect 8300 19116 8352 19168
rect 10140 19184 10192 19236
rect 12440 19295 12492 19304
rect 12440 19261 12449 19295
rect 12449 19261 12483 19295
rect 12483 19261 12492 19295
rect 13820 19320 13872 19372
rect 12440 19252 12492 19261
rect 13084 19252 13136 19304
rect 14188 19320 14240 19372
rect 17776 19388 17828 19440
rect 18512 19388 18564 19440
rect 13176 19184 13228 19236
rect 13912 19184 13964 19236
rect 11060 19116 11112 19168
rect 11888 19116 11940 19168
rect 12256 19116 12308 19168
rect 13268 19116 13320 19168
rect 14464 19184 14516 19236
rect 15844 19252 15896 19304
rect 16488 19320 16540 19372
rect 17500 19252 17552 19304
rect 15752 19184 15804 19236
rect 18144 19227 18196 19236
rect 18144 19193 18153 19227
rect 18153 19193 18187 19227
rect 18187 19193 18196 19227
rect 18144 19184 18196 19193
rect 18236 19227 18288 19236
rect 18236 19193 18245 19227
rect 18245 19193 18279 19227
rect 18279 19193 18288 19227
rect 18236 19184 18288 19193
rect 19984 19252 20036 19304
rect 20444 19252 20496 19304
rect 23572 19252 23624 19304
rect 14740 19116 14792 19168
rect 15476 19116 15528 19168
rect 15660 19159 15712 19168
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 17408 19116 17460 19168
rect 18604 19116 18656 19168
rect 19524 19159 19576 19168
rect 19524 19125 19533 19159
rect 19533 19125 19567 19159
rect 19567 19125 19576 19159
rect 19524 19116 19576 19125
rect 20352 19116 20404 19168
rect 20812 19116 20864 19168
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 20 18912 72 18964
rect 5724 18912 5776 18964
rect 7288 18912 7340 18964
rect 2136 18844 2188 18896
rect 3608 18844 3660 18896
rect 2228 18776 2280 18828
rect 2044 18640 2096 18692
rect 3240 18776 3292 18828
rect 3884 18776 3936 18828
rect 4344 18844 4396 18896
rect 4436 18776 4488 18828
rect 5908 18844 5960 18896
rect 7564 18844 7616 18896
rect 6184 18819 6236 18828
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 7196 18776 7248 18828
rect 7656 18819 7708 18828
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 3792 18708 3844 18760
rect 3884 18683 3936 18692
rect 3884 18649 3893 18683
rect 3893 18649 3927 18683
rect 3927 18649 3936 18683
rect 5356 18708 5408 18760
rect 6460 18708 6512 18760
rect 7656 18785 7665 18819
rect 7665 18785 7699 18819
rect 7699 18785 7708 18819
rect 7656 18776 7708 18785
rect 8392 18912 8444 18964
rect 8576 18912 8628 18964
rect 7840 18844 7892 18896
rect 12624 18912 12676 18964
rect 13176 18912 13228 18964
rect 14188 18912 14240 18964
rect 15844 18912 15896 18964
rect 10324 18844 10376 18896
rect 12072 18887 12124 18896
rect 12072 18853 12081 18887
rect 12081 18853 12115 18887
rect 12115 18853 12124 18887
rect 12072 18844 12124 18853
rect 7564 18708 7616 18760
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 8576 18708 8628 18760
rect 9680 18776 9732 18828
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 11428 18776 11480 18828
rect 12808 18844 12860 18896
rect 12624 18776 12676 18828
rect 13084 18819 13136 18828
rect 9956 18708 10008 18760
rect 3884 18640 3936 18649
rect 6184 18640 6236 18692
rect 6552 18640 6604 18692
rect 1676 18615 1728 18624
rect 1676 18581 1685 18615
rect 1685 18581 1719 18615
rect 1719 18581 1728 18615
rect 1676 18572 1728 18581
rect 4804 18572 4856 18624
rect 5540 18572 5592 18624
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 8392 18572 8444 18624
rect 8944 18572 8996 18624
rect 11152 18640 11204 18692
rect 12532 18708 12584 18760
rect 12072 18640 12124 18692
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 13912 18844 13964 18896
rect 14924 18844 14976 18896
rect 16028 18887 16080 18896
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 15016 18776 15068 18828
rect 15200 18776 15252 18828
rect 16028 18853 16037 18887
rect 16037 18853 16071 18887
rect 16071 18853 16080 18887
rect 16028 18844 16080 18853
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 17224 18776 17276 18828
rect 17408 18844 17460 18896
rect 18144 18912 18196 18964
rect 20812 18844 20864 18896
rect 16396 18708 16448 18760
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 13820 18640 13872 18692
rect 14188 18640 14240 18692
rect 18236 18776 18288 18828
rect 18420 18776 18472 18828
rect 19432 18819 19484 18828
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 19616 18708 19668 18760
rect 20628 18708 20680 18760
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 12808 18572 12860 18624
rect 14096 18572 14148 18624
rect 14556 18572 14608 18624
rect 16028 18572 16080 18624
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 3424 18411 3476 18420
rect 3424 18377 3448 18411
rect 3448 18377 3476 18411
rect 3424 18368 3476 18377
rect 3608 18368 3660 18420
rect 3884 18411 3936 18420
rect 3884 18377 3893 18411
rect 3893 18377 3927 18411
rect 3927 18377 3936 18411
rect 3884 18368 3936 18377
rect 3976 18368 4028 18420
rect 4344 18411 4396 18420
rect 4344 18377 4353 18411
rect 4353 18377 4387 18411
rect 4387 18377 4396 18411
rect 4344 18368 4396 18377
rect 3240 18300 3292 18352
rect 5908 18411 5960 18420
rect 5908 18377 5917 18411
rect 5917 18377 5951 18411
rect 5951 18377 5960 18411
rect 5908 18368 5960 18377
rect 6184 18411 6236 18420
rect 6184 18377 6193 18411
rect 6193 18377 6227 18411
rect 6227 18377 6236 18411
rect 6184 18368 6236 18377
rect 7564 18368 7616 18420
rect 9496 18368 9548 18420
rect 9680 18368 9732 18420
rect 9956 18368 10008 18420
rect 11060 18368 11112 18420
rect 11152 18368 11204 18420
rect 12348 18368 12400 18420
rect 4896 18300 4948 18352
rect 3332 18232 3384 18284
rect 3976 18232 4028 18284
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 2044 18164 2096 18216
rect 3424 18164 3476 18216
rect 4252 18164 4304 18216
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 5448 18232 5500 18284
rect 10232 18300 10284 18352
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 7380 18232 7432 18284
rect 7564 18232 7616 18284
rect 7196 18164 7248 18216
rect 940 18028 992 18080
rect 2780 18096 2832 18148
rect 3240 18139 3292 18148
rect 3240 18105 3249 18139
rect 3249 18105 3283 18139
rect 3283 18105 3292 18139
rect 3240 18096 3292 18105
rect 3700 18096 3752 18148
rect 7012 18096 7064 18148
rect 7564 18139 7616 18148
rect 7564 18105 7573 18139
rect 7573 18105 7607 18139
rect 7607 18105 7616 18139
rect 7564 18096 7616 18105
rect 4344 18028 4396 18080
rect 7840 18164 7892 18216
rect 11428 18232 11480 18284
rect 7840 18071 7892 18080
rect 7840 18037 7849 18071
rect 7849 18037 7883 18071
rect 7883 18037 7892 18071
rect 7840 18028 7892 18037
rect 8300 18096 8352 18148
rect 9036 18164 9088 18216
rect 9956 18164 10008 18216
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 15200 18368 15252 18420
rect 15476 18368 15528 18420
rect 16948 18411 17000 18420
rect 16948 18377 16957 18411
rect 16957 18377 16991 18411
rect 16991 18377 17000 18411
rect 16948 18368 17000 18377
rect 19248 18368 19300 18420
rect 19708 18368 19760 18420
rect 20076 18368 20128 18420
rect 14096 18300 14148 18352
rect 16856 18300 16908 18352
rect 18512 18300 18564 18352
rect 14556 18232 14608 18284
rect 19800 18232 19852 18284
rect 20260 18300 20312 18352
rect 12900 18207 12952 18216
rect 8852 18028 8904 18080
rect 10048 18096 10100 18148
rect 10600 18096 10652 18148
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 14464 18207 14516 18216
rect 12716 18096 12768 18148
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 14740 18096 14792 18148
rect 16304 18164 16356 18216
rect 18144 18164 18196 18216
rect 18328 18164 18380 18216
rect 20812 18300 20864 18352
rect 22192 18164 22244 18216
rect 9588 18028 9640 18080
rect 10232 18028 10284 18080
rect 11060 18028 11112 18080
rect 11796 18028 11848 18080
rect 12348 18028 12400 18080
rect 13820 18028 13872 18080
rect 14096 18071 14148 18080
rect 14096 18037 14105 18071
rect 14105 18037 14139 18071
rect 14139 18037 14148 18071
rect 14096 18028 14148 18037
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 15200 18028 15252 18080
rect 16764 18096 16816 18148
rect 17224 18096 17276 18148
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 17868 18028 17920 18080
rect 18420 18028 18472 18080
rect 19248 18028 19300 18080
rect 20536 18096 20588 18148
rect 20628 18096 20680 18148
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 1676 17824 1728 17876
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 3148 17756 3200 17808
rect 3332 17756 3384 17808
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 2872 17688 2924 17740
rect 4712 17824 4764 17876
rect 6644 17867 6696 17876
rect 6644 17833 6653 17867
rect 6653 17833 6687 17867
rect 6687 17833 6696 17867
rect 6644 17824 6696 17833
rect 6828 17824 6880 17876
rect 7472 17824 7524 17876
rect 8300 17824 8352 17876
rect 8852 17824 8904 17876
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 11520 17824 11572 17876
rect 12440 17824 12492 17876
rect 15568 17824 15620 17876
rect 16304 17867 16356 17876
rect 16304 17833 16313 17867
rect 16313 17833 16347 17867
rect 16347 17833 16356 17867
rect 16304 17824 16356 17833
rect 17592 17824 17644 17876
rect 18052 17824 18104 17876
rect 18328 17824 18380 17876
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 19984 17824 20036 17876
rect 4620 17756 4672 17808
rect 10324 17756 10376 17808
rect 10876 17756 10928 17808
rect 4896 17688 4948 17740
rect 5264 17688 5316 17740
rect 6828 17731 6880 17740
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 3700 17620 3752 17672
rect 5172 17620 5224 17672
rect 2228 17552 2280 17604
rect 4252 17552 4304 17604
rect 1492 17484 1544 17536
rect 3240 17484 3292 17536
rect 4068 17484 4120 17536
rect 4436 17484 4488 17536
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 6920 17688 6972 17740
rect 5632 17663 5684 17672
rect 5632 17629 5641 17663
rect 5641 17629 5675 17663
rect 5675 17629 5684 17663
rect 5632 17620 5684 17629
rect 6276 17620 6328 17672
rect 5816 17552 5868 17604
rect 9220 17688 9272 17740
rect 9680 17688 9732 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 11612 17731 11664 17740
rect 11612 17697 11621 17731
rect 11621 17697 11655 17731
rect 11655 17697 11664 17731
rect 11612 17688 11664 17697
rect 12716 17756 12768 17808
rect 12900 17756 12952 17808
rect 12624 17731 12676 17740
rect 12624 17697 12633 17731
rect 12633 17697 12667 17731
rect 12667 17697 12676 17731
rect 12624 17688 12676 17697
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 13544 17688 13596 17740
rect 14924 17756 14976 17808
rect 13820 17688 13872 17740
rect 14464 17688 14516 17740
rect 14648 17688 14700 17740
rect 15476 17731 15528 17740
rect 15476 17697 15485 17731
rect 15485 17697 15519 17731
rect 15519 17697 15528 17731
rect 15476 17688 15528 17697
rect 17500 17731 17552 17740
rect 5724 17484 5776 17536
rect 7656 17527 7708 17536
rect 7656 17493 7665 17527
rect 7665 17493 7699 17527
rect 7699 17493 7708 17527
rect 12808 17620 12860 17672
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 15108 17620 15160 17672
rect 17500 17697 17509 17731
rect 17509 17697 17543 17731
rect 17543 17697 17552 17731
rect 17500 17688 17552 17697
rect 18604 17688 18656 17740
rect 19064 17756 19116 17808
rect 20076 17756 20128 17808
rect 20812 17688 20864 17740
rect 21456 17731 21508 17740
rect 21456 17697 21465 17731
rect 21465 17697 21499 17731
rect 21499 17697 21508 17731
rect 21456 17688 21508 17697
rect 10048 17552 10100 17604
rect 10876 17552 10928 17604
rect 15844 17552 15896 17604
rect 21456 17552 21508 17604
rect 7656 17484 7708 17493
rect 8852 17484 8904 17536
rect 9312 17484 9364 17536
rect 9956 17484 10008 17536
rect 12624 17484 12676 17536
rect 14556 17527 14608 17536
rect 14556 17493 14565 17527
rect 14565 17493 14599 17527
rect 14599 17493 14608 17527
rect 14556 17484 14608 17493
rect 16764 17527 16816 17536
rect 16764 17493 16773 17527
rect 16773 17493 16807 17527
rect 16807 17493 16816 17527
rect 16764 17484 16816 17493
rect 18604 17484 18656 17536
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 20 17459 72 17468
rect 20 17425 29 17459
rect 29 17425 63 17459
rect 63 17425 72 17459
rect 20 17416 72 17425
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 2228 17280 2280 17332
rect 2688 17280 2740 17332
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 4344 17280 4396 17332
rect 6184 17280 6236 17332
rect 6460 17280 6512 17332
rect 8116 17280 8168 17332
rect 8300 17280 8352 17332
rect 2044 17212 2096 17264
rect 4712 17212 4764 17264
rect 6828 17212 6880 17264
rect 7472 17255 7524 17264
rect 7472 17221 7481 17255
rect 7481 17221 7515 17255
rect 7515 17221 7524 17255
rect 9220 17280 9272 17332
rect 9680 17280 9732 17332
rect 13544 17323 13596 17332
rect 13544 17289 13553 17323
rect 13553 17289 13587 17323
rect 13587 17289 13596 17323
rect 13544 17280 13596 17289
rect 7472 17212 7524 17221
rect 2412 17076 2464 17128
rect 2872 17076 2924 17128
rect 4160 17144 4212 17196
rect 4252 17144 4304 17196
rect 3976 17076 4028 17128
rect 4436 17076 4488 17128
rect 6184 17144 6236 17196
rect 7012 17144 7064 17196
rect 7380 17144 7432 17196
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 9680 17144 9732 17196
rect 10876 17144 10928 17196
rect 5724 17119 5776 17128
rect 5724 17085 5733 17119
rect 5733 17085 5767 17119
rect 5767 17085 5776 17119
rect 5724 17076 5776 17085
rect 7840 17076 7892 17128
rect 11612 17212 11664 17264
rect 12624 17212 12676 17264
rect 13360 17212 13412 17264
rect 17500 17280 17552 17332
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 18696 17280 18748 17332
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 19340 17280 19392 17332
rect 21364 17323 21416 17332
rect 11244 17144 11296 17196
rect 4344 17051 4396 17060
rect 4344 17017 4353 17051
rect 4353 17017 4387 17051
rect 4387 17017 4396 17051
rect 4344 17008 4396 17017
rect 4896 17008 4948 17060
rect 5264 17008 5316 17060
rect 5908 17051 5960 17060
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 4436 16983 4488 16992
rect 4436 16949 4445 16983
rect 4445 16949 4479 16983
rect 4479 16949 4488 16983
rect 4436 16940 4488 16949
rect 5172 16940 5224 16992
rect 5448 16940 5500 16992
rect 5908 17017 5917 17051
rect 5917 17017 5951 17051
rect 5951 17017 5960 17051
rect 5908 17008 5960 17017
rect 7012 17051 7064 17060
rect 7012 17017 7021 17051
rect 7021 17017 7055 17051
rect 7055 17017 7064 17051
rect 7012 17008 7064 17017
rect 8484 17008 8536 17060
rect 11796 17076 11848 17128
rect 6828 16940 6880 16992
rect 7196 16940 7248 16992
rect 8300 16983 8352 16992
rect 8300 16949 8309 16983
rect 8309 16949 8343 16983
rect 8343 16949 8352 16983
rect 11612 17008 11664 17060
rect 8300 16940 8352 16949
rect 11060 16940 11112 16992
rect 12716 17076 12768 17128
rect 14464 17119 14516 17128
rect 14464 17085 14473 17119
rect 14473 17085 14507 17119
rect 14507 17085 14516 17119
rect 14464 17076 14516 17085
rect 15844 17144 15896 17196
rect 15936 17144 15988 17196
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 17776 17076 17828 17128
rect 21364 17289 21373 17323
rect 21373 17289 21407 17323
rect 21407 17289 21416 17323
rect 21364 17280 21416 17289
rect 21456 17280 21508 17332
rect 20260 17076 20312 17128
rect 13176 17051 13228 17060
rect 13176 17017 13185 17051
rect 13185 17017 13219 17051
rect 13219 17017 13228 17051
rect 13176 17008 13228 17017
rect 13544 17008 13596 17060
rect 15476 17008 15528 17060
rect 15936 17008 15988 17060
rect 16304 17051 16356 17060
rect 16304 17017 16313 17051
rect 16313 17017 16347 17051
rect 16347 17017 16356 17051
rect 16304 17008 16356 17017
rect 18696 17008 18748 17060
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15016 16940 15068 16992
rect 15384 16940 15436 16992
rect 19524 16940 19576 16992
rect 20812 16940 20864 16992
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 664 16779 716 16788
rect 664 16745 673 16779
rect 673 16745 707 16779
rect 707 16745 716 16779
rect 664 16736 716 16745
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 2412 16779 2464 16788
rect 2412 16745 2421 16779
rect 2421 16745 2455 16779
rect 2455 16745 2464 16779
rect 2412 16736 2464 16745
rect 3976 16736 4028 16788
rect 6092 16668 6144 16720
rect 6920 16668 6972 16720
rect 7288 16668 7340 16720
rect 7840 16668 7892 16720
rect 8116 16668 8168 16720
rect 8576 16668 8628 16720
rect 8944 16668 8996 16720
rect 10324 16736 10376 16788
rect 10876 16736 10928 16788
rect 12716 16736 12768 16788
rect 14464 16736 14516 16788
rect 15108 16779 15160 16788
rect 15108 16745 15117 16779
rect 15117 16745 15151 16779
rect 15151 16745 15160 16779
rect 15108 16736 15160 16745
rect 15384 16736 15436 16788
rect 18328 16779 18380 16788
rect 18328 16745 18337 16779
rect 18337 16745 18371 16779
rect 18371 16745 18380 16779
rect 18328 16736 18380 16745
rect 18880 16779 18932 16788
rect 18880 16745 18889 16779
rect 18889 16745 18923 16779
rect 18923 16745 18932 16779
rect 18880 16736 18932 16745
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 2136 16600 2188 16652
rect 3332 16600 3384 16652
rect 4528 16600 4580 16652
rect 5356 16600 5408 16652
rect 5448 16600 5500 16652
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 11152 16600 11204 16652
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 11612 16600 11664 16652
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 13912 16668 13964 16720
rect 17868 16668 17920 16720
rect 20720 16668 20772 16720
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 16028 16600 16080 16652
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 17224 16600 17276 16652
rect 18696 16643 18748 16652
rect 2228 16532 2280 16584
rect 6828 16532 6880 16584
rect 7472 16532 7524 16584
rect 9312 16532 9364 16584
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 8484 16464 8536 16516
rect 9220 16464 9272 16516
rect 9588 16464 9640 16516
rect 12624 16532 12676 16584
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 14464 16532 14516 16584
rect 16396 16532 16448 16584
rect 18696 16609 18705 16643
rect 18705 16609 18739 16643
rect 18739 16609 18748 16643
rect 18696 16600 18748 16609
rect 19432 16532 19484 16584
rect 20812 16532 20864 16584
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 11152 16464 11204 16516
rect 14832 16464 14884 16516
rect 4160 16396 4212 16448
rect 5724 16396 5776 16448
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 7012 16396 7064 16448
rect 7656 16396 7708 16448
rect 8760 16396 8812 16448
rect 9036 16396 9088 16448
rect 9312 16396 9364 16448
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 12624 16396 12676 16448
rect 13912 16396 13964 16448
rect 15108 16396 15160 16448
rect 17592 16396 17644 16448
rect 17776 16396 17828 16448
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 2136 16192 2188 16244
rect 3332 16192 3384 16244
rect 3700 16192 3752 16244
rect 112 16124 164 16176
rect 3608 16124 3660 16176
rect 4160 16124 4212 16176
rect 4436 16235 4488 16244
rect 4436 16201 4445 16235
rect 4445 16201 4479 16235
rect 4479 16201 4488 16235
rect 4436 16192 4488 16201
rect 4528 16192 4580 16244
rect 6000 16192 6052 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 6828 16124 6880 16176
rect 8392 16124 8444 16176
rect 8760 16124 8812 16176
rect 112 15988 164 16040
rect 1768 15988 1820 16040
rect 8208 16056 8260 16108
rect 4620 15988 4672 16040
rect 6092 15988 6144 16040
rect 2780 15963 2832 15972
rect 2780 15929 2789 15963
rect 2789 15929 2823 15963
rect 2823 15929 2832 15963
rect 2780 15920 2832 15929
rect 3332 15963 3384 15972
rect 3332 15929 3341 15963
rect 3341 15929 3375 15963
rect 3375 15929 3384 15963
rect 3332 15920 3384 15929
rect 4160 15963 4212 15972
rect 4160 15929 4169 15963
rect 4169 15929 4203 15963
rect 4203 15929 4212 15963
rect 4160 15920 4212 15929
rect 3700 15852 3752 15904
rect 5080 15852 5132 15904
rect 6368 15920 6420 15972
rect 6092 15852 6144 15904
rect 6920 15852 6972 15904
rect 7012 15852 7064 15904
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 8116 15920 8168 15972
rect 7840 15852 7892 15904
rect 8392 15852 8444 15904
rect 9128 15920 9180 15972
rect 9956 16124 10008 16176
rect 10784 16192 10836 16244
rect 11244 16192 11296 16244
rect 10692 16124 10744 16176
rect 11612 16124 11664 16176
rect 9496 16056 9548 16108
rect 9864 16056 9916 16108
rect 11428 16099 11480 16108
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 10508 15988 10560 16040
rect 11152 15988 11204 16040
rect 12072 16056 12124 16108
rect 12992 16056 13044 16108
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 15568 16192 15620 16244
rect 16028 16192 16080 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 17500 16192 17552 16244
rect 18696 16192 18748 16244
rect 20260 16192 20312 16244
rect 15476 16124 15528 16176
rect 18972 16124 19024 16176
rect 19156 16124 19208 16176
rect 16948 16056 17000 16108
rect 17684 16056 17736 16108
rect 15108 15988 15160 16040
rect 15936 15988 15988 16040
rect 11520 15920 11572 15972
rect 10692 15852 10744 15904
rect 11060 15852 11112 15904
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 12808 15852 12860 15904
rect 13176 15852 13228 15904
rect 15568 15920 15620 15972
rect 16672 15988 16724 16040
rect 18696 15988 18748 16040
rect 20720 16056 20772 16108
rect 19800 15988 19852 16040
rect 16396 15920 16448 15972
rect 18236 15920 18288 15972
rect 18972 15920 19024 15972
rect 19340 15920 19392 15972
rect 21640 15988 21692 16040
rect 19708 15852 19760 15904
rect 20812 15852 20864 15904
rect 21456 15852 21508 15904
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 1768 15648 1820 15700
rect 2780 15648 2832 15700
rect 4620 15691 4672 15700
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 2596 15580 2648 15632
rect 2964 15623 3016 15632
rect 2964 15589 2973 15623
rect 2973 15589 3007 15623
rect 3007 15589 3016 15623
rect 2964 15580 3016 15589
rect 4620 15657 4629 15691
rect 4629 15657 4663 15691
rect 4663 15657 4672 15691
rect 4620 15648 4672 15657
rect 5356 15691 5408 15700
rect 5356 15657 5365 15691
rect 5365 15657 5399 15691
rect 5399 15657 5408 15691
rect 5356 15648 5408 15657
rect 9956 15648 10008 15700
rect 13452 15648 13504 15700
rect 16028 15648 16080 15700
rect 1124 15512 1176 15564
rect 1768 15512 1820 15564
rect 3516 15512 3568 15564
rect 4252 15512 4304 15564
rect 4896 15580 4948 15632
rect 5172 15580 5224 15632
rect 6000 15580 6052 15632
rect 6644 15580 6696 15632
rect 8392 15580 8444 15632
rect 8484 15580 8536 15632
rect 8760 15580 8812 15632
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 10968 15580 11020 15632
rect 11152 15580 11204 15632
rect 12624 15580 12676 15632
rect 6184 15512 6236 15564
rect 13176 15580 13228 15632
rect 14832 15580 14884 15632
rect 18144 15648 18196 15700
rect 19432 15691 19484 15700
rect 19432 15657 19441 15691
rect 19441 15657 19475 15691
rect 19475 15657 19484 15691
rect 19432 15648 19484 15657
rect 12900 15512 12952 15564
rect 14648 15512 14700 15564
rect 15108 15512 15160 15564
rect 15568 15512 15620 15564
rect 17040 15512 17092 15564
rect 19984 15580 20036 15632
rect 17500 15512 17552 15564
rect 1400 15444 1452 15496
rect 2320 15444 2372 15496
rect 2964 15444 3016 15496
rect 3884 15444 3936 15496
rect 4160 15444 4212 15496
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 4988 15444 5040 15496
rect 6552 15444 6604 15496
rect 6644 15444 6696 15496
rect 7840 15444 7892 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 11428 15444 11480 15496
rect 756 15376 808 15428
rect 1124 15376 1176 15428
rect 3056 15376 3108 15428
rect 6276 15376 6328 15428
rect 3240 15308 3292 15360
rect 3700 15308 3752 15360
rect 3976 15308 4028 15360
rect 4160 15308 4212 15360
rect 5356 15308 5408 15360
rect 6552 15308 6604 15360
rect 10048 15376 10100 15428
rect 10324 15419 10376 15428
rect 10324 15385 10333 15419
rect 10333 15385 10367 15419
rect 10367 15385 10376 15419
rect 10324 15376 10376 15385
rect 12072 15444 12124 15496
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 15660 15444 15712 15496
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 17684 15444 17736 15496
rect 18236 15512 18288 15564
rect 18880 15512 18932 15564
rect 19156 15512 19208 15564
rect 20168 15512 20220 15564
rect 20812 15512 20864 15564
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19064 15444 19116 15453
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 8116 15308 8168 15360
rect 9680 15308 9732 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 11152 15308 11204 15360
rect 18144 15376 18196 15428
rect 12808 15308 12860 15360
rect 15568 15308 15620 15360
rect 15936 15308 15988 15360
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 16856 15308 16908 15360
rect 17684 15308 17736 15360
rect 17776 15308 17828 15360
rect 19432 15308 19484 15360
rect 20168 15351 20220 15360
rect 20168 15317 20177 15351
rect 20177 15317 20211 15351
rect 20211 15317 20220 15351
rect 20168 15308 20220 15317
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 2872 15104 2924 15156
rect 3792 15104 3844 15156
rect 3976 15104 4028 15156
rect 4252 15104 4304 15156
rect 6184 15104 6236 15156
rect 6460 15104 6512 15156
rect 1584 15079 1636 15088
rect 1584 15045 1593 15079
rect 1593 15045 1627 15079
rect 1627 15045 1636 15079
rect 1584 15036 1636 15045
rect 2044 15036 2096 15088
rect 2228 14968 2280 15020
rect 3148 14968 3200 15020
rect 3792 14968 3844 15020
rect 296 14900 348 14952
rect 2044 14900 2096 14952
rect 5172 15036 5224 15088
rect 6828 15036 6880 15088
rect 8392 15079 8444 15088
rect 8392 15045 8401 15079
rect 8401 15045 8435 15079
rect 8435 15045 8444 15079
rect 8392 15036 8444 15045
rect 7840 14968 7892 15020
rect 6276 14900 6328 14952
rect 1216 14832 1268 14884
rect 5080 14832 5132 14884
rect 5264 14832 5316 14884
rect 6552 14832 6604 14884
rect 2596 14764 2648 14816
rect 4436 14764 4488 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 6000 14764 6052 14816
rect 6828 14764 6880 14816
rect 7840 14832 7892 14884
rect 8576 15036 8628 15088
rect 9128 15036 9180 15088
rect 10508 15104 10560 15156
rect 11244 15147 11296 15156
rect 11244 15113 11253 15147
rect 11253 15113 11287 15147
rect 11287 15113 11296 15147
rect 11244 15104 11296 15113
rect 9772 15036 9824 15088
rect 15568 15104 15620 15156
rect 16212 15104 16264 15156
rect 16948 15104 17000 15156
rect 17500 15104 17552 15156
rect 20812 15104 20864 15156
rect 21732 15147 21784 15156
rect 21732 15113 21741 15147
rect 21741 15113 21775 15147
rect 21775 15113 21784 15147
rect 21732 15104 21784 15113
rect 10324 14968 10376 15020
rect 12808 14968 12860 15020
rect 20628 15036 20680 15088
rect 11244 14900 11296 14952
rect 12164 14900 12216 14952
rect 15108 14900 15160 14952
rect 15844 14900 15896 14952
rect 16212 14943 16264 14952
rect 8760 14875 8812 14884
rect 8760 14841 8769 14875
rect 8769 14841 8803 14875
rect 8803 14841 8812 14875
rect 8760 14832 8812 14841
rect 9128 14832 9180 14884
rect 9864 14832 9916 14884
rect 9956 14764 10008 14816
rect 10324 14875 10376 14884
rect 10324 14841 10333 14875
rect 10333 14841 10367 14875
rect 10367 14841 10376 14875
rect 10324 14832 10376 14841
rect 10968 14832 11020 14884
rect 14188 14832 14240 14884
rect 11152 14764 11204 14816
rect 11428 14764 11480 14816
rect 14004 14764 14056 14816
rect 15016 14832 15068 14884
rect 16212 14909 16221 14943
rect 16221 14909 16255 14943
rect 16255 14909 16264 14943
rect 16212 14900 16264 14909
rect 17500 14900 17552 14952
rect 18880 14900 18932 14952
rect 19524 14900 19576 14952
rect 19984 14900 20036 14952
rect 21732 14900 21784 14952
rect 18144 14875 18196 14884
rect 15844 14764 15896 14816
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 18144 14841 18153 14875
rect 18153 14841 18187 14875
rect 18187 14841 18196 14875
rect 18144 14832 18196 14841
rect 18236 14875 18288 14884
rect 18236 14841 18245 14875
rect 18245 14841 18279 14875
rect 18279 14841 18288 14875
rect 18788 14875 18840 14884
rect 18236 14832 18288 14841
rect 18788 14841 18797 14875
rect 18797 14841 18831 14875
rect 18831 14841 18840 14875
rect 18788 14832 18840 14841
rect 296 14696 348 14748
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 572 14603 624 14612
rect 572 14569 581 14603
rect 581 14569 615 14603
rect 615 14569 624 14603
rect 572 14560 624 14569
rect 1860 14560 1912 14612
rect 2044 14560 2096 14612
rect 3332 14560 3384 14612
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 4988 14560 5040 14612
rect 5172 14603 5224 14612
rect 5172 14569 5181 14603
rect 5181 14569 5215 14603
rect 5215 14569 5224 14603
rect 5172 14560 5224 14569
rect 5264 14560 5316 14612
rect 2596 14535 2648 14544
rect 2596 14501 2605 14535
rect 2605 14501 2639 14535
rect 2639 14501 2648 14535
rect 2596 14492 2648 14501
rect 2688 14492 2740 14544
rect 3516 14492 3568 14544
rect 572 14424 624 14476
rect 1308 14424 1360 14476
rect 3700 14424 3752 14476
rect 5448 14492 5500 14544
rect 6276 14560 6328 14612
rect 8208 14603 8260 14612
rect 8208 14569 8217 14603
rect 8217 14569 8251 14603
rect 8251 14569 8260 14603
rect 8208 14560 8260 14569
rect 8392 14492 8444 14544
rect 8760 14560 8812 14612
rect 8852 14560 8904 14612
rect 9864 14560 9916 14612
rect 10416 14560 10468 14612
rect 12808 14603 12860 14612
rect 12808 14569 12817 14603
rect 12817 14569 12851 14603
rect 12851 14569 12860 14603
rect 12808 14560 12860 14569
rect 13912 14560 13964 14612
rect 14188 14560 14240 14612
rect 15752 14560 15804 14612
rect 17316 14560 17368 14612
rect 18052 14560 18104 14612
rect 4712 14356 4764 14408
rect 5448 14356 5500 14408
rect 5908 14424 5960 14476
rect 8576 14424 8628 14476
rect 10324 14492 10376 14544
rect 14740 14535 14792 14544
rect 14740 14501 14749 14535
rect 14749 14501 14783 14535
rect 14783 14501 14792 14535
rect 14740 14492 14792 14501
rect 16028 14492 16080 14544
rect 16488 14492 16540 14544
rect 16856 14492 16908 14544
rect 18512 14535 18564 14544
rect 18512 14501 18521 14535
rect 18521 14501 18555 14535
rect 18555 14501 18564 14535
rect 18512 14492 18564 14501
rect 19432 14492 19484 14544
rect 19984 14492 20036 14544
rect 20260 14492 20312 14544
rect 20720 14492 20772 14544
rect 9128 14424 9180 14476
rect 9588 14424 9640 14476
rect 13360 14424 13412 14476
rect 13636 14424 13688 14476
rect 14556 14424 14608 14476
rect 15568 14424 15620 14476
rect 15752 14424 15804 14476
rect 16580 14424 16632 14476
rect 20812 14424 20864 14476
rect 7656 14356 7708 14408
rect 7932 14356 7984 14408
rect 8208 14356 8260 14408
rect 8392 14356 8444 14408
rect 9956 14356 10008 14408
rect 10784 14356 10836 14408
rect 12256 14356 12308 14408
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 1952 14331 2004 14340
rect 1952 14297 1961 14331
rect 1961 14297 1995 14331
rect 1995 14297 2004 14331
rect 1952 14288 2004 14297
rect 2412 14288 2464 14340
rect 2688 14288 2740 14340
rect 3700 14288 3752 14340
rect 3884 14331 3936 14340
rect 3884 14297 3893 14331
rect 3893 14297 3927 14331
rect 3927 14297 3936 14331
rect 3884 14288 3936 14297
rect 4804 14288 4856 14340
rect 5908 14288 5960 14340
rect 9588 14288 9640 14340
rect 9864 14288 9916 14340
rect 15476 14288 15528 14340
rect 15936 14288 15988 14340
rect 1860 14220 1912 14272
rect 4436 14220 4488 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 6368 14220 6420 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 6828 14263 6880 14272
rect 6828 14229 6837 14263
rect 6837 14229 6871 14263
rect 6871 14229 6880 14263
rect 6828 14220 6880 14229
rect 7932 14220 7984 14272
rect 9220 14220 9272 14272
rect 10692 14220 10744 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 12164 14220 12216 14272
rect 14740 14220 14792 14272
rect 16488 14220 16540 14272
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17776 14356 17828 14408
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 19800 14356 19852 14408
rect 16948 14288 17000 14340
rect 20444 14288 20496 14340
rect 18236 14220 18288 14272
rect 21272 14288 21324 14340
rect 21364 14220 21416 14272
rect 22008 14263 22060 14272
rect 22008 14229 22017 14263
rect 22017 14229 22051 14263
rect 22051 14229 22060 14263
rect 22008 14220 22060 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 1308 14016 1360 14068
rect 2228 14016 2280 14068
rect 2504 14016 2556 14068
rect 3148 14016 3200 14068
rect 7012 14016 7064 14068
rect 8760 14016 8812 14068
rect 9312 14016 9364 14068
rect 10600 14016 10652 14068
rect 11336 14016 11388 14068
rect 11612 14016 11664 14068
rect 12440 14016 12492 14068
rect 14188 14016 14240 14068
rect 14556 14016 14608 14068
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 15292 14016 15344 14068
rect 18236 14016 18288 14068
rect 19156 14059 19208 14068
rect 19156 14025 19165 14059
rect 19165 14025 19199 14059
rect 19199 14025 19208 14059
rect 19156 14016 19208 14025
rect 2320 13948 2372 14000
rect 3516 13948 3568 14000
rect 4436 13991 4488 14000
rect 1124 13880 1176 13932
rect 1308 13880 1360 13932
rect 2136 13880 2188 13932
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 4804 13948 4856 14000
rect 4620 13880 4672 13932
rect 2780 13812 2832 13864
rect 4896 13812 4948 13864
rect 5724 13948 5776 14000
rect 6184 13948 6236 14000
rect 5448 13880 5500 13932
rect 1124 13676 1176 13728
rect 2044 13676 2096 13728
rect 3516 13676 3568 13728
rect 3700 13719 3752 13728
rect 3700 13685 3709 13719
rect 3709 13685 3743 13719
rect 3743 13685 3752 13719
rect 3700 13676 3752 13685
rect 5080 13744 5132 13796
rect 5724 13744 5776 13796
rect 6276 13744 6328 13796
rect 7564 13880 7616 13932
rect 7012 13744 7064 13796
rect 7564 13744 7616 13796
rect 7840 13880 7892 13932
rect 8576 13948 8628 14000
rect 8944 13948 8996 14000
rect 9680 13948 9732 14000
rect 10416 13880 10468 13932
rect 16764 13948 16816 14000
rect 17408 13948 17460 14000
rect 18696 13948 18748 14000
rect 20812 14016 20864 14068
rect 15108 13880 15160 13932
rect 16948 13880 17000 13932
rect 17316 13880 17368 13932
rect 9128 13812 9180 13864
rect 11888 13812 11940 13864
rect 12900 13812 12952 13864
rect 14188 13812 14240 13864
rect 14832 13812 14884 13864
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 16580 13812 16632 13864
rect 17868 13812 17920 13864
rect 19800 13855 19852 13864
rect 19800 13821 19809 13855
rect 19809 13821 19843 13855
rect 19843 13821 19852 13855
rect 19800 13812 19852 13821
rect 20996 13880 21048 13932
rect 23480 14016 23532 14068
rect 23572 13948 23624 14000
rect 21364 13812 21416 13864
rect 5448 13676 5500 13728
rect 6460 13719 6512 13728
rect 6460 13685 6469 13719
rect 6469 13685 6503 13719
rect 6503 13685 6512 13719
rect 6460 13676 6512 13685
rect 7380 13676 7432 13728
rect 7656 13676 7708 13728
rect 8852 13744 8904 13796
rect 9404 13744 9456 13796
rect 10692 13744 10744 13796
rect 8208 13676 8260 13728
rect 8484 13676 8536 13728
rect 9680 13676 9732 13728
rect 10416 13676 10468 13728
rect 12808 13676 12860 13728
rect 13176 13676 13228 13728
rect 15568 13744 15620 13796
rect 14740 13676 14792 13728
rect 15476 13676 15528 13728
rect 16856 13676 16908 13728
rect 17868 13676 17920 13728
rect 18236 13787 18288 13796
rect 18236 13753 18245 13787
rect 18245 13753 18279 13787
rect 18279 13753 18288 13787
rect 18236 13744 18288 13753
rect 18328 13676 18380 13728
rect 19340 13676 19392 13728
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 1124 13472 1176 13524
rect 2596 13472 2648 13524
rect 2504 13404 2556 13456
rect 3700 13404 3752 13456
rect 3884 13404 3936 13456
rect 4896 13404 4948 13456
rect 6000 13472 6052 13524
rect 5632 13404 5684 13456
rect 8392 13472 8444 13524
rect 10784 13472 10836 13524
rect 11060 13472 11112 13524
rect 8760 13404 8812 13456
rect 10416 13404 10468 13456
rect 11888 13404 11940 13456
rect 11980 13404 12032 13456
rect 12256 13472 12308 13524
rect 15936 13472 15988 13524
rect 18052 13472 18104 13524
rect 1492 13336 1544 13388
rect 1584 13336 1636 13388
rect 1860 13336 1912 13388
rect 4344 13336 4396 13388
rect 4436 13336 4488 13388
rect 7012 13379 7064 13388
rect 7012 13345 7030 13379
rect 7030 13345 7064 13379
rect 7012 13336 7064 13345
rect 7380 13336 7432 13388
rect 12348 13404 12400 13456
rect 13176 13404 13228 13456
rect 16672 13447 16724 13456
rect 16672 13413 16681 13447
rect 16681 13413 16715 13447
rect 16715 13413 16724 13447
rect 16672 13404 16724 13413
rect 18236 13447 18288 13456
rect 18236 13413 18245 13447
rect 18245 13413 18279 13447
rect 18279 13413 18288 13447
rect 18236 13404 18288 13413
rect 18512 13472 18564 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 20904 13472 20956 13524
rect 12440 13336 12492 13388
rect 13912 13336 13964 13388
rect 14372 13336 14424 13388
rect 2320 13268 2372 13320
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 388 13200 440 13252
rect 1124 13200 1176 13252
rect 2044 13200 2096 13252
rect 2504 13200 2556 13252
rect 6460 13268 6512 13320
rect 9588 13268 9640 13320
rect 9956 13268 10008 13320
rect 12164 13268 12216 13320
rect 12256 13268 12308 13320
rect 13268 13268 13320 13320
rect 4620 13200 4672 13252
rect 4988 13200 5040 13252
rect 8576 13243 8628 13252
rect 8576 13209 8585 13243
rect 8585 13209 8619 13243
rect 8619 13209 8628 13243
rect 8576 13200 8628 13209
rect 12072 13243 12124 13252
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 2320 13132 2372 13184
rect 3332 13132 3384 13184
rect 3608 13132 3660 13184
rect 4436 13132 4488 13184
rect 4712 13132 4764 13184
rect 7656 13132 7708 13184
rect 8024 13132 8076 13184
rect 8392 13132 8444 13184
rect 8852 13132 8904 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 11244 13175 11296 13184
rect 11244 13141 11253 13175
rect 11253 13141 11287 13175
rect 11287 13141 11296 13175
rect 11244 13132 11296 13141
rect 12072 13209 12081 13243
rect 12081 13209 12115 13243
rect 12115 13209 12124 13243
rect 12072 13200 12124 13209
rect 12440 13200 12492 13252
rect 15568 13336 15620 13388
rect 18880 13336 18932 13388
rect 19432 13336 19484 13388
rect 20812 13336 20864 13388
rect 20996 13336 21048 13388
rect 22100 13336 22152 13388
rect 17316 13268 17368 13320
rect 18512 13268 18564 13320
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 14556 13175 14608 13184
rect 14556 13141 14565 13175
rect 14565 13141 14599 13175
rect 14599 13141 14608 13175
rect 14556 13132 14608 13141
rect 14648 13132 14700 13184
rect 15200 13132 15252 13184
rect 15292 13132 15344 13184
rect 18328 13200 18380 13252
rect 22560 13200 22612 13252
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 16580 13132 16632 13184
rect 16856 13132 16908 13184
rect 17776 13132 17828 13184
rect 18420 13132 18472 13184
rect 21916 13175 21968 13184
rect 21916 13141 21925 13175
rect 21925 13141 21959 13175
rect 21959 13141 21968 13175
rect 21916 13132 21968 13141
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 1584 12928 1636 12980
rect 1768 12928 1820 12980
rect 4436 12928 4488 12980
rect 5816 12928 5868 12980
rect 6828 12928 6880 12980
rect 8760 12928 8812 12980
rect 9220 12928 9272 12980
rect 9588 12928 9640 12980
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 2964 12860 3016 12912
rect 3424 12903 3476 12912
rect 3424 12869 3433 12903
rect 3433 12869 3467 12903
rect 3467 12869 3476 12903
rect 3424 12860 3476 12869
rect 3884 12860 3936 12912
rect 5448 12860 5500 12912
rect 7012 12860 7064 12912
rect 7656 12860 7708 12912
rect 9312 12860 9364 12912
rect 10508 12860 10560 12912
rect 12072 12928 12124 12980
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 13912 12928 13964 12980
rect 14096 12928 14148 12980
rect 16948 12928 17000 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20812 12928 20864 12980
rect 21548 12928 21600 12980
rect 22100 12971 22152 12980
rect 22100 12937 22109 12971
rect 22109 12937 22143 12971
rect 22143 12937 22152 12971
rect 22100 12928 22152 12937
rect 11704 12860 11756 12912
rect 11980 12860 12032 12912
rect 14372 12860 14424 12912
rect 18236 12860 18288 12912
rect 20 12792 72 12844
rect 1768 12792 1820 12844
rect 3148 12792 3200 12844
rect 3240 12792 3292 12844
rect 3516 12792 3568 12844
rect 5632 12792 5684 12844
rect 6552 12792 6604 12844
rect 7380 12792 7432 12844
rect 9404 12792 9456 12844
rect 9864 12792 9916 12844
rect 3332 12724 3384 12776
rect 3884 12724 3936 12776
rect 1952 12656 2004 12708
rect 1676 12588 1728 12640
rect 3148 12699 3200 12708
rect 3148 12665 3157 12699
rect 3157 12665 3191 12699
rect 3191 12665 3200 12699
rect 3148 12656 3200 12665
rect 3240 12656 3292 12708
rect 4344 12724 4396 12776
rect 3976 12588 4028 12640
rect 4804 12656 4856 12708
rect 4896 12699 4948 12708
rect 4896 12665 4905 12699
rect 4905 12665 4939 12699
rect 4939 12665 4948 12699
rect 4896 12656 4948 12665
rect 5724 12656 5776 12708
rect 6828 12656 6880 12708
rect 7748 12656 7800 12708
rect 8208 12656 8260 12708
rect 5632 12588 5684 12640
rect 6000 12588 6052 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 7380 12588 7432 12640
rect 8576 12588 8628 12640
rect 9312 12656 9364 12708
rect 13636 12792 13688 12844
rect 16764 12792 16816 12844
rect 21456 12860 21508 12912
rect 22652 12860 22704 12912
rect 18788 12835 18840 12844
rect 10876 12699 10928 12708
rect 10876 12665 10885 12699
rect 10885 12665 10919 12699
rect 10919 12665 10928 12699
rect 10876 12656 10928 12665
rect 10416 12588 10468 12640
rect 10600 12588 10652 12640
rect 11428 12588 11480 12640
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14096 12724 14148 12776
rect 14372 12724 14424 12776
rect 15292 12724 15344 12776
rect 15568 12724 15620 12776
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 20168 12767 20220 12776
rect 14924 12656 14976 12708
rect 16028 12699 16080 12708
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 12348 12588 12400 12640
rect 14096 12588 14148 12640
rect 16028 12665 16031 12699
rect 16031 12665 16065 12699
rect 16065 12665 16080 12699
rect 16028 12656 16080 12665
rect 17868 12656 17920 12708
rect 16580 12588 16632 12640
rect 16672 12588 16724 12640
rect 19248 12656 19300 12708
rect 20168 12733 20177 12767
rect 20177 12733 20211 12767
rect 20211 12733 20220 12767
rect 20168 12724 20220 12733
rect 20536 12724 20588 12776
rect 20720 12656 20772 12708
rect 18696 12588 18748 12640
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 2136 12384 2188 12436
rect 3240 12384 3292 12436
rect 6460 12384 6512 12436
rect 8024 12384 8076 12436
rect 2872 12316 2924 12368
rect 4160 12316 4212 12368
rect 6000 12316 6052 12368
rect 6276 12359 6328 12368
rect 6276 12325 6285 12359
rect 6285 12325 6319 12359
rect 6319 12325 6328 12359
rect 6276 12316 6328 12325
rect 7012 12316 7064 12368
rect 7748 12316 7800 12368
rect 8576 12384 8628 12436
rect 11704 12427 11756 12436
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 9864 12316 9916 12368
rect 13452 12427 13504 12436
rect 1400 12248 1452 12300
rect 2412 12248 2464 12300
rect 3148 12248 3200 12300
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 4344 12180 4396 12232
rect 2412 12112 2464 12164
rect 2136 12044 2188 12096
rect 3240 12044 3292 12096
rect 3884 12044 3936 12096
rect 4252 12044 4304 12096
rect 4528 12044 4580 12096
rect 4896 12180 4948 12232
rect 5540 12180 5592 12232
rect 5724 12180 5776 12232
rect 7472 12248 7524 12300
rect 8944 12248 8996 12300
rect 6276 12180 6328 12232
rect 6920 12180 6972 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 8392 12180 8444 12232
rect 9036 12180 9088 12232
rect 11060 12248 11112 12300
rect 11704 12248 11756 12300
rect 12348 12248 12400 12300
rect 12992 12316 13044 12368
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 13912 12384 13964 12436
rect 16120 12384 16172 12436
rect 18144 12384 18196 12436
rect 18328 12384 18380 12436
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 20444 12384 20496 12436
rect 15016 12316 15068 12368
rect 10048 12180 10100 12232
rect 10876 12180 10928 12232
rect 13728 12248 13780 12300
rect 15568 12316 15620 12368
rect 16764 12316 16816 12368
rect 17500 12316 17552 12368
rect 15936 12248 15988 12300
rect 17224 12248 17276 12300
rect 17776 12248 17828 12300
rect 19432 12248 19484 12300
rect 19800 12248 19852 12300
rect 20812 12248 20864 12300
rect 21456 12248 21508 12300
rect 4804 12112 4856 12164
rect 5540 12087 5592 12096
rect 5540 12053 5549 12087
rect 5549 12053 5583 12087
rect 5583 12053 5592 12087
rect 5540 12044 5592 12053
rect 6736 12044 6788 12096
rect 11336 12112 11388 12164
rect 17408 12180 17460 12232
rect 17592 12180 17644 12232
rect 13636 12112 13688 12164
rect 13912 12112 13964 12164
rect 18512 12112 18564 12164
rect 7748 12044 7800 12096
rect 9312 12044 9364 12096
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 10692 12044 10744 12096
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 11152 12044 11204 12096
rect 14648 12044 14700 12096
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 17868 12087 17920 12096
rect 17868 12053 17877 12087
rect 17877 12053 17911 12087
rect 17911 12053 17920 12087
rect 17868 12044 17920 12053
rect 19524 12044 19576 12096
rect 21640 12044 21692 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 3976 11840 4028 11892
rect 4160 11840 4212 11892
rect 6276 11840 6328 11892
rect 6920 11840 6972 11892
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 11888 11840 11940 11892
rect 20 11772 72 11824
rect 6368 11772 6420 11824
rect 7932 11772 7984 11824
rect 12348 11772 12400 11824
rect 14188 11840 14240 11892
rect 16488 11840 16540 11892
rect 17500 11840 17552 11892
rect 18236 11840 18288 11892
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 19616 11840 19668 11892
rect 204 11704 256 11756
rect 2596 11704 2648 11756
rect 4528 11704 4580 11756
rect 940 11568 992 11620
rect 1400 11568 1452 11620
rect 3608 11636 3660 11688
rect 4344 11636 4396 11688
rect 6460 11704 6512 11756
rect 5448 11636 5500 11688
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 2872 11543 2924 11552
rect 1768 11500 1820 11509
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 3608 11500 3660 11552
rect 3884 11500 3936 11552
rect 4068 11568 4120 11620
rect 4896 11611 4948 11620
rect 4896 11577 4905 11611
rect 4905 11577 4939 11611
rect 4939 11577 4948 11611
rect 4896 11568 4948 11577
rect 6736 11704 6788 11756
rect 8852 11704 8904 11756
rect 9772 11704 9824 11756
rect 10416 11636 10468 11688
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 12808 11704 12860 11756
rect 13452 11704 13504 11756
rect 4804 11500 4856 11552
rect 5908 11500 5960 11552
rect 6276 11500 6328 11552
rect 8484 11500 8536 11552
rect 10324 11568 10376 11620
rect 11888 11636 11940 11688
rect 14832 11704 14884 11756
rect 15568 11704 15620 11756
rect 16120 11704 16172 11756
rect 19800 11772 19852 11824
rect 18420 11704 18472 11756
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 20168 11704 20220 11756
rect 20812 11840 20864 11892
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 21732 11840 21784 11892
rect 21456 11772 21508 11824
rect 21364 11704 21416 11756
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 21732 11636 21784 11688
rect 13084 11568 13136 11620
rect 14096 11568 14148 11620
rect 16120 11568 16172 11620
rect 17592 11568 17644 11620
rect 18144 11611 18196 11620
rect 18144 11577 18153 11611
rect 18153 11577 18187 11611
rect 18187 11577 18196 11611
rect 18144 11568 18196 11577
rect 18236 11611 18288 11620
rect 18236 11577 18245 11611
rect 18245 11577 18279 11611
rect 18279 11577 18288 11611
rect 18236 11568 18288 11577
rect 19800 11611 19852 11620
rect 19800 11577 19809 11611
rect 19809 11577 19843 11611
rect 19843 11577 19852 11611
rect 19800 11568 19852 11577
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 12440 11500 12492 11552
rect 13636 11500 13688 11552
rect 14648 11500 14700 11552
rect 15016 11500 15068 11552
rect 18604 11500 18656 11552
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 848 11296 900 11348
rect 1768 11228 1820 11280
rect 204 11160 256 11212
rect 3516 11296 3568 11348
rect 3884 11296 3936 11348
rect 4344 11296 4396 11348
rect 4896 11296 4948 11348
rect 4068 11228 4120 11280
rect 7196 11296 7248 11348
rect 7748 11296 7800 11348
rect 8576 11296 8628 11348
rect 9312 11296 9364 11348
rect 9864 11339 9916 11348
rect 9864 11305 9873 11339
rect 9873 11305 9907 11339
rect 9907 11305 9916 11339
rect 9864 11296 9916 11305
rect 10876 11296 10928 11348
rect 11980 11339 12032 11348
rect 5908 11228 5960 11280
rect 6552 11228 6604 11280
rect 4344 11160 4396 11212
rect 4252 11092 4304 11144
rect 5264 11160 5316 11212
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 9036 11228 9088 11280
rect 9220 11228 9272 11280
rect 11980 11305 11989 11339
rect 11989 11305 12023 11339
rect 12023 11305 12032 11339
rect 11980 11296 12032 11305
rect 12072 11296 12124 11348
rect 13084 11296 13136 11348
rect 13452 11296 13504 11348
rect 13728 11296 13780 11348
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 17868 11296 17920 11348
rect 19800 11296 19852 11348
rect 20168 11296 20220 11348
rect 20628 11296 20680 11348
rect 8852 11160 8904 11212
rect 10416 11160 10468 11212
rect 7748 11092 7800 11144
rect 11060 11228 11112 11280
rect 12624 11271 12676 11280
rect 12624 11237 12633 11271
rect 12633 11237 12667 11271
rect 12667 11237 12676 11271
rect 12624 11228 12676 11237
rect 12808 11228 12860 11280
rect 12900 11228 12952 11280
rect 13360 11228 13412 11280
rect 17776 11228 17828 11280
rect 18880 11228 18932 11280
rect 19892 11228 19944 11280
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 17592 11160 17644 11212
rect 20812 11160 20864 11212
rect 21732 11160 21784 11212
rect 4528 11067 4580 11076
rect 4528 11033 4537 11067
rect 4537 11033 4571 11067
rect 4571 11033 4580 11067
rect 4528 11024 4580 11033
rect 4804 11024 4856 11076
rect 5264 11067 5316 11076
rect 5264 11033 5273 11067
rect 5273 11033 5307 11067
rect 5307 11033 5316 11067
rect 5264 11024 5316 11033
rect 6736 11024 6788 11076
rect 7932 11024 7984 11076
rect 1768 10956 1820 11008
rect 3700 10956 3752 11008
rect 5724 10956 5776 11008
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 8116 10956 8168 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 9312 10956 9364 11008
rect 9496 10956 9548 11008
rect 10048 10956 10100 11008
rect 10876 11024 10928 11076
rect 13268 11092 13320 11144
rect 15292 11092 15344 11144
rect 15936 11092 15988 11144
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 11336 11024 11388 11076
rect 13176 11067 13228 11076
rect 13176 11033 13185 11067
rect 13185 11033 13219 11067
rect 13219 11033 13228 11067
rect 13176 11024 13228 11033
rect 13360 10956 13412 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 17316 10999 17368 11008
rect 17316 10965 17325 10999
rect 17325 10965 17359 10999
rect 17359 10965 17368 10999
rect 17316 10956 17368 10965
rect 18236 10956 18288 11008
rect 18604 10956 18656 11008
rect 20720 10956 20772 11008
rect 22284 10999 22336 11008
rect 22284 10965 22293 10999
rect 22293 10965 22327 10999
rect 22327 10965 22336 10999
rect 22284 10956 22336 10965
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 1216 10752 1268 10804
rect 2688 10752 2740 10804
rect 4160 10752 4212 10804
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 5908 10752 5960 10804
rect 7748 10752 7800 10804
rect 8760 10752 8812 10804
rect 9404 10752 9456 10804
rect 11060 10752 11112 10804
rect 11704 10752 11756 10804
rect 11980 10752 12032 10804
rect 13360 10752 13412 10804
rect 13912 10752 13964 10804
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 16120 10752 16172 10804
rect 17592 10795 17644 10804
rect 17592 10761 17601 10795
rect 17601 10761 17635 10795
rect 17635 10761 17644 10795
rect 17592 10752 17644 10761
rect 18328 10752 18380 10804
rect 18880 10752 18932 10804
rect 19616 10752 19668 10804
rect 20260 10752 20312 10804
rect 3976 10684 4028 10736
rect 9036 10684 9088 10736
rect 9496 10684 9548 10736
rect 10876 10684 10928 10736
rect 7564 10659 7616 10668
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2504 10412 2556 10464
rect 3884 10548 3936 10600
rect 4528 10548 4580 10600
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8116 10616 8168 10668
rect 9128 10616 9180 10668
rect 9772 10616 9824 10668
rect 5080 10548 5132 10600
rect 5448 10548 5500 10600
rect 8484 10548 8536 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10416 10616 10468 10668
rect 13452 10684 13504 10736
rect 17684 10684 17736 10736
rect 20444 10684 20496 10736
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 3884 10412 3936 10464
rect 4344 10412 4396 10464
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5448 10412 5500 10464
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 9772 10480 9824 10532
rect 12808 10616 12860 10668
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 16212 10616 16264 10668
rect 17960 10616 18012 10668
rect 15292 10548 15344 10600
rect 12532 10523 12584 10532
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 12900 10480 12952 10532
rect 13176 10523 13228 10532
rect 13176 10489 13185 10523
rect 13185 10489 13219 10523
rect 13219 10489 13228 10523
rect 13176 10480 13228 10489
rect 14648 10523 14700 10532
rect 14648 10489 14657 10523
rect 14657 10489 14691 10523
rect 14691 10489 14700 10523
rect 14648 10480 14700 10489
rect 16120 10480 16172 10532
rect 16580 10480 16632 10532
rect 18236 10523 18288 10532
rect 18236 10489 18245 10523
rect 18245 10489 18279 10523
rect 18279 10489 18288 10523
rect 18236 10480 18288 10489
rect 18788 10523 18840 10532
rect 18788 10489 18797 10523
rect 18797 10489 18831 10523
rect 18831 10489 18840 10523
rect 18788 10480 18840 10489
rect 7748 10412 7800 10464
rect 8484 10412 8536 10464
rect 10048 10412 10100 10464
rect 10876 10412 10928 10464
rect 11704 10412 11756 10464
rect 17776 10412 17828 10464
rect 20812 10752 20864 10804
rect 21732 10795 21784 10804
rect 21732 10761 21741 10795
rect 21741 10761 21775 10795
rect 21775 10761 21784 10795
rect 21732 10752 21784 10761
rect 23480 10684 23532 10736
rect 20536 10480 20588 10532
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 3700 10251 3752 10260
rect 3700 10217 3709 10251
rect 3709 10217 3743 10251
rect 3743 10217 3752 10251
rect 3700 10208 3752 10217
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 4620 10208 4672 10260
rect 4804 10208 4856 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 6092 10208 6144 10260
rect 6552 10208 6604 10260
rect 3516 10140 3568 10192
rect 4528 10140 4580 10192
rect 5172 10140 5224 10192
rect 7840 10208 7892 10260
rect 9956 10208 10008 10260
rect 10600 10208 10652 10260
rect 11520 10208 11572 10260
rect 12440 10208 12492 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 8576 10140 8628 10192
rect 9312 10140 9364 10192
rect 11152 10140 11204 10192
rect 13176 10208 13228 10260
rect 13452 10208 13504 10260
rect 14648 10208 14700 10260
rect 15752 10208 15804 10260
rect 16212 10208 16264 10260
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 16764 10208 16816 10260
rect 12808 10140 12860 10192
rect 13636 10140 13688 10192
rect 2780 10072 2832 10124
rect 4160 10072 4212 10124
rect 5816 10072 5868 10124
rect 6920 10072 6972 10124
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 8760 10072 8812 10124
rect 9680 10072 9732 10124
rect 572 9936 624 9988
rect 3884 10004 3936 10056
rect 5264 10004 5316 10056
rect 5448 10004 5500 10056
rect 8024 10004 8076 10056
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 10876 10072 10928 10124
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 13176 10072 13228 10124
rect 10416 10004 10468 10056
rect 12256 10004 12308 10056
rect 2780 9936 2832 9988
rect 4068 9936 4120 9988
rect 572 9732 624 9784
rect 572 9634 624 9686
rect 3516 9868 3568 9920
rect 5080 9936 5132 9988
rect 9772 9936 9824 9988
rect 13452 10004 13504 10056
rect 14096 10140 14148 10192
rect 14832 10140 14884 10192
rect 17408 10183 17460 10192
rect 14740 10072 14792 10124
rect 15936 10072 15988 10124
rect 16856 10072 16908 10124
rect 17408 10149 17417 10183
rect 17417 10149 17451 10183
rect 17451 10149 17460 10183
rect 17408 10140 17460 10149
rect 18052 10208 18104 10260
rect 20444 10251 20496 10260
rect 20444 10217 20453 10251
rect 20453 10217 20487 10251
rect 20487 10217 20496 10251
rect 20444 10208 20496 10217
rect 20536 10208 20588 10260
rect 17868 10140 17920 10192
rect 18788 10140 18840 10192
rect 19064 10140 19116 10192
rect 17592 10072 17644 10124
rect 17776 10115 17828 10124
rect 17776 10081 17794 10115
rect 17794 10081 17828 10115
rect 17776 10072 17828 10081
rect 19984 10072 20036 10124
rect 20812 10072 20864 10124
rect 21732 10072 21784 10124
rect 18788 10047 18840 10056
rect 18788 10013 18797 10047
rect 18797 10013 18831 10047
rect 18831 10013 18840 10047
rect 18788 10004 18840 10013
rect 12992 9936 13044 9988
rect 13636 9979 13688 9988
rect 13636 9945 13645 9979
rect 13645 9945 13679 9979
rect 13679 9945 13688 9979
rect 13636 9936 13688 9945
rect 16856 9936 16908 9988
rect 18696 9936 18748 9988
rect 18880 9936 18932 9988
rect 20168 9936 20220 9988
rect 5632 9868 5684 9920
rect 6460 9868 6512 9920
rect 6644 9868 6696 9920
rect 6736 9868 6788 9920
rect 7012 9868 7064 9920
rect 8024 9868 8076 9920
rect 8300 9911 8352 9920
rect 8300 9877 8309 9911
rect 8309 9877 8343 9911
rect 8343 9877 8352 9911
rect 8300 9868 8352 9877
rect 8484 9868 8536 9920
rect 9036 9868 9088 9920
rect 9864 9868 9916 9920
rect 10048 9868 10100 9920
rect 10692 9868 10744 9920
rect 12440 9868 12492 9920
rect 15108 9868 15160 9920
rect 15292 9868 15344 9920
rect 16764 9868 16816 9920
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 2320 9707 2372 9716
rect 2320 9673 2329 9707
rect 2329 9673 2363 9707
rect 2363 9673 2372 9707
rect 2320 9664 2372 9673
rect 3056 9664 3108 9716
rect 3700 9664 3752 9716
rect 4068 9664 4120 9716
rect 4436 9664 4488 9716
rect 4620 9664 4672 9716
rect 5724 9664 5776 9716
rect 6644 9664 6696 9716
rect 2504 9596 2556 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 1768 9528 1820 9580
rect 2044 9528 2096 9580
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 3424 9596 3476 9648
rect 4344 9596 4396 9648
rect 4712 9639 4764 9648
rect 4712 9605 4721 9639
rect 4721 9605 4755 9639
rect 4755 9605 4764 9639
rect 4712 9596 4764 9605
rect 5264 9596 5316 9648
rect 7104 9596 7156 9648
rect 7472 9639 7524 9648
rect 7472 9605 7481 9639
rect 7481 9605 7515 9639
rect 7515 9605 7524 9639
rect 7472 9596 7524 9605
rect 9036 9664 9088 9716
rect 9680 9707 9732 9716
rect 9680 9673 9689 9707
rect 9689 9673 9723 9707
rect 9723 9673 9732 9707
rect 9680 9664 9732 9673
rect 10508 9664 10560 9716
rect 12716 9664 12768 9716
rect 13728 9664 13780 9716
rect 13912 9664 13964 9716
rect 14648 9664 14700 9716
rect 16304 9664 16356 9716
rect 17132 9707 17184 9716
rect 17132 9673 17141 9707
rect 17141 9673 17175 9707
rect 17175 9673 17184 9707
rect 17132 9664 17184 9673
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 18144 9664 18196 9716
rect 20812 9664 20864 9716
rect 22008 9664 22060 9716
rect 4436 9528 4488 9580
rect 5632 9528 5684 9580
rect 8208 9528 8260 9580
rect 11888 9596 11940 9648
rect 12164 9596 12216 9648
rect 14740 9596 14792 9648
rect 20536 9596 20588 9648
rect 21732 9596 21784 9648
rect 11060 9571 11112 9580
rect 11060 9537 11069 9571
rect 11069 9537 11103 9571
rect 11103 9537 11112 9571
rect 11060 9528 11112 9537
rect 17316 9528 17368 9580
rect 17592 9528 17644 9580
rect 18604 9528 18656 9580
rect 19984 9528 20036 9580
rect 1492 9460 1544 9512
rect 5080 9460 5132 9512
rect 6092 9460 6144 9512
rect 6276 9460 6328 9512
rect 8024 9460 8076 9512
rect 8576 9460 8628 9512
rect 9680 9460 9732 9512
rect 2504 9324 2556 9376
rect 4068 9392 4120 9444
rect 4436 9435 4488 9444
rect 4436 9401 4445 9435
rect 4445 9401 4479 9435
rect 4479 9401 4488 9435
rect 4436 9392 4488 9401
rect 4804 9392 4856 9444
rect 6920 9435 6972 9444
rect 6276 9324 6328 9376
rect 6920 9401 6929 9435
rect 6929 9401 6963 9435
rect 6963 9401 6972 9435
rect 6920 9392 6972 9401
rect 7104 9392 7156 9444
rect 8300 9392 8352 9444
rect 8024 9324 8076 9376
rect 10600 9392 10652 9444
rect 14464 9460 14516 9512
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 16948 9460 17000 9512
rect 17868 9460 17920 9512
rect 15108 9392 15160 9444
rect 16304 9435 16356 9444
rect 16304 9401 16313 9435
rect 16313 9401 16347 9435
rect 16347 9401 16356 9435
rect 18144 9435 18196 9444
rect 16304 9392 16356 9401
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 18236 9435 18288 9444
rect 18236 9401 18245 9435
rect 18245 9401 18279 9435
rect 18279 9401 18288 9435
rect 18236 9392 18288 9401
rect 18420 9392 18472 9444
rect 18880 9392 18932 9444
rect 19800 9460 19852 9512
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 10508 9324 10560 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 17868 9324 17920 9376
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 20996 9392 21048 9444
rect 21548 9392 21600 9444
rect 22008 9392 22060 9444
rect 20260 9324 20312 9376
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 1308 9120 1360 9172
rect 1216 9052 1268 9104
rect 2044 9052 2096 9104
rect 2320 9052 2372 9104
rect 3240 9120 3292 9172
rect 4436 9120 4488 9172
rect 5448 9120 5500 9172
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 4896 9052 4948 9104
rect 4988 9095 5040 9104
rect 4988 9061 4997 9095
rect 4997 9061 5031 9095
rect 5031 9061 5040 9095
rect 4988 9052 5040 9061
rect 1584 8984 1636 9036
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 6184 9052 6236 9104
rect 5448 8984 5500 9036
rect 6000 8984 6052 9036
rect 112 8959 164 8968
rect 112 8925 121 8959
rect 121 8925 155 8959
rect 155 8925 164 8959
rect 112 8916 164 8925
rect 1032 8848 1084 8900
rect 1768 8848 1820 8900
rect 2320 8916 2372 8968
rect 3148 8916 3200 8968
rect 4988 8916 5040 8968
rect 6644 8916 6696 8968
rect 4804 8848 4856 8900
rect 6276 8891 6328 8900
rect 6276 8857 6285 8891
rect 6285 8857 6319 8891
rect 6319 8857 6328 8891
rect 6276 8848 6328 8857
rect 1400 8780 1452 8832
rect 2964 8780 3016 8832
rect 3240 8780 3292 8832
rect 4712 8780 4764 8832
rect 6644 8780 6696 8832
rect 6828 9052 6880 9104
rect 7564 9052 7616 9104
rect 8024 9120 8076 9172
rect 8668 9120 8720 9172
rect 10140 9120 10192 9172
rect 10324 9120 10376 9172
rect 10876 9120 10928 9172
rect 12716 9120 12768 9172
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8116 8984 8168 9036
rect 8760 8984 8812 9036
rect 6828 8916 6880 8968
rect 10232 8984 10284 9036
rect 11704 9052 11756 9104
rect 13360 9120 13412 9172
rect 13728 9120 13780 9172
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 14556 9120 14608 9172
rect 16304 9120 16356 9172
rect 17776 9120 17828 9172
rect 14832 9052 14884 9104
rect 16580 9052 16632 9104
rect 18052 9095 18104 9104
rect 18052 9061 18061 9095
rect 18061 9061 18095 9095
rect 18095 9061 18104 9095
rect 18052 9052 18104 9061
rect 19064 9120 19116 9172
rect 19248 9120 19300 9172
rect 21916 9120 21968 9172
rect 18604 9052 18656 9104
rect 19340 9052 19392 9104
rect 19616 9052 19668 9104
rect 20996 9095 21048 9104
rect 20996 9061 21005 9095
rect 21005 9061 21039 9095
rect 21039 9061 21048 9095
rect 20996 9052 21048 9061
rect 21088 9095 21140 9104
rect 21088 9061 21097 9095
rect 21097 9061 21131 9095
rect 21131 9061 21140 9095
rect 21088 9052 21140 9061
rect 13636 8984 13688 9036
rect 13912 8984 13964 9036
rect 9772 8916 9824 8968
rect 11980 8916 12032 8968
rect 12256 8916 12308 8968
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 13268 8916 13320 8968
rect 14280 8916 14332 8968
rect 14648 8916 14700 8968
rect 15108 8916 15160 8968
rect 16856 8984 16908 9036
rect 19064 8984 19116 9036
rect 19524 8984 19576 9036
rect 19800 8984 19852 9036
rect 7472 8891 7524 8900
rect 7472 8857 7481 8891
rect 7481 8857 7515 8891
rect 7515 8857 7524 8891
rect 7472 8848 7524 8857
rect 7748 8848 7800 8900
rect 13636 8848 13688 8900
rect 14464 8848 14516 8900
rect 17960 8916 18012 8968
rect 18696 8848 18748 8900
rect 19616 8916 19668 8968
rect 21640 8848 21692 8900
rect 9128 8780 9180 8832
rect 9864 8823 9916 8832
rect 9864 8789 9873 8823
rect 9873 8789 9907 8823
rect 9907 8789 9916 8823
rect 9864 8780 9916 8789
rect 10232 8780 10284 8832
rect 12164 8780 12216 8832
rect 13728 8823 13780 8832
rect 13728 8789 13737 8823
rect 13737 8789 13771 8823
rect 13771 8789 13780 8823
rect 13728 8780 13780 8789
rect 15016 8780 15068 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 17316 8823 17368 8832
rect 17316 8789 17325 8823
rect 17325 8789 17359 8823
rect 17359 8789 17368 8823
rect 17316 8780 17368 8789
rect 18328 8780 18380 8832
rect 19616 8823 19668 8832
rect 19616 8789 19625 8823
rect 19625 8789 19659 8823
rect 19659 8789 19668 8823
rect 19616 8780 19668 8789
rect 19892 8780 19944 8832
rect 20536 8780 20588 8832
rect 21916 8823 21968 8832
rect 21916 8789 21925 8823
rect 21925 8789 21959 8823
rect 21959 8789 21968 8823
rect 21916 8780 21968 8789
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 1400 8576 1452 8628
rect 1952 8576 2004 8628
rect 3240 8576 3292 8628
rect 3516 8576 3568 8628
rect 3792 8576 3844 8628
rect 112 8508 164 8560
rect 4712 8508 4764 8560
rect 8024 8576 8076 8628
rect 10692 8576 10744 8628
rect 10876 8576 10928 8628
rect 11520 8576 11572 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 13360 8576 13412 8628
rect 13636 8576 13688 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 15108 8619 15160 8628
rect 13820 8576 13872 8585
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 9864 8508 9916 8560
rect 11060 8551 11112 8560
rect 11060 8517 11069 8551
rect 11069 8517 11103 8551
rect 11103 8517 11112 8551
rect 11060 8508 11112 8517
rect 11796 8508 11848 8560
rect 3148 8440 3200 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 20 8304 72 8356
rect 2964 8372 3016 8424
rect 4252 8440 4304 8492
rect 4436 8440 4488 8492
rect 7380 8440 7432 8492
rect 8852 8440 8904 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 3516 8372 3568 8424
rect 940 8236 992 8288
rect 2412 8304 2464 8356
rect 2872 8347 2924 8356
rect 2872 8313 2881 8347
rect 2881 8313 2915 8347
rect 2915 8313 2924 8347
rect 2872 8304 2924 8313
rect 3240 8347 3292 8356
rect 3240 8313 3249 8347
rect 3249 8313 3283 8347
rect 3283 8313 3292 8347
rect 3240 8304 3292 8313
rect 4344 8372 4396 8424
rect 4160 8304 4212 8356
rect 4252 8304 4304 8356
rect 5080 8372 5132 8424
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 2964 8236 3016 8288
rect 3792 8236 3844 8288
rect 4712 8236 4764 8288
rect 5172 8236 5224 8288
rect 5632 8304 5684 8356
rect 8208 8304 8260 8356
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 8484 8347 8536 8356
rect 8484 8313 8493 8347
rect 8493 8313 8527 8347
rect 8527 8313 8536 8347
rect 8484 8304 8536 8313
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 7104 8236 7156 8288
rect 7380 8236 7432 8288
rect 9864 8304 9916 8356
rect 10508 8440 10560 8492
rect 11428 8440 11480 8492
rect 12716 8440 12768 8492
rect 13636 8440 13688 8492
rect 11520 8372 11572 8424
rect 12256 8372 12308 8424
rect 10508 8347 10560 8356
rect 10508 8313 10511 8347
rect 10511 8313 10545 8347
rect 10545 8313 10560 8347
rect 10508 8304 10560 8313
rect 13176 8347 13228 8356
rect 11428 8279 11480 8288
rect 11428 8245 11437 8279
rect 11437 8245 11471 8279
rect 11471 8245 11480 8279
rect 11428 8236 11480 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 13176 8313 13185 8347
rect 13185 8313 13219 8347
rect 13219 8313 13228 8347
rect 14556 8508 14608 8560
rect 15476 8576 15528 8628
rect 16580 8576 16632 8628
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 18788 8576 18840 8628
rect 18880 8576 18932 8628
rect 19800 8576 19852 8628
rect 20812 8576 20864 8628
rect 14280 8440 14332 8492
rect 19892 8508 19944 8560
rect 20996 8508 21048 8560
rect 21916 8576 21968 8628
rect 21548 8508 21600 8560
rect 14924 8372 14976 8424
rect 15476 8440 15528 8492
rect 17868 8440 17920 8492
rect 19248 8440 19300 8492
rect 20444 8440 20496 8492
rect 15936 8372 15988 8424
rect 17224 8372 17276 8424
rect 19064 8372 19116 8424
rect 21732 8415 21784 8424
rect 21732 8381 21741 8415
rect 21741 8381 21775 8415
rect 21775 8381 21784 8415
rect 21732 8372 21784 8381
rect 13176 8304 13228 8313
rect 12164 8236 12216 8245
rect 12716 8236 12768 8288
rect 17316 8304 17368 8356
rect 16028 8236 16080 8288
rect 17776 8279 17828 8288
rect 17776 8245 17785 8279
rect 17785 8245 17819 8279
rect 17819 8245 17828 8279
rect 17776 8236 17828 8245
rect 18420 8304 18472 8356
rect 19340 8236 19392 8288
rect 19800 8347 19852 8356
rect 19800 8313 19809 8347
rect 19809 8313 19843 8347
rect 19843 8313 19852 8347
rect 19800 8304 19852 8313
rect 22100 8304 22152 8356
rect 21272 8236 21324 8288
rect 22468 8279 22520 8288
rect 22468 8245 22477 8279
rect 22477 8245 22511 8279
rect 22511 8245 22520 8279
rect 22468 8236 22520 8245
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 6920 8032 6972 8084
rect 7288 8032 7340 8084
rect 8300 8032 8352 8084
rect 9404 8032 9456 8084
rect 10508 8032 10560 8084
rect 2136 7964 2188 8016
rect 2412 7964 2464 8016
rect 3056 8007 3108 8016
rect 3056 7973 3065 8007
rect 3065 7973 3099 8007
rect 3099 7973 3108 8007
rect 3056 7964 3108 7973
rect 4896 7964 4948 8016
rect 6552 8007 6604 8016
rect 4160 7896 4212 7948
rect 1952 7828 2004 7880
rect 664 7760 716 7812
rect 1400 7760 1452 7812
rect 3148 7828 3200 7880
rect 5356 7896 5408 7948
rect 6552 7973 6561 8007
rect 6561 7973 6595 8007
rect 6595 7973 6604 8007
rect 6552 7964 6604 7973
rect 7748 7964 7800 8016
rect 7840 7964 7892 8016
rect 11152 8032 11204 8084
rect 11060 8007 11112 8016
rect 2688 7803 2740 7812
rect 2688 7769 2697 7803
rect 2697 7769 2731 7803
rect 2731 7769 2740 7803
rect 2688 7760 2740 7769
rect 3240 7760 3292 7812
rect 6276 7828 6328 7880
rect 1492 7692 1544 7744
rect 2964 7692 3016 7744
rect 4436 7692 4488 7744
rect 6000 7760 6052 7812
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 7564 7896 7616 7948
rect 8116 7896 8168 7948
rect 8392 7896 8444 7948
rect 11060 7973 11069 8007
rect 11069 7973 11103 8007
rect 11103 7973 11112 8007
rect 11060 7964 11112 7973
rect 12532 8032 12584 8084
rect 12348 7964 12400 8016
rect 13452 8032 13504 8084
rect 14004 8032 14056 8084
rect 14740 8032 14792 8084
rect 15660 8032 15712 8084
rect 13084 8007 13136 8016
rect 13084 7973 13093 8007
rect 13093 7973 13127 8007
rect 13127 7973 13136 8007
rect 13084 7964 13136 7973
rect 13360 7964 13412 8016
rect 13636 8007 13688 8016
rect 13636 7973 13645 8007
rect 13645 7973 13679 8007
rect 13679 7973 13688 8007
rect 13636 7964 13688 7973
rect 14464 7964 14516 8016
rect 14648 7964 14700 8016
rect 15936 7964 15988 8016
rect 17776 8032 17828 8084
rect 19340 8032 19392 8084
rect 20812 8032 20864 8084
rect 8852 7896 8904 7948
rect 9496 7896 9548 7948
rect 11704 7896 11756 7948
rect 13176 7896 13228 7948
rect 15660 7896 15712 7948
rect 15844 7896 15896 7948
rect 16396 8007 16448 8016
rect 16396 7973 16399 8007
rect 16399 7973 16433 8007
rect 16433 7973 16448 8007
rect 16396 7964 16448 7973
rect 16580 7964 16632 8016
rect 17868 7964 17920 8016
rect 19984 7964 20036 8016
rect 20996 8007 21048 8016
rect 20996 7973 21005 8007
rect 21005 7973 21039 8007
rect 21039 7973 21048 8007
rect 20996 7964 21048 7973
rect 6736 7828 6788 7880
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11152 7828 11204 7880
rect 14188 7871 14240 7880
rect 6920 7760 6972 7812
rect 11060 7760 11112 7812
rect 11336 7760 11388 7812
rect 12532 7760 12584 7812
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 16580 7828 16632 7880
rect 18052 7828 18104 7880
rect 19432 7896 19484 7948
rect 20444 7896 20496 7948
rect 19800 7828 19852 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 7380 7692 7432 7744
rect 8208 7692 8260 7744
rect 8760 7692 8812 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 10140 7692 10192 7744
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 11888 7692 11940 7701
rect 13452 7692 13504 7744
rect 14648 7692 14700 7744
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 14832 7692 14884 7701
rect 14924 7692 14976 7744
rect 15936 7735 15988 7744
rect 15936 7701 15945 7735
rect 15945 7701 15979 7735
rect 15979 7701 15988 7735
rect 15936 7692 15988 7701
rect 18788 7692 18840 7744
rect 19340 7735 19392 7744
rect 19340 7701 19349 7735
rect 19349 7701 19383 7735
rect 19383 7701 19392 7735
rect 19340 7692 19392 7701
rect 21272 7692 21324 7744
rect 21732 7692 21784 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 3240 7488 3292 7540
rect 4160 7420 4212 7472
rect 1216 7352 1268 7404
rect 1584 7352 1636 7404
rect 2964 7352 3016 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 5356 7488 5408 7540
rect 6920 7488 6972 7540
rect 7288 7488 7340 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8484 7488 8536 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 4344 7420 4396 7472
rect 6644 7420 6696 7472
rect 7564 7420 7616 7472
rect 10048 7420 10100 7472
rect 2320 7284 2372 7336
rect 940 7148 992 7200
rect 1676 7216 1728 7268
rect 2688 7216 2740 7268
rect 2320 7148 2372 7200
rect 3056 7216 3108 7268
rect 6736 7352 6788 7404
rect 7656 7352 7708 7404
rect 10876 7352 10928 7404
rect 10968 7352 11020 7404
rect 14648 7420 14700 7472
rect 13728 7352 13780 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15844 7488 15896 7540
rect 16396 7488 16448 7540
rect 15568 7352 15620 7404
rect 17316 7488 17368 7540
rect 20076 7488 20128 7540
rect 20812 7488 20864 7540
rect 19064 7420 19116 7472
rect 19248 7420 19300 7472
rect 20628 7420 20680 7472
rect 23572 7420 23624 7472
rect 19984 7352 20036 7404
rect 20260 7352 20312 7404
rect 23204 7352 23256 7404
rect 6184 7284 6236 7336
rect 3240 7148 3292 7200
rect 3608 7148 3660 7200
rect 5080 7216 5132 7268
rect 5540 7216 5592 7268
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 12348 7284 12400 7336
rect 7380 7216 7432 7268
rect 8208 7216 8260 7268
rect 8576 7216 8628 7268
rect 4436 7148 4488 7200
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 8668 7148 8720 7200
rect 10508 7148 10560 7200
rect 11060 7216 11112 7268
rect 18880 7284 18932 7336
rect 19432 7284 19484 7336
rect 20536 7284 20588 7336
rect 11428 7148 11480 7200
rect 12164 7148 12216 7200
rect 14280 7216 14332 7268
rect 14648 7259 14700 7268
rect 14648 7225 14657 7259
rect 14657 7225 14691 7259
rect 14691 7225 14700 7259
rect 14648 7216 14700 7225
rect 16580 7259 16632 7268
rect 16580 7225 16589 7259
rect 16589 7225 16623 7259
rect 16623 7225 16632 7259
rect 18328 7259 18380 7268
rect 16580 7216 16632 7225
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 13820 7148 13872 7200
rect 15568 7148 15620 7200
rect 16856 7148 16908 7200
rect 18328 7225 18337 7259
rect 18337 7225 18371 7259
rect 18371 7225 18380 7259
rect 18328 7216 18380 7225
rect 19064 7216 19116 7268
rect 19892 7259 19944 7268
rect 19892 7225 19901 7259
rect 19901 7225 19935 7259
rect 19935 7225 19944 7259
rect 19892 7216 19944 7225
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 17960 7148 18012 7200
rect 21916 7148 21968 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 2504 6944 2556 6996
rect 3424 6944 3476 6996
rect 2044 6876 2096 6928
rect 2964 6876 3016 6928
rect 3240 6919 3292 6928
rect 3240 6885 3249 6919
rect 3249 6885 3283 6919
rect 3283 6885 3292 6919
rect 3976 6944 4028 6996
rect 3240 6876 3292 6885
rect 4344 6876 4396 6928
rect 4988 6944 5040 6996
rect 5540 6944 5592 6996
rect 1860 6740 1912 6792
rect 2412 6740 2464 6792
rect 3884 6808 3936 6860
rect 5356 6876 5408 6928
rect 6000 6919 6052 6928
rect 6000 6885 6009 6919
rect 6009 6885 6043 6919
rect 6043 6885 6052 6919
rect 6000 6876 6052 6885
rect 6828 6944 6880 6996
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 8668 6944 8720 6996
rect 12164 6987 12216 6996
rect 12164 6953 12173 6987
rect 12173 6953 12207 6987
rect 12207 6953 12216 6987
rect 12164 6944 12216 6953
rect 13544 6944 13596 6996
rect 15016 6987 15068 6996
rect 15016 6953 15025 6987
rect 15025 6953 15059 6987
rect 15059 6953 15068 6987
rect 15016 6944 15068 6953
rect 16488 6944 16540 6996
rect 17684 6944 17736 6996
rect 18052 6944 18104 6996
rect 18328 6944 18380 6996
rect 19892 6944 19944 6996
rect 6644 6919 6696 6928
rect 6644 6885 6653 6919
rect 6653 6885 6687 6919
rect 6687 6885 6696 6919
rect 6644 6876 6696 6885
rect 7656 6876 7708 6928
rect 8392 6876 8444 6928
rect 8760 6876 8812 6928
rect 11152 6876 11204 6928
rect 13452 6876 13504 6928
rect 13820 6919 13872 6928
rect 13820 6885 13829 6919
rect 13829 6885 13863 6919
rect 13863 6885 13872 6919
rect 13820 6876 13872 6885
rect 14372 6876 14424 6928
rect 15108 6876 15160 6928
rect 16396 6876 16448 6928
rect 17776 6876 17828 6928
rect 19064 6876 19116 6928
rect 20812 6876 20864 6928
rect 4988 6740 5040 6792
rect 7932 6808 7984 6860
rect 8208 6808 8260 6860
rect 10508 6808 10560 6860
rect 11980 6808 12032 6860
rect 8484 6740 8536 6792
rect 9588 6740 9640 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10692 6740 10744 6792
rect 13544 6740 13596 6792
rect 13820 6740 13872 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 5080 6715 5132 6724
rect 3240 6604 3292 6656
rect 3884 6604 3936 6656
rect 3976 6604 4028 6656
rect 4160 6604 4212 6656
rect 5080 6681 5089 6715
rect 5089 6681 5123 6715
rect 5123 6681 5132 6715
rect 5080 6672 5132 6681
rect 5632 6672 5684 6724
rect 6828 6672 6880 6724
rect 8300 6672 8352 6724
rect 10140 6672 10192 6724
rect 10968 6672 11020 6724
rect 15016 6672 15068 6724
rect 16028 6808 16080 6860
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 17776 6740 17828 6792
rect 20720 6740 20772 6792
rect 4712 6604 4764 6656
rect 6092 6604 6144 6656
rect 7840 6604 7892 6656
rect 10692 6604 10744 6656
rect 10876 6604 10928 6656
rect 11520 6604 11572 6656
rect 11888 6604 11940 6656
rect 13728 6604 13780 6656
rect 15292 6604 15344 6656
rect 19616 6672 19668 6724
rect 21640 6672 21692 6724
rect 18236 6604 18288 6656
rect 20076 6647 20128 6656
rect 20076 6613 20085 6647
rect 20085 6613 20119 6647
rect 20119 6613 20128 6647
rect 20076 6604 20128 6613
rect 22100 6604 22152 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 756 6400 808 6452
rect 2412 6400 2464 6452
rect 3056 6443 3108 6452
rect 3056 6409 3065 6443
rect 3065 6409 3099 6443
rect 3099 6409 3108 6443
rect 3056 6400 3108 6409
rect 1400 6332 1452 6384
rect 2596 6332 2648 6384
rect 2688 6332 2740 6384
rect 5632 6400 5684 6452
rect 6000 6400 6052 6452
rect 6276 6400 6328 6452
rect 7104 6400 7156 6452
rect 9312 6400 9364 6452
rect 12256 6443 12308 6452
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 13452 6400 13504 6452
rect 13544 6400 13596 6452
rect 14004 6400 14056 6452
rect 15016 6400 15068 6452
rect 16396 6400 16448 6452
rect 16580 6400 16632 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18512 6400 18564 6452
rect 18696 6400 18748 6452
rect 3976 6332 4028 6384
rect 5080 6332 5132 6384
rect 2228 6264 2280 6316
rect 2872 6264 2924 6316
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 1860 6128 1912 6180
rect 2044 6128 2096 6180
rect 3240 6171 3292 6180
rect 3240 6137 3249 6171
rect 3249 6137 3283 6171
rect 3283 6137 3292 6171
rect 3240 6128 3292 6137
rect 3424 6128 3476 6180
rect 4436 6264 4488 6316
rect 5816 6332 5868 6384
rect 7196 6332 7248 6384
rect 7748 6332 7800 6384
rect 7840 6332 7892 6384
rect 13636 6332 13688 6384
rect 14280 6332 14332 6384
rect 14648 6332 14700 6384
rect 18880 6332 18932 6384
rect 19064 6375 19116 6384
rect 19064 6341 19073 6375
rect 19073 6341 19107 6375
rect 19107 6341 19116 6375
rect 19064 6332 19116 6341
rect 20076 6332 20128 6384
rect 20352 6400 20404 6452
rect 21456 6400 21508 6452
rect 20812 6332 20864 6384
rect 21548 6332 21600 6384
rect 22008 6375 22060 6384
rect 22008 6341 22017 6375
rect 22017 6341 22051 6375
rect 22051 6341 22060 6375
rect 22008 6332 22060 6341
rect 9404 6264 9456 6316
rect 12164 6264 12216 6316
rect 5632 6239 5684 6248
rect 5632 6205 5641 6239
rect 5641 6205 5675 6239
rect 5675 6205 5684 6239
rect 5632 6196 5684 6205
rect 4344 6128 4396 6180
rect 4436 6060 4488 6112
rect 4620 6060 4672 6112
rect 5632 6060 5684 6112
rect 6092 6060 6144 6112
rect 7840 6196 7892 6248
rect 8208 6196 8260 6248
rect 11796 6196 11848 6248
rect 13912 6264 13964 6316
rect 19340 6264 19392 6316
rect 15108 6239 15160 6248
rect 7196 6128 7248 6180
rect 7288 6060 7340 6112
rect 7472 6060 7524 6112
rect 9036 6128 9088 6180
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 10232 6128 10284 6180
rect 9772 6060 9824 6112
rect 10692 6060 10744 6112
rect 10968 6171 11020 6180
rect 10968 6137 10977 6171
rect 10977 6137 11011 6171
rect 11011 6137 11020 6171
rect 10968 6128 11020 6137
rect 11152 6128 11204 6180
rect 12992 6171 13044 6180
rect 12992 6137 13001 6171
rect 13001 6137 13035 6171
rect 13035 6137 13044 6171
rect 12992 6128 13044 6137
rect 13360 6128 13412 6180
rect 13452 6128 13504 6180
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 14280 6128 14332 6180
rect 14464 6128 14516 6180
rect 16396 6128 16448 6180
rect 19248 6196 19300 6248
rect 20720 6196 20772 6248
rect 11060 6060 11112 6112
rect 11704 6060 11756 6112
rect 11980 6060 12032 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 17316 6060 17368 6112
rect 18052 6060 18104 6112
rect 18236 6171 18288 6180
rect 18236 6137 18245 6171
rect 18245 6137 18279 6171
rect 18279 6137 18288 6171
rect 18236 6128 18288 6137
rect 18420 6060 18472 6112
rect 18512 6060 18564 6112
rect 19524 6128 19576 6180
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 1860 5788 1912 5840
rect 2228 5788 2280 5840
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 4068 5856 4120 5908
rect 3148 5788 3200 5840
rect 4344 5831 4396 5840
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 4344 5797 4353 5831
rect 4353 5797 4387 5831
rect 4387 5797 4396 5831
rect 4344 5788 4396 5797
rect 4436 5788 4488 5840
rect 4068 5720 4120 5772
rect 2872 5652 2924 5704
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 1768 5584 1820 5636
rect 3700 5584 3752 5636
rect 4712 5652 4764 5704
rect 3976 5584 4028 5636
rect 8208 5856 8260 5908
rect 8392 5856 8444 5908
rect 10140 5856 10192 5908
rect 10232 5856 10284 5908
rect 5540 5788 5592 5840
rect 6000 5831 6052 5840
rect 6000 5797 6009 5831
rect 6009 5797 6043 5831
rect 6043 5797 6052 5831
rect 6000 5788 6052 5797
rect 6276 5831 6328 5840
rect 6276 5797 6285 5831
rect 6285 5797 6319 5831
rect 6319 5797 6328 5831
rect 6276 5788 6328 5797
rect 6552 5788 6604 5840
rect 9496 5788 9548 5840
rect 13544 5856 13596 5908
rect 13728 5856 13780 5908
rect 14740 5856 14792 5908
rect 16580 5899 16632 5908
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 18236 5856 18288 5908
rect 18328 5856 18380 5908
rect 21364 5856 21416 5908
rect 10692 5788 10744 5840
rect 12164 5788 12216 5840
rect 12716 5831 12768 5840
rect 12716 5797 12725 5831
rect 12725 5797 12759 5831
rect 12759 5797 12768 5831
rect 12716 5788 12768 5797
rect 14188 5788 14240 5840
rect 15660 5831 15712 5840
rect 15660 5797 15669 5831
rect 15669 5797 15703 5831
rect 15703 5797 15712 5831
rect 15660 5788 15712 5797
rect 16028 5788 16080 5840
rect 17776 5788 17828 5840
rect 19064 5788 19116 5840
rect 20444 5788 20496 5840
rect 21640 5831 21692 5840
rect 21640 5797 21649 5831
rect 21649 5797 21683 5831
rect 21683 5797 21692 5831
rect 21640 5788 21692 5797
rect 6920 5720 6972 5772
rect 7288 5763 7340 5772
rect 7288 5729 7297 5763
rect 7297 5729 7331 5763
rect 7331 5729 7340 5763
rect 7288 5720 7340 5729
rect 7656 5720 7708 5772
rect 7932 5720 7984 5772
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 10600 5720 10652 5772
rect 5172 5652 5224 5704
rect 8852 5652 8904 5704
rect 6000 5584 6052 5636
rect 6276 5584 6328 5636
rect 9680 5584 9732 5636
rect 9956 5652 10008 5704
rect 13084 5720 13136 5772
rect 15016 5720 15068 5772
rect 16304 5720 16356 5772
rect 16488 5720 16540 5772
rect 12808 5652 12860 5704
rect 13452 5652 13504 5704
rect 16764 5652 16816 5704
rect 11796 5584 11848 5636
rect 12348 5584 12400 5636
rect 13084 5584 13136 5636
rect 13728 5584 13780 5636
rect 4620 5516 4672 5568
rect 6368 5516 6420 5568
rect 8392 5559 8444 5568
rect 8392 5525 8401 5559
rect 8401 5525 8435 5559
rect 8435 5525 8444 5559
rect 8392 5516 8444 5525
rect 10600 5516 10652 5568
rect 11152 5516 11204 5568
rect 14832 5584 14884 5636
rect 17868 5720 17920 5772
rect 17408 5652 17460 5704
rect 17500 5652 17552 5704
rect 19616 5652 19668 5704
rect 22100 5652 22152 5704
rect 14188 5559 14240 5568
rect 14188 5525 14197 5559
rect 14197 5525 14231 5559
rect 14231 5525 14240 5559
rect 14188 5516 14240 5525
rect 15384 5516 15436 5568
rect 16580 5516 16632 5568
rect 17316 5584 17368 5636
rect 17684 5627 17736 5636
rect 17684 5593 17693 5627
rect 17693 5593 17727 5627
rect 17727 5593 17736 5627
rect 17684 5584 17736 5593
rect 18328 5584 18380 5636
rect 18972 5516 19024 5568
rect 19156 5516 19208 5568
rect 19524 5559 19576 5568
rect 19524 5525 19533 5559
rect 19533 5525 19567 5559
rect 19567 5525 19576 5559
rect 19524 5516 19576 5525
rect 20260 5584 20312 5636
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 296 5312 348 5364
rect 3056 5312 3108 5364
rect 9128 5312 9180 5364
rect 12808 5312 12860 5364
rect 2780 5244 2832 5296
rect 3148 5176 3200 5228
rect 1952 5108 2004 5160
rect 2504 5108 2556 5160
rect 3240 5108 3292 5160
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 3976 5151 4028 5160
rect 3976 5117 3985 5151
rect 3985 5117 4019 5151
rect 4019 5117 4028 5151
rect 3976 5108 4028 5117
rect 4436 5151 4488 5160
rect 4436 5117 4445 5151
rect 4445 5117 4479 5151
rect 4479 5117 4488 5151
rect 4436 5108 4488 5117
rect 5080 5244 5132 5296
rect 5632 5244 5684 5296
rect 7472 5244 7524 5296
rect 8576 5244 8628 5296
rect 9312 5244 9364 5296
rect 9864 5244 9916 5296
rect 10508 5244 10560 5296
rect 7840 5219 7892 5228
rect 2136 5040 2188 5092
rect 3608 5040 3660 5092
rect 4620 5040 4672 5092
rect 5264 5083 5316 5092
rect 5264 5049 5273 5083
rect 5273 5049 5307 5083
rect 5307 5049 5316 5083
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 9496 5176 9548 5228
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 9772 5176 9824 5228
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 12072 5244 12124 5296
rect 15660 5312 15712 5364
rect 20812 5312 20864 5364
rect 14372 5176 14424 5228
rect 15752 5244 15804 5296
rect 16120 5244 16172 5296
rect 17408 5244 17460 5296
rect 17500 5244 17552 5296
rect 17868 5244 17920 5296
rect 19064 5244 19116 5296
rect 19800 5244 19852 5296
rect 20628 5244 20680 5296
rect 18328 5176 18380 5228
rect 15660 5151 15712 5160
rect 5264 5040 5316 5049
rect 5632 5040 5684 5092
rect 6000 5083 6052 5092
rect 1952 4972 2004 5024
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 4344 4972 4396 5024
rect 6000 5049 6009 5083
rect 6009 5049 6043 5083
rect 6043 5049 6052 5083
rect 6000 5040 6052 5049
rect 6368 5040 6420 5092
rect 6644 5040 6696 5092
rect 7012 5083 7064 5092
rect 7012 5049 7021 5083
rect 7021 5049 7055 5083
rect 7055 5049 7064 5083
rect 7012 5040 7064 5049
rect 8300 5040 8352 5092
rect 12072 5040 12124 5092
rect 13084 5040 13136 5092
rect 6736 4972 6788 5024
rect 8116 4972 8168 5024
rect 8392 4972 8444 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 12624 4972 12676 5024
rect 12900 4972 12952 5024
rect 13636 4972 13688 5024
rect 15016 5040 15068 5092
rect 15660 5117 15669 5151
rect 15669 5117 15703 5151
rect 15703 5117 15712 5151
rect 15660 5108 15712 5117
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 17684 5108 17736 5160
rect 18972 5108 19024 5160
rect 16488 5040 16540 5092
rect 17500 5040 17552 5092
rect 22744 5108 22796 5160
rect 16120 4972 16172 5024
rect 16856 4972 16908 5024
rect 17592 4972 17644 5024
rect 20444 4972 20496 5024
rect 22008 5015 22060 5024
rect 22008 4981 22017 5015
rect 22017 4981 22051 5015
rect 22051 4981 22060 5015
rect 22008 4972 22060 4981
rect 22192 4972 22244 5024
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 1768 4811 1820 4820
rect 1768 4777 1777 4811
rect 1777 4777 1811 4811
rect 1811 4777 1820 4811
rect 1768 4768 1820 4777
rect 3424 4768 3476 4820
rect 4344 4768 4396 4820
rect 5356 4768 5408 4820
rect 5632 4768 5684 4820
rect 6368 4768 6420 4820
rect 2780 4700 2832 4752
rect 3884 4700 3936 4752
rect 4620 4700 4672 4752
rect 4804 4700 4856 4752
rect 6644 4743 6696 4752
rect 388 4632 440 4684
rect 3516 4632 3568 4684
rect 4528 4675 4580 4684
rect 1492 4564 1544 4616
rect 3976 4564 4028 4616
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 5172 4632 5224 4684
rect 5356 4632 5408 4684
rect 5540 4632 5592 4684
rect 4436 4564 4488 4616
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 5632 4564 5684 4616
rect 6184 4607 6236 4616
rect 4252 4496 4304 4548
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6276 4564 6328 4616
rect 6644 4709 6653 4743
rect 6653 4709 6687 4743
rect 6687 4709 6696 4743
rect 6644 4700 6696 4709
rect 7380 4768 7432 4820
rect 8484 4768 8536 4820
rect 11060 4768 11112 4820
rect 14096 4768 14148 4820
rect 14372 4768 14424 4820
rect 16856 4768 16908 4820
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 17868 4768 17920 4820
rect 7104 4700 7156 4752
rect 7288 4700 7340 4752
rect 7564 4743 7616 4752
rect 7564 4709 7573 4743
rect 7573 4709 7607 4743
rect 7607 4709 7616 4743
rect 7564 4700 7616 4709
rect 8116 4743 8168 4752
rect 8116 4709 8125 4743
rect 8125 4709 8159 4743
rect 8159 4709 8168 4743
rect 8116 4700 8168 4709
rect 8300 4700 8352 4752
rect 4436 4428 4488 4480
rect 4528 4428 4580 4480
rect 4712 4428 4764 4480
rect 5632 4428 5684 4480
rect 7656 4564 7708 4616
rect 7196 4539 7248 4548
rect 7196 4505 7205 4539
rect 7205 4505 7239 4539
rect 7239 4505 7248 4539
rect 7196 4496 7248 4505
rect 7748 4496 7800 4548
rect 8668 4700 8720 4752
rect 11152 4700 11204 4752
rect 12624 4700 12676 4752
rect 13268 4743 13320 4752
rect 13268 4709 13277 4743
rect 13277 4709 13311 4743
rect 13311 4709 13320 4743
rect 13268 4700 13320 4709
rect 14188 4700 14240 4752
rect 9496 4632 9548 4684
rect 12256 4632 12308 4684
rect 13084 4632 13136 4684
rect 14464 4632 14516 4684
rect 8576 4564 8628 4616
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 9864 4564 9916 4616
rect 12808 4564 12860 4616
rect 13636 4564 13688 4616
rect 15292 4564 15344 4616
rect 8576 4428 8628 4480
rect 9588 4496 9640 4548
rect 13544 4496 13596 4548
rect 16304 4700 16356 4752
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 19432 4700 19484 4752
rect 20812 4700 20864 4752
rect 21640 4743 21692 4752
rect 21640 4709 21649 4743
rect 21649 4709 21683 4743
rect 21683 4709 21692 4743
rect 21640 4700 21692 4709
rect 17592 4564 17644 4616
rect 19064 4564 19116 4616
rect 19984 4632 20036 4684
rect 20168 4675 20220 4684
rect 20168 4641 20177 4675
rect 20177 4641 20211 4675
rect 20211 4641 20220 4675
rect 20168 4632 20220 4641
rect 20352 4632 20404 4684
rect 20628 4632 20680 4684
rect 20076 4564 20128 4616
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 21916 4564 21968 4616
rect 16212 4496 16264 4548
rect 12164 4428 12216 4480
rect 12624 4428 12676 4480
rect 13360 4428 13412 4480
rect 13728 4428 13780 4480
rect 14096 4428 14148 4480
rect 14832 4428 14884 4480
rect 15568 4428 15620 4480
rect 18972 4496 19024 4548
rect 17684 4428 17736 4480
rect 18144 4428 18196 4480
rect 19616 4428 19668 4480
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 2688 4199 2740 4208
rect 2688 4165 2697 4199
rect 2697 4165 2731 4199
rect 2731 4165 2740 4199
rect 2688 4156 2740 4165
rect 4344 4156 4396 4208
rect 3056 4088 3108 4140
rect 7104 4224 7156 4276
rect 7380 4156 7432 4208
rect 8116 4224 8168 4276
rect 9312 4224 9364 4276
rect 8852 4156 8904 4208
rect 9588 4156 9640 4208
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 3332 4020 3384 4072
rect 3884 4020 3936 4072
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 5908 4020 5960 4072
rect 6184 4020 6236 4072
rect 6552 4020 6604 4072
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 7196 4020 7248 4072
rect 7564 4020 7616 4072
rect 1768 3884 1820 3936
rect 3240 3884 3292 3936
rect 3332 3884 3384 3936
rect 3700 3952 3752 4004
rect 6736 3952 6788 4004
rect 8116 3952 8168 4004
rect 8668 3995 8720 4004
rect 8668 3961 8677 3995
rect 8677 3961 8711 3995
rect 8711 3961 8720 3995
rect 8668 3952 8720 3961
rect 9220 3952 9272 4004
rect 4804 3884 4856 3936
rect 5264 3884 5316 3936
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6644 3884 6696 3936
rect 6828 3884 6880 3936
rect 7196 3884 7248 3936
rect 7748 3884 7800 3936
rect 8300 3884 8352 3936
rect 10324 3995 10376 4004
rect 10324 3961 10333 3995
rect 10333 3961 10367 3995
rect 10367 3961 10376 3995
rect 13636 4224 13688 4276
rect 13912 4224 13964 4276
rect 14648 4224 14700 4276
rect 15108 4224 15160 4276
rect 11796 4199 11848 4208
rect 11796 4165 11805 4199
rect 11805 4165 11839 4199
rect 11839 4165 11848 4199
rect 11796 4156 11848 4165
rect 13268 4156 13320 4208
rect 14832 4199 14884 4208
rect 14832 4165 14841 4199
rect 14841 4165 14875 4199
rect 14875 4165 14884 4199
rect 14832 4156 14884 4165
rect 16304 4224 16356 4276
rect 16856 4224 16908 4276
rect 19064 4224 19116 4276
rect 19524 4224 19576 4276
rect 11152 4088 11204 4140
rect 11980 4088 12032 4140
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 14740 4088 14792 4140
rect 16212 4088 16264 4140
rect 17408 4131 17460 4140
rect 11244 4020 11296 4072
rect 10324 3952 10376 3961
rect 11060 3884 11112 3936
rect 11244 3884 11296 3936
rect 11612 4020 11664 4072
rect 12256 4020 12308 4072
rect 12716 4020 12768 4072
rect 14280 4020 14332 4072
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 18788 4088 18840 4140
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 13636 3995 13688 4004
rect 13636 3961 13645 3995
rect 13645 3961 13679 3995
rect 13679 3961 13688 3995
rect 13636 3952 13688 3961
rect 15016 3952 15068 4004
rect 15292 3952 15344 4004
rect 14372 3884 14424 3936
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 17960 3952 18012 4004
rect 18144 3995 18196 4004
rect 18144 3961 18153 3995
rect 18153 3961 18187 3995
rect 18187 3961 18196 3995
rect 18144 3952 18196 3961
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 18788 3952 18840 4004
rect 19800 4156 19852 4208
rect 20812 4224 20864 4276
rect 21640 4224 21692 4276
rect 21916 4224 21968 4276
rect 22376 4267 22428 4276
rect 22376 4233 22385 4267
rect 22385 4233 22419 4267
rect 22419 4233 22428 4267
rect 22376 4224 22428 4233
rect 18972 4020 19024 4072
rect 16488 3884 16540 3936
rect 20352 4020 20404 4072
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 19616 3884 19668 3936
rect 19800 3995 19852 4004
rect 19800 3961 19809 3995
rect 19809 3961 19843 3995
rect 19843 3961 19852 3995
rect 19800 3952 19852 3961
rect 19892 3884 19944 3936
rect 21732 3884 21784 3936
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 3240 3680 3292 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 5356 3680 5408 3732
rect 7012 3680 7064 3732
rect 8300 3680 8352 3732
rect 9956 3680 10008 3732
rect 10692 3680 10744 3732
rect 2872 3612 2924 3664
rect 1032 3544 1084 3596
rect 1952 3544 2004 3596
rect 4068 3544 4120 3596
rect 2688 3476 2740 3528
rect 4160 3408 4212 3460
rect 5264 3612 5316 3664
rect 6368 3655 6420 3664
rect 6368 3621 6377 3655
rect 6377 3621 6411 3655
rect 6411 3621 6420 3655
rect 6368 3612 6420 3621
rect 7748 3612 7800 3664
rect 7932 3612 7984 3664
rect 9036 3612 9088 3664
rect 9864 3612 9916 3664
rect 5816 3544 5868 3596
rect 9128 3587 9180 3596
rect 5724 3476 5776 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7472 3476 7524 3528
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 9496 3544 9548 3596
rect 9680 3587 9732 3596
rect 9680 3553 9724 3587
rect 9724 3553 9732 3587
rect 9680 3544 9732 3553
rect 11704 3612 11756 3664
rect 12900 3680 12952 3732
rect 13268 3680 13320 3732
rect 13636 3680 13688 3732
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 15476 3723 15528 3732
rect 15476 3689 15485 3723
rect 15485 3689 15519 3723
rect 15519 3689 15528 3723
rect 15476 3680 15528 3689
rect 16120 3680 16172 3732
rect 15752 3612 15804 3664
rect 17408 3680 17460 3732
rect 16856 3612 16908 3664
rect 18052 3680 18104 3732
rect 19156 3723 19208 3732
rect 19156 3689 19165 3723
rect 19165 3689 19199 3723
rect 19199 3689 19208 3723
rect 19156 3680 19208 3689
rect 19708 3723 19760 3732
rect 19708 3689 19717 3723
rect 19717 3689 19751 3723
rect 19751 3689 19760 3723
rect 19708 3680 19760 3689
rect 20536 3723 20588 3732
rect 20536 3689 20545 3723
rect 20545 3689 20579 3723
rect 20579 3689 20588 3723
rect 20536 3680 20588 3689
rect 20628 3680 20680 3732
rect 18236 3612 18288 3664
rect 20444 3612 20496 3664
rect 20812 3612 20864 3664
rect 10232 3476 10284 3528
rect 10692 3544 10744 3596
rect 11152 3544 11204 3596
rect 13912 3544 13964 3596
rect 15568 3544 15620 3596
rect 16120 3544 16172 3596
rect 16212 3544 16264 3596
rect 18052 3544 18104 3596
rect 18328 3544 18380 3596
rect 18696 3544 18748 3596
rect 6736 3408 6788 3460
rect 7656 3408 7708 3460
rect 9588 3408 9640 3460
rect 10784 3476 10836 3528
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 13728 3476 13780 3528
rect 16580 3476 16632 3528
rect 19432 3476 19484 3528
rect 20720 3476 20772 3528
rect 21180 3476 21232 3528
rect 10968 3408 11020 3460
rect 11060 3408 11112 3460
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 8760 3340 8812 3392
rect 11428 3340 11480 3392
rect 11704 3383 11756 3392
rect 11704 3349 11713 3383
rect 11713 3349 11747 3383
rect 11747 3349 11756 3383
rect 11704 3340 11756 3349
rect 13636 3408 13688 3460
rect 21916 3476 21968 3528
rect 14280 3340 14332 3392
rect 15752 3340 15804 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 18144 3340 18196 3392
rect 19524 3383 19576 3392
rect 19524 3349 19533 3383
rect 19533 3349 19567 3383
rect 19567 3349 19576 3383
rect 19524 3340 19576 3349
rect 22284 3383 22336 3392
rect 22284 3349 22293 3383
rect 22293 3349 22327 3383
rect 22327 3349 22336 3383
rect 22284 3340 22336 3349
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 1124 3068 1176 3120
rect 7288 3136 7340 3188
rect 7564 3136 7616 3188
rect 8208 3136 8260 3188
rect 9496 3136 9548 3188
rect 10692 3136 10744 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 6552 3068 6604 3120
rect 7104 3000 7156 3052
rect 9772 3068 9824 3120
rect 9956 3111 10008 3120
rect 9956 3077 9965 3111
rect 9965 3077 9999 3111
rect 9999 3077 10008 3111
rect 9956 3068 10008 3077
rect 10048 3068 10100 3120
rect 12072 3136 12124 3188
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 9404 3000 9456 3052
rect 10416 3000 10468 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 11336 3000 11388 3052
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 2504 2932 2556 2984
rect 3976 2864 4028 2916
rect 4528 2864 4580 2916
rect 6368 2932 6420 2984
rect 6460 2975 6512 2984
rect 6460 2941 6469 2975
rect 6469 2941 6503 2975
rect 6503 2941 6512 2975
rect 6460 2932 6512 2941
rect 5724 2907 5776 2916
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 3332 2839 3384 2848
rect 3332 2805 3341 2839
rect 3341 2805 3375 2839
rect 3375 2805 3384 2839
rect 3332 2796 3384 2805
rect 5356 2839 5408 2848
rect 5356 2805 5365 2839
rect 5365 2805 5399 2839
rect 5399 2805 5408 2839
rect 5356 2796 5408 2805
rect 5724 2873 5733 2907
rect 5733 2873 5767 2907
rect 5767 2873 5776 2907
rect 5724 2864 5776 2873
rect 6000 2864 6052 2916
rect 7196 2932 7248 2984
rect 7472 2932 7524 2984
rect 11796 3068 11848 3120
rect 13268 3111 13320 3120
rect 13268 3077 13277 3111
rect 13277 3077 13311 3111
rect 13311 3077 13320 3111
rect 13268 3068 13320 3077
rect 14372 3136 14424 3188
rect 17868 3136 17920 3188
rect 15292 3068 15344 3120
rect 15660 3111 15712 3120
rect 15660 3077 15669 3111
rect 15669 3077 15703 3111
rect 15703 3077 15712 3111
rect 15660 3068 15712 3077
rect 15752 3068 15804 3120
rect 17316 3068 17368 3120
rect 13544 3000 13596 3052
rect 13728 3000 13780 3052
rect 14740 3000 14792 3052
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 18512 3068 18564 3120
rect 19064 3000 19116 3052
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 19892 3000 19944 3052
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 7748 2864 7800 2916
rect 6460 2796 6512 2848
rect 6828 2796 6880 2848
rect 7012 2796 7064 2848
rect 8208 2864 8260 2916
rect 8944 2864 8996 2916
rect 9220 2864 9272 2916
rect 10324 2907 10376 2916
rect 10324 2873 10333 2907
rect 10333 2873 10367 2907
rect 10367 2873 10376 2907
rect 10324 2864 10376 2873
rect 11152 2907 11204 2916
rect 11152 2873 11161 2907
rect 11161 2873 11195 2907
rect 11195 2873 11204 2907
rect 11152 2864 11204 2873
rect 12348 2864 12400 2916
rect 12624 2932 12676 2984
rect 13360 2932 13412 2984
rect 14464 2932 14516 2984
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 13544 2907 13596 2916
rect 9680 2796 9732 2848
rect 11060 2796 11112 2848
rect 11244 2796 11296 2848
rect 11796 2796 11848 2848
rect 12164 2796 12216 2848
rect 13544 2873 13553 2907
rect 13553 2873 13587 2907
rect 13587 2873 13596 2907
rect 13544 2864 13596 2873
rect 13728 2864 13780 2916
rect 15108 2907 15160 2916
rect 15108 2873 15117 2907
rect 15117 2873 15151 2907
rect 15151 2873 15160 2907
rect 15108 2864 15160 2873
rect 15568 2864 15620 2916
rect 15844 2864 15896 2916
rect 17868 2864 17920 2916
rect 18144 2907 18196 2916
rect 18144 2873 18153 2907
rect 18153 2873 18187 2907
rect 18187 2873 18196 2907
rect 18144 2864 18196 2873
rect 18236 2907 18288 2916
rect 18236 2873 18245 2907
rect 18245 2873 18279 2907
rect 18279 2873 18288 2907
rect 18236 2864 18288 2873
rect 19524 2864 19576 2916
rect 22100 2907 22152 2916
rect 13820 2796 13872 2848
rect 16120 2796 16172 2848
rect 16856 2796 16908 2848
rect 18328 2796 18380 2848
rect 19340 2796 19392 2848
rect 22100 2873 22109 2907
rect 22109 2873 22143 2907
rect 22143 2873 22152 2907
rect 22100 2864 22152 2873
rect 20812 2796 20864 2848
rect 21364 2839 21416 2848
rect 21364 2805 21373 2839
rect 21373 2805 21407 2839
rect 21407 2805 21416 2839
rect 21364 2796 21416 2805
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 2596 2592 2648 2644
rect 6184 2592 6236 2644
rect 1768 2567 1820 2576
rect 1768 2533 1771 2567
rect 1771 2533 1805 2567
rect 1805 2533 1820 2567
rect 1768 2524 1820 2533
rect 2780 2524 2832 2576
rect 3976 2524 4028 2576
rect 5724 2524 5776 2576
rect 204 2456 256 2508
rect 3516 2456 3568 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 6092 2499 6144 2508
rect 6092 2465 6101 2499
rect 6101 2465 6135 2499
rect 6135 2465 6144 2499
rect 6092 2456 6144 2465
rect 7012 2524 7064 2576
rect 8024 2592 8076 2644
rect 10600 2592 10652 2644
rect 7656 2524 7708 2576
rect 8116 2567 8168 2576
rect 8116 2533 8125 2567
rect 8125 2533 8159 2567
rect 8159 2533 8168 2567
rect 8116 2524 8168 2533
rect 8852 2567 8904 2576
rect 8852 2533 8861 2567
rect 8861 2533 8895 2567
rect 8895 2533 8904 2567
rect 8852 2524 8904 2533
rect 8944 2567 8996 2576
rect 8944 2533 8953 2567
rect 8953 2533 8987 2567
rect 8987 2533 8996 2567
rect 9496 2567 9548 2576
rect 8944 2524 8996 2533
rect 9496 2533 9505 2567
rect 9505 2533 9539 2567
rect 9539 2533 9548 2567
rect 9496 2524 9548 2533
rect 9864 2567 9916 2576
rect 9864 2533 9873 2567
rect 9873 2533 9907 2567
rect 9907 2533 9916 2567
rect 9864 2524 9916 2533
rect 10140 2524 10192 2576
rect 12164 2592 12216 2644
rect 14004 2635 14056 2644
rect 11980 2524 12032 2576
rect 7840 2456 7892 2508
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 14740 2592 14792 2644
rect 12808 2567 12860 2576
rect 12808 2533 12817 2567
rect 12817 2533 12851 2567
rect 12851 2533 12860 2567
rect 17316 2592 17368 2644
rect 17684 2635 17736 2644
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 18696 2592 18748 2644
rect 21824 2592 21876 2644
rect 12808 2524 12860 2533
rect 16120 2524 16172 2576
rect 16672 2524 16724 2576
rect 18420 2567 18472 2576
rect 18420 2533 18429 2567
rect 18429 2533 18463 2567
rect 18463 2533 18472 2567
rect 18420 2524 18472 2533
rect 18512 2567 18564 2576
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 18880 2524 18932 2576
rect 13360 2456 13412 2508
rect 848 2388 900 2440
rect 4252 2320 4304 2372
rect 480 2252 532 2304
rect 5448 2252 5500 2304
rect 5540 2252 5592 2304
rect 7564 2388 7616 2440
rect 8392 2320 8444 2372
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 11612 2388 11664 2440
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 12900 2388 12952 2440
rect 14740 2456 14792 2508
rect 15844 2456 15896 2508
rect 18236 2456 18288 2508
rect 19064 2499 19116 2508
rect 19064 2465 19073 2499
rect 19073 2465 19107 2499
rect 19107 2465 19116 2499
rect 19064 2456 19116 2465
rect 20260 2456 20312 2508
rect 21272 2456 21324 2508
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 10048 2252 10100 2304
rect 15568 2320 15620 2372
rect 16856 2363 16908 2372
rect 16856 2329 16865 2363
rect 16865 2329 16899 2363
rect 16899 2329 16908 2363
rect 16856 2320 16908 2329
rect 18512 2320 18564 2372
rect 19248 2320 19300 2372
rect 13452 2252 13504 2304
rect 13544 2252 13596 2304
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 14740 2295 14792 2304
rect 14740 2261 14749 2295
rect 14749 2261 14783 2295
rect 14783 2261 14792 2295
rect 14740 2252 14792 2261
rect 18788 2252 18840 2304
rect 19708 2295 19760 2304
rect 19708 2261 19717 2295
rect 19717 2261 19751 2295
rect 19751 2261 19760 2295
rect 19708 2252 19760 2261
rect 19800 2252 19852 2304
rect 21732 2295 21784 2304
rect 21732 2261 21741 2295
rect 21741 2261 21775 2295
rect 21775 2261 21784 2295
rect 21732 2252 21784 2261
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 6276 2048 6328 2100
rect 11520 2048 11572 2100
rect 12072 2048 12124 2100
rect 16212 2048 16264 2100
rect 112 1980 164 2032
rect 4804 1980 4856 2032
rect 940 1912 992 1964
rect 6736 1980 6788 2032
rect 8944 1980 8996 2032
rect 14464 1980 14516 2032
rect 22192 1980 22244 2032
rect 5356 1912 5408 1964
rect 15384 1912 15436 1964
rect 4712 1844 4764 1896
rect 9312 1844 9364 1896
rect 11704 1844 11756 1896
rect 4252 1776 4304 1828
rect 10140 1776 10192 1828
rect 2412 76 2464 128
rect 16764 76 16816 128
rect 17408 76 17460 128
rect 14464 8 14516 60
rect 21364 8 21416 60
<< metal2 >>
rect 938 23610 994 24000
rect 2778 23610 2834 24000
rect 4618 23610 4674 24000
rect 6458 23610 6514 24000
rect 938 23582 1256 23610
rect 938 23520 994 23582
rect 846 23216 902 23225
rect 846 23151 902 23160
rect 572 22976 624 22982
rect 572 22918 624 22924
rect 386 21584 442 21593
rect 386 21519 442 21528
rect 202 20632 258 20641
rect 202 20567 258 20576
rect 112 20256 164 20262
rect 18 20224 74 20233
rect 112 20198 164 20204
rect 18 20159 74 20168
rect 32 18970 60 20159
rect 20 18964 72 18970
rect 20 18906 72 18912
rect 20 17468 72 17474
rect 20 17410 72 17416
rect 32 14657 60 17410
rect 124 17105 152 20198
rect 110 17096 166 17105
rect 110 17031 166 17040
rect 110 16280 166 16289
rect 110 16215 166 16224
rect 124 16182 152 16215
rect 112 16176 164 16182
rect 112 16118 164 16124
rect 112 16040 164 16046
rect 112 15982 164 15988
rect 18 14648 74 14657
rect 18 14583 74 14592
rect 32 12850 60 14583
rect 20 12844 72 12850
rect 20 12786 72 12792
rect 18 12608 74 12617
rect 18 12543 74 12552
rect 32 11937 60 12543
rect 18 11928 74 11937
rect 18 11863 74 11872
rect 20 11824 72 11830
rect 20 11766 72 11772
rect 32 11529 60 11766
rect 18 11520 74 11529
rect 18 11455 74 11464
rect 124 8974 152 15982
rect 216 11762 244 20567
rect 294 17368 350 17377
rect 294 17303 350 17312
rect 308 14958 336 17303
rect 296 14952 348 14958
rect 296 14894 348 14900
rect 296 14748 348 14754
rect 296 14690 348 14696
rect 204 11756 256 11762
rect 204 11698 256 11704
rect 204 11212 256 11218
rect 204 11154 256 11160
rect 112 8968 164 8974
rect 112 8910 164 8916
rect 112 8560 164 8566
rect 112 8502 164 8508
rect 20 8356 72 8362
rect 20 8298 72 8304
rect 32 5137 60 8298
rect 124 7449 152 8502
rect 110 7440 166 7449
rect 110 7375 166 7384
rect 18 5128 74 5137
rect 18 5063 74 5072
rect 32 4154 60 5063
rect 32 4126 152 4154
rect 124 2038 152 4126
rect 216 2514 244 11154
rect 308 5370 336 14690
rect 400 13258 428 21519
rect 478 19952 534 19961
rect 478 19887 534 19896
rect 388 13252 440 13258
rect 388 13194 440 13200
rect 386 12880 442 12889
rect 386 12815 442 12824
rect 296 5364 348 5370
rect 296 5306 348 5312
rect 400 4690 428 12815
rect 388 4684 440 4690
rect 388 4626 440 4632
rect 204 2508 256 2514
rect 204 2450 256 2456
rect 492 2310 520 19887
rect 584 17592 612 22918
rect 754 22672 810 22681
rect 754 22607 810 22616
rect 584 17564 704 17592
rect 570 17504 626 17513
rect 570 17439 626 17448
rect 584 14618 612 17439
rect 676 17377 704 17564
rect 662 17368 718 17377
rect 662 17303 718 17312
rect 664 16788 716 16794
rect 664 16730 716 16736
rect 676 16697 704 16730
rect 662 16688 718 16697
rect 662 16623 718 16632
rect 662 16552 718 16561
rect 662 16487 718 16496
rect 572 14612 624 14618
rect 572 14554 624 14560
rect 572 14476 624 14482
rect 572 14418 624 14424
rect 584 9994 612 14418
rect 572 9988 624 9994
rect 572 9930 624 9936
rect 570 9888 626 9897
rect 570 9823 626 9832
rect 584 9790 612 9823
rect 572 9784 624 9790
rect 572 9726 624 9732
rect 572 9686 624 9692
rect 572 9628 624 9634
rect 480 2304 532 2310
rect 480 2246 532 2252
rect 112 2032 164 2038
rect 112 1974 164 1980
rect 584 1601 612 9628
rect 676 7818 704 16487
rect 768 15434 796 22607
rect 860 18057 888 23151
rect 1124 22908 1176 22914
rect 1124 22850 1176 22856
rect 940 22840 992 22846
rect 940 22782 992 22788
rect 952 18329 980 22782
rect 1032 22228 1084 22234
rect 1032 22170 1084 22176
rect 938 18320 994 18329
rect 938 18255 994 18264
rect 940 18080 992 18086
rect 846 18048 902 18057
rect 940 18022 992 18028
rect 846 17983 902 17992
rect 846 16824 902 16833
rect 846 16759 902 16768
rect 756 15428 808 15434
rect 756 15370 808 15376
rect 754 14512 810 14521
rect 754 14447 810 14456
rect 664 7812 716 7818
rect 664 7754 716 7760
rect 768 6458 796 14447
rect 860 11506 888 16759
rect 952 11626 980 18022
rect 940 11620 992 11626
rect 940 11562 992 11568
rect 860 11478 980 11506
rect 848 11348 900 11354
rect 848 11290 900 11296
rect 756 6452 808 6458
rect 756 6394 808 6400
rect 860 2446 888 11290
rect 952 8294 980 11478
rect 1044 8906 1072 22170
rect 1136 15570 1164 22850
rect 1228 21418 1256 23582
rect 2778 23594 2912 23610
rect 2778 23588 2924 23594
rect 2778 23582 2872 23588
rect 2778 23520 2834 23582
rect 2872 23530 2924 23536
rect 4618 23582 4936 23610
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 1398 22944 1454 22953
rect 1398 22879 1454 22888
rect 1306 22400 1362 22409
rect 1306 22335 1362 22344
rect 1216 21412 1268 21418
rect 1216 21354 1268 21360
rect 1216 19712 1268 19718
rect 1216 19654 1268 19660
rect 1228 19310 1256 19654
rect 1216 19304 1268 19310
rect 1216 19246 1268 19252
rect 1228 16969 1256 19246
rect 1214 16960 1270 16969
rect 1214 16895 1270 16904
rect 1124 15564 1176 15570
rect 1124 15506 1176 15512
rect 1124 15428 1176 15434
rect 1124 15370 1176 15376
rect 1136 13938 1164 15370
rect 1216 14884 1268 14890
rect 1216 14826 1268 14832
rect 1124 13932 1176 13938
rect 1124 13874 1176 13880
rect 1124 13728 1176 13734
rect 1124 13670 1176 13676
rect 1136 13530 1164 13670
rect 1124 13524 1176 13530
rect 1124 13466 1176 13472
rect 1122 13288 1178 13297
rect 1122 13223 1124 13232
rect 1176 13223 1178 13232
rect 1124 13194 1176 13200
rect 1032 8900 1084 8906
rect 1032 8842 1084 8848
rect 1136 8786 1164 13194
rect 1228 12345 1256 14826
rect 1320 14482 1348 22335
rect 1412 21486 1440 22879
rect 1674 22808 1730 22817
rect 1674 22743 1730 22752
rect 2044 22772 2096 22778
rect 1492 22568 1544 22574
rect 1492 22510 1544 22516
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21146 1440 21422
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 1504 18408 1532 22510
rect 1582 21312 1638 21321
rect 1582 21247 1638 21256
rect 1412 18380 1532 18408
rect 1412 15502 1440 18380
rect 1490 18320 1546 18329
rect 1490 18255 1546 18264
rect 1504 17542 1532 18255
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1320 14074 1348 14418
rect 1308 14068 1360 14074
rect 1308 14010 1360 14016
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1214 12336 1270 12345
rect 1214 12271 1270 12280
rect 1214 10976 1270 10985
rect 1214 10911 1270 10920
rect 1228 10810 1256 10911
rect 1216 10804 1268 10810
rect 1216 10746 1268 10752
rect 1214 9208 1270 9217
rect 1320 9178 1348 13874
rect 1412 12306 1440 14991
rect 1504 13394 1532 16934
rect 1596 16794 1624 21247
rect 1688 20058 1716 22743
rect 2044 22714 2096 22720
rect 1860 22704 1912 22710
rect 1860 22646 1912 22652
rect 1768 21004 1820 21010
rect 1768 20946 1820 20952
rect 1780 20058 1808 20946
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 18222 1716 18566
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1582 15192 1638 15201
rect 1582 15127 1638 15136
rect 1596 15094 1624 15127
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 13394 1624 14311
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1688 13274 1716 17818
rect 1780 16046 1808 19790
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1780 15706 1808 15982
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1504 13246 1716 13274
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1400 11620 1452 11626
rect 1400 11562 1452 11568
rect 1412 11121 1440 11562
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1412 9586 1440 11047
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1504 9518 1532 13246
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1596 10713 1624 12922
rect 1688 12646 1716 13126
rect 1780 12986 1808 15506
rect 1872 14618 1900 22646
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1964 14464 1992 22578
rect 2056 19145 2084 22714
rect 2240 21690 2268 22986
rect 2596 21888 2648 21894
rect 2596 21830 2648 21836
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 2608 21418 2636 21830
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2136 21344 2188 21350
rect 2136 21286 2188 21292
rect 2318 21312 2374 21321
rect 2148 20233 2176 21286
rect 2318 21247 2374 21256
rect 2226 21176 2282 21185
rect 2226 21111 2282 21120
rect 2134 20224 2190 20233
rect 2134 20159 2190 20168
rect 2134 20088 2190 20097
rect 2134 20023 2190 20032
rect 2148 19446 2176 20023
rect 2240 19825 2268 21111
rect 2332 19922 2360 21247
rect 2608 21078 2636 21354
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2412 20868 2464 20874
rect 2412 20810 2464 20816
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2226 19816 2282 19825
rect 2226 19751 2282 19760
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2240 19514 2268 19654
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2042 19136 2098 19145
rect 2042 19071 2098 19080
rect 2148 18986 2176 19246
rect 2056 18958 2176 18986
rect 2056 18698 2084 18958
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2044 18692 2096 18698
rect 2044 18634 2096 18640
rect 2056 18222 2084 18634
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 2056 16794 2084 17206
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2042 16688 2098 16697
rect 2148 16658 2176 18838
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2240 17610 2268 18770
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2226 17504 2282 17513
rect 2226 17439 2282 17448
rect 2240 17338 2268 17439
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2226 17096 2282 17105
rect 2226 17031 2282 17040
rect 2042 16623 2098 16632
rect 2136 16652 2188 16658
rect 2056 15094 2084 16623
rect 2136 16594 2188 16600
rect 2148 16250 2176 16594
rect 2240 16590 2268 17031
rect 2332 16674 2360 19654
rect 2424 17241 2452 20810
rect 2608 19922 2636 21014
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2792 20777 2820 20946
rect 2778 20768 2834 20777
rect 2778 20703 2834 20712
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2504 19780 2556 19786
rect 2504 19722 2556 19728
rect 2516 19689 2544 19722
rect 2502 19680 2558 19689
rect 2502 19615 2558 19624
rect 2608 19446 2636 19858
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2410 17232 2466 17241
rect 2410 17167 2466 17176
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2424 16794 2452 17070
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2332 16646 2452 16674
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2226 16280 2282 16289
rect 2136 16244 2188 16250
rect 2226 16215 2282 16224
rect 2136 16186 2188 16192
rect 2044 15088 2096 15094
rect 2044 15030 2096 15036
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 2056 14618 2084 14894
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 1964 14436 2084 14464
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1860 14272 1912 14278
rect 1964 14249 1992 14282
rect 1860 14214 1912 14220
rect 1950 14240 2006 14249
rect 1872 13512 1900 14214
rect 1950 14175 2006 14184
rect 2056 13814 2084 14436
rect 2148 13938 2176 16186
rect 2240 15026 2268 16215
rect 2318 16144 2374 16153
rect 2318 16079 2374 16088
rect 2332 15638 2360 16079
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2240 14929 2268 14962
rect 2226 14920 2282 14929
rect 2226 14855 2282 14864
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2056 13786 2176 13814
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 1872 13484 1992 13512
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 12640 1728 12646
rect 1780 12617 1808 12786
rect 1676 12582 1728 12588
rect 1766 12608 1822 12617
rect 1582 10704 1638 10713
rect 1582 10639 1638 10648
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1490 9344 1546 9353
rect 1490 9279 1546 9288
rect 1214 9143 1270 9152
rect 1308 9172 1360 9178
rect 1228 9110 1256 9143
rect 1308 9114 1360 9120
rect 1216 9104 1268 9110
rect 1216 9046 1268 9052
rect 1214 8936 1270 8945
rect 1214 8871 1270 8880
rect 1044 8758 1164 8786
rect 940 8288 992 8294
rect 940 8230 992 8236
rect 940 7200 992 7206
rect 940 7142 992 7148
rect 848 2440 900 2446
rect 848 2382 900 2388
rect 952 1970 980 7142
rect 1044 3602 1072 8758
rect 1122 8392 1178 8401
rect 1122 8327 1178 8336
rect 1032 3596 1084 3602
rect 1032 3538 1084 3544
rect 1136 3126 1164 8327
rect 1228 7410 1256 8871
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 8634 1440 8774
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8129 1440 8366
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1400 7812 1452 7818
rect 1400 7754 1452 7760
rect 1216 7404 1268 7410
rect 1216 7346 1268 7352
rect 1412 6390 1440 7754
rect 1504 7750 1532 9279
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1596 7410 1624 8978
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1400 6384 1452 6390
rect 1596 6361 1624 7346
rect 1688 7274 1716 12582
rect 1766 12543 1822 12552
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1780 11286 1808 11494
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1780 11014 1808 11222
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10470 1808 10950
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 8906 1808 9522
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1780 8809 1808 8842
rect 1766 8800 1822 8809
rect 1766 8735 1822 8744
rect 1872 8242 1900 13330
rect 1964 12714 1992 13484
rect 2056 13258 2084 13670
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2148 13002 2176 13786
rect 2056 12974 2176 13002
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1950 12064 2006 12073
rect 1950 11999 2006 12008
rect 1964 8634 1992 11999
rect 2056 9586 2084 12974
rect 2134 12744 2190 12753
rect 2134 12679 2190 12688
rect 2148 12442 2176 12679
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 9897 2176 12038
rect 2134 9888 2190 9897
rect 2134 9823 2190 9832
rect 2134 9752 2190 9761
rect 2134 9687 2190 9696
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2042 9208 2098 9217
rect 2042 9143 2098 9152
rect 2056 9110 2084 9143
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 2148 8956 2176 9687
rect 2056 8928 2176 8956
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1950 8528 2006 8537
rect 1950 8463 2006 8472
rect 1780 8214 1900 8242
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1674 6624 1730 6633
rect 1674 6559 1730 6568
rect 1400 6326 1452 6332
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1688 6254 1716 6559
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1490 6080 1546 6089
rect 1490 6015 1546 6024
rect 1504 4622 1532 6015
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1124 3120 1176 3126
rect 1124 3062 1176 3068
rect 1412 3058 1440 3703
rect 1688 3233 1716 6190
rect 1780 5642 1808 8214
rect 1964 7886 1992 8463
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 2056 7732 2084 8928
rect 2134 8664 2190 8673
rect 2134 8599 2190 8608
rect 2148 8022 2176 8599
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2134 7848 2190 7857
rect 2134 7783 2190 7792
rect 1964 7704 2084 7732
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 1872 6798 1900 7375
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1872 5846 1900 6122
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1768 4820 1820 4826
rect 1872 4808 1900 5782
rect 1964 5166 1992 7704
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2056 6769 2084 6870
rect 2042 6760 2098 6769
rect 2042 6695 2098 6704
rect 2056 6186 2084 6695
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 2148 5098 2176 7783
rect 2240 6322 2268 14010
rect 2332 14006 2360 15438
rect 2424 14346 2452 16646
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2410 14104 2466 14113
rect 2516 14074 2544 18702
rect 2700 18465 2728 20198
rect 2792 19446 2820 20703
rect 2884 19718 2912 23530
rect 4618 23520 4674 23582
rect 3700 23180 3752 23186
rect 3700 23122 3752 23128
rect 3712 23089 3740 23122
rect 3698 23080 3754 23089
rect 3698 23015 3754 23024
rect 3700 22364 3752 22370
rect 3700 22306 3752 22312
rect 3240 22296 3292 22302
rect 3240 22238 3292 22244
rect 3054 21448 3110 21457
rect 3054 21383 3110 21392
rect 3148 21412 3200 21418
rect 3068 19854 3096 21383
rect 3148 21354 3200 21360
rect 3160 21078 3188 21354
rect 3148 21072 3200 21078
rect 3148 21014 3200 21020
rect 3056 19848 3108 19854
rect 2962 19816 3018 19825
rect 3056 19790 3108 19796
rect 2962 19751 3018 19760
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 2780 19346 2832 19352
rect 2780 19288 2832 19294
rect 2686 18456 2742 18465
rect 2608 18414 2686 18442
rect 2608 15722 2636 18414
rect 2686 18391 2742 18400
rect 2792 18154 2820 19288
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2686 18048 2742 18057
rect 2884 18034 2912 19110
rect 2686 17983 2742 17992
rect 2792 18006 2912 18034
rect 2700 17746 2728 17983
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2700 17338 2728 17682
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2792 16980 2820 18006
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2884 17338 2912 17682
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2884 17134 2912 17274
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2792 16952 2912 16980
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2608 15694 2728 15722
rect 2792 15706 2820 15914
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2608 14822 2636 15574
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14550 2636 14758
rect 2700 14550 2728 15694
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2778 15192 2834 15201
rect 2884 15162 2912 16952
rect 2976 15638 3004 19751
rect 3252 19553 3280 22238
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 3436 21350 3464 21558
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3436 21010 3464 21286
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3436 20602 3464 20946
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3332 20528 3384 20534
rect 3332 20470 3384 20476
rect 3238 19544 3294 19553
rect 3056 19508 3108 19514
rect 3238 19479 3294 19488
rect 3056 19450 3108 19456
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 3068 15586 3096 19450
rect 3146 19136 3202 19145
rect 3146 19071 3202 19080
rect 3160 17814 3188 19071
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3252 18358 3280 18770
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3344 18290 3372 20470
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3436 19718 3464 20334
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 18426 3464 19654
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 3148 17808 3200 17814
rect 3148 17750 3200 17756
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 15881 3188 17614
rect 3252 17542 3280 18090
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3344 16658 3372 17750
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 16250 3372 16594
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 3332 15972 3384 15978
rect 3146 15872 3202 15881
rect 3146 15807 3202 15816
rect 3068 15558 3188 15586
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2778 15127 2834 15136
rect 2872 15156 2924 15162
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2410 14039 2466 14048
rect 2504 14068 2556 14074
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2332 13326 2360 13942
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 9722 2360 13126
rect 2424 12306 2452 14039
rect 2504 14010 2556 14016
rect 2608 13814 2636 14486
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2516 13786 2636 13814
rect 2516 13462 2544 13786
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2332 9110 2360 9658
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2332 7342 2360 8910
rect 2424 8362 2452 12106
rect 2516 11257 2544 13194
rect 2608 11762 2636 13466
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2594 11656 2650 11665
rect 2594 11591 2650 11600
rect 2502 11248 2558 11257
rect 2502 11183 2558 11192
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9654 2544 10406
rect 2608 9674 2636 11591
rect 2700 10810 2728 14282
rect 2792 13870 2820 15127
rect 2872 15098 2924 15104
rect 2976 14532 3004 15438
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 2884 14504 3004 14532
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2884 13410 2912 14504
rect 2962 14240 3018 14249
rect 2962 14175 3018 14184
rect 2792 13382 2912 13410
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2686 10704 2742 10713
rect 2686 10639 2742 10648
rect 2700 10305 2728 10639
rect 2686 10296 2742 10305
rect 2686 10231 2742 10240
rect 2792 10130 2820 13382
rect 2872 13320 2924 13326
rect 2976 13308 3004 14175
rect 2924 13280 3004 13308
rect 2872 13262 2924 13268
rect 2884 12374 2912 13262
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 10169 2912 11494
rect 2870 10160 2926 10169
rect 2780 10124 2832 10130
rect 2870 10095 2926 10104
rect 2780 10066 2832 10072
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2504 9648 2556 9654
rect 2608 9646 2728 9674
rect 2504 9590 2556 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2608 9489 2636 9522
rect 2594 9480 2650 9489
rect 2594 9415 2650 9424
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2424 8022 2452 8298
rect 2516 8129 2544 9318
rect 2608 8401 2636 9415
rect 2700 9042 2728 9646
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2594 8392 2650 8401
rect 2594 8327 2650 8336
rect 2502 8120 2558 8129
rect 2502 8055 2558 8064
rect 2412 8016 2464 8022
rect 2464 7976 2544 8004
rect 2412 7958 2464 7964
rect 2410 7712 2466 7721
rect 2410 7647 2466 7656
rect 2424 7546 2452 7647
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2226 5944 2282 5953
rect 2226 5879 2282 5888
rect 2240 5846 2268 5879
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2136 5092 2188 5098
rect 2136 5034 2188 5040
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1820 4780 1900 4808
rect 1768 4762 1820 4768
rect 1780 3942 1808 4762
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3738 1808 3878
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1674 3224 1730 3233
rect 1674 3159 1730 3168
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1780 2854 1808 3674
rect 1964 3602 1992 4966
rect 2332 4049 2360 7142
rect 2516 7002 2544 7976
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2424 6458 2452 6734
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2608 6390 2636 8327
rect 2700 8265 2728 8978
rect 2686 8256 2742 8265
rect 2686 8191 2742 8200
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2700 7274 2728 7754
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2686 6488 2742 6497
rect 2686 6423 2742 6432
rect 2700 6390 2728 6423
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2686 6080 2742 6089
rect 2686 6015 2742 6024
rect 2700 5778 2728 6015
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2792 5302 2820 9930
rect 2976 9761 3004 12854
rect 2962 9752 3018 9761
rect 3068 9722 3096 15370
rect 3160 15026 3188 15558
rect 3252 15366 3280 15943
rect 3332 15914 3384 15920
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3238 15192 3294 15201
rect 3238 15127 3294 15136
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3160 12850 3188 14010
rect 3252 12850 3280 15127
rect 3344 14793 3372 15914
rect 3330 14784 3386 14793
rect 3330 14719 3386 14728
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3344 13190 3372 14554
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3436 12918 3464 18158
rect 3528 15570 3556 20878
rect 3606 20632 3662 20641
rect 3606 20567 3662 20576
rect 3620 20398 3648 20567
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3712 20262 3740 22306
rect 4068 22160 4120 22166
rect 4908 22137 4936 23582
rect 6288 23582 6514 23610
rect 4068 22102 4120 22108
rect 4894 22128 4950 22137
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 3896 20346 3924 21898
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3988 20874 4016 21422
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 3896 20318 4016 20346
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3700 19984 3752 19990
rect 3700 19926 3752 19932
rect 3608 19780 3660 19786
rect 3608 19722 3660 19728
rect 3620 18902 3648 19722
rect 3712 19242 3740 19926
rect 3700 19236 3752 19242
rect 3700 19178 3752 19184
rect 3804 19122 3832 19994
rect 3896 19514 3924 20198
rect 3988 20097 4016 20318
rect 3974 20088 4030 20097
rect 3974 20023 4030 20032
rect 3988 19990 4016 20023
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3988 19310 4016 19790
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3712 19094 3832 19122
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3608 18896 3660 18902
rect 3608 18838 3660 18844
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3620 16182 3648 18362
rect 3712 18154 3740 19094
rect 3896 19009 3924 19110
rect 3882 19000 3938 19009
rect 3882 18935 3938 18944
rect 3896 18834 3924 18935
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3700 18148 3752 18154
rect 3700 18090 3752 18096
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 3712 16250 3740 17614
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3608 16176 3660 16182
rect 3608 16118 3660 16124
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 14006 3556 14486
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3514 13832 3570 13841
rect 3514 13767 3570 13776
rect 3528 13734 3556 13767
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3620 13308 3648 16118
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15473 3740 15846
rect 3698 15464 3754 15473
rect 3698 15399 3754 15408
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3712 14482 3740 15302
rect 3804 15162 3832 18702
rect 3884 18692 3936 18698
rect 3884 18634 3936 18640
rect 3896 18426 3924 18634
rect 3988 18426 4016 19246
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3896 17882 3924 18362
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3988 17762 4016 18226
rect 4080 17785 4108 22102
rect 4894 22063 4950 22072
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4436 21684 4488 21690
rect 4356 21644 4436 21672
rect 4252 21616 4304 21622
rect 4252 21558 4304 21564
rect 4264 21146 4292 21558
rect 4252 21140 4304 21146
rect 4252 21082 4304 21088
rect 4160 20528 4212 20534
rect 4264 20516 4292 21082
rect 4356 21078 4384 21644
rect 4436 21626 4488 21632
rect 4724 21622 4752 21830
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4344 21072 4396 21078
rect 4620 21072 4672 21078
rect 4344 21014 4396 21020
rect 4434 21040 4490 21049
rect 4620 21014 4672 21020
rect 4434 20975 4490 20984
rect 4448 20942 4476 20975
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4344 20868 4396 20874
rect 4344 20810 4396 20816
rect 4212 20488 4292 20516
rect 4160 20470 4212 20476
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4172 19990 4200 20266
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 4264 19718 4292 20488
rect 4356 19904 4384 20810
rect 4448 20788 4476 20878
rect 4528 20800 4580 20806
rect 4448 20760 4528 20788
rect 4448 20448 4476 20760
rect 4528 20742 4580 20748
rect 4632 20602 4660 21014
rect 4724 20874 4752 21286
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4724 20777 4752 20810
rect 4710 20768 4766 20777
rect 4710 20703 4766 20712
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4620 20460 4672 20466
rect 4448 20420 4620 20448
rect 4620 20402 4672 20408
rect 4710 20088 4766 20097
rect 4710 20023 4766 20032
rect 4528 19916 4580 19922
rect 4356 19876 4528 19904
rect 4528 19858 4580 19864
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4540 19417 4568 19858
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4526 19408 4582 19417
rect 4632 19378 4660 19654
rect 4724 19446 4752 20023
rect 4816 19854 4844 21490
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5092 21146 5120 21286
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5460 20913 5488 21286
rect 5446 20904 5502 20913
rect 5356 20868 5408 20874
rect 5446 20839 5502 20848
rect 5356 20810 5408 20816
rect 5368 20777 5396 20810
rect 5448 20800 5500 20806
rect 5354 20768 5410 20777
rect 4956 20700 5252 20720
rect 5552 20788 5580 21898
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5920 21146 5948 21626
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 5816 21072 5868 21078
rect 5816 21014 5868 21020
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5500 20760 5580 20788
rect 5448 20742 5500 20748
rect 5354 20703 5410 20712
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4908 20262 4936 20402
rect 4988 20324 5040 20330
rect 4988 20266 5040 20272
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 5000 20058 5028 20266
rect 5460 20262 5488 20538
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4816 19514 4844 19790
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 5460 19514 5488 20198
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 4712 19440 4764 19446
rect 5264 19440 5316 19446
rect 4712 19382 4764 19388
rect 4802 19408 4858 19417
rect 4526 19343 4582 19352
rect 4620 19372 4672 19378
rect 5264 19382 5316 19388
rect 4802 19343 4858 19352
rect 4620 19314 4672 19320
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 3896 17734 4016 17762
rect 4066 17776 4122 17785
rect 3896 16674 3924 17734
rect 4066 17711 4122 17720
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3988 16794 4016 17070
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3896 16646 4016 16674
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3804 14618 3832 14962
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3896 14498 3924 15438
rect 3988 15366 4016 16646
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3804 14470 3924 14498
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3712 14249 3740 14282
rect 3698 14240 3754 14249
rect 3698 14175 3754 14184
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3712 13462 3740 13670
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3620 13280 3740 13308
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3422 12744 3478 12753
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3160 12481 3188 12650
rect 3146 12472 3202 12481
rect 3252 12442 3280 12650
rect 3146 12407 3202 12416
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3160 11558 3188 12242
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2962 9687 3018 9696
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3054 9072 3110 9081
rect 3054 9007 3110 9016
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8430 3004 8774
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 6322 2912 8298
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7993 3004 8230
rect 3068 8022 3096 9007
rect 3160 8974 3188 11494
rect 3252 9489 3280 12038
rect 3238 9480 3294 9489
rect 3238 9415 3294 9424
rect 3252 9178 3280 9415
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3238 8936 3294 8945
rect 3238 8871 3294 8880
rect 3252 8838 3280 8871
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3056 8016 3108 8022
rect 2962 7984 3018 7993
rect 3056 7958 3108 7964
rect 2962 7919 3018 7928
rect 3160 7886 3188 8434
rect 3252 8362 3280 8570
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 8265 3280 8298
rect 3238 8256 3294 8265
rect 3238 8191 3294 8200
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7410 3004 7686
rect 3146 7576 3202 7585
rect 3252 7546 3280 7754
rect 3146 7511 3202 7520
rect 3240 7540 3292 7546
rect 3160 7410 3188 7511
rect 3240 7482 3292 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2962 7168 3018 7177
rect 2962 7103 3018 7112
rect 2976 6934 3004 7103
rect 2964 6928 3016 6934
rect 3068 6905 3096 7210
rect 2964 6870 3016 6876
rect 3054 6896 3110 6905
rect 3054 6831 3110 6840
rect 3068 6458 3096 6831
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2870 6216 2926 6225
rect 2870 6151 2926 6160
rect 2884 5710 2912 6151
rect 3160 5846 3188 7346
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6934 3280 7142
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6186 3280 6598
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2516 4078 2544 5102
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4758 2820 4966
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2686 4312 2742 4321
rect 2686 4247 2742 4256
rect 2700 4214 2728 4247
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2504 4072 2556 4078
rect 2318 4040 2374 4049
rect 2504 4014 2556 4020
rect 2318 3975 2374 3984
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 2961 2360 3334
rect 2410 3088 2466 3097
rect 2410 3023 2466 3032
rect 2424 2990 2452 3023
rect 2516 2990 2544 4014
rect 2884 3670 2912 5646
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3068 4146 3096 5306
rect 3160 5234 3188 5646
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2872 3664 2924 3670
rect 2686 3632 2742 3641
rect 2872 3606 2924 3612
rect 2686 3567 2742 3576
rect 2700 3534 2728 3567
rect 2688 3528 2740 3534
rect 2594 3496 2650 3505
rect 2688 3470 2740 3476
rect 2594 3431 2650 3440
rect 2412 2984 2464 2990
rect 2318 2952 2374 2961
rect 2412 2926 2464 2932
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2318 2887 2374 2896
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1780 2582 1808 2790
rect 1768 2576 1820 2582
rect 1768 2518 1820 2524
rect 940 1964 992 1970
rect 940 1906 992 1912
rect 570 1592 626 1601
rect 570 1527 626 1536
rect 294 96 350 105
rect 478 82 534 480
rect 350 54 534 82
rect 294 31 350 40
rect 478 0 534 54
rect 1398 82 1454 480
rect 1780 82 1808 2518
rect 2332 1737 2360 2790
rect 2608 2650 2636 3431
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2792 2582 2820 2790
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 3160 1873 3188 5170
rect 3252 5166 3280 5714
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3344 4078 3372 12718
rect 3422 12679 3478 12688
rect 3436 10554 3464 12679
rect 3528 11558 3556 12786
rect 3620 11694 3648 13126
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3528 11354 3556 11494
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3436 10526 3556 10554
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 9654 3464 10406
rect 3528 10198 3556 10526
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3422 9208 3478 9217
rect 3422 9143 3478 9152
rect 3436 7449 3464 9143
rect 3528 8634 3556 9862
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3436 7177 3464 7375
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3436 6186 3464 6938
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3436 4826 3464 6122
rect 3528 5166 3556 8366
rect 3620 7206 3648 11494
rect 3712 11014 3740 13280
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 10266 3740 10406
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3712 8673 3740 9658
rect 3698 8664 3754 8673
rect 3804 8634 3832 14470
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3896 13569 3924 14282
rect 3882 13560 3938 13569
rect 3882 13495 3938 13504
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3896 12918 3924 13398
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3884 12776 3936 12782
rect 3988 12764 4016 15098
rect 3936 12736 4016 12764
rect 3884 12718 3936 12724
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11558 3924 12038
rect 3988 11898 4016 12582
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4080 11626 4108 17478
rect 4172 17202 4200 19246
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18222 4292 19110
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4356 18601 4384 18838
rect 4448 18834 4476 19246
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4342 18592 4398 18601
rect 4342 18527 4398 18536
rect 4356 18426 4384 18527
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4356 18086 4384 18362
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4342 17776 4398 17785
rect 4342 17711 4398 17720
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4264 17202 4292 17546
rect 4356 17338 4384 17711
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4448 17134 4476 17478
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4250 16960 4306 16969
rect 4250 16895 4306 16904
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16182 4200 16390
rect 4160 16176 4212 16182
rect 4160 16118 4212 16124
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4172 15502 4200 15914
rect 4264 15570 4292 16895
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 12481 4200 15302
rect 4264 15162 4292 15506
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4250 14920 4306 14929
rect 4250 14855 4306 14864
rect 4158 12472 4214 12481
rect 4158 12407 4214 12416
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4172 12238 4200 12310
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4264 12102 4292 14855
rect 4356 13512 4384 17002
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4448 16250 4476 16934
rect 4540 16658 4568 19246
rect 4816 19009 4844 19343
rect 4802 19000 4858 19009
rect 4802 18935 4858 18944
rect 4804 18624 4856 18630
rect 5276 18612 5304 19382
rect 5354 19272 5410 19281
rect 5354 19207 5410 19216
rect 5368 18766 5396 19207
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5552 18630 5580 19994
rect 5540 18624 5592 18630
rect 5276 18584 5396 18612
rect 4804 18566 4856 18572
rect 4710 18456 4766 18465
rect 4710 18391 4766 18400
rect 4724 17882 4752 18391
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4540 16250 4568 16594
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4448 15473 4476 16186
rect 4434 15464 4490 15473
rect 4434 15399 4490 15408
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14278 4476 14758
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4434 14104 4490 14113
rect 4434 14039 4490 14048
rect 4448 14006 4476 14039
rect 4436 14000 4488 14006
rect 4540 13988 4568 16186
rect 4632 16046 4660 17750
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4632 15706 4660 15982
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4724 14414 4752 17206
rect 4816 15502 4844 18566
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 5368 18408 5396 18584
rect 5540 18566 5592 18572
rect 5184 18380 5396 18408
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4908 17746 4936 18294
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4908 17524 4936 17682
rect 5184 17678 5212 18380
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5276 17746 5304 18158
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4883 17496 4936 17524
rect 4883 17320 4911 17496
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 4883 17292 4936 17320
rect 4908 17066 4936 17292
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 4908 16969 4936 17002
rect 5172 16992 5224 16998
rect 4894 16960 4950 16969
rect 5276 16969 5304 17002
rect 5172 16934 5224 16940
rect 5262 16960 5318 16969
rect 4894 16895 4950 16904
rect 5184 16368 5212 16934
rect 5262 16895 5318 16904
rect 5368 16658 5396 18226
rect 5460 16998 5488 18226
rect 5644 17762 5672 20810
rect 5736 20602 5764 20878
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5736 19718 5764 20266
rect 5828 19990 5856 21014
rect 5920 20942 5948 21082
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5908 20528 5960 20534
rect 5908 20470 5960 20476
rect 5920 20058 5948 20470
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5736 18970 5764 19110
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5828 18873 5856 19314
rect 5920 19242 5948 19994
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 5908 18896 5960 18902
rect 5814 18864 5870 18873
rect 5908 18838 5960 18844
rect 5814 18799 5870 18808
rect 5920 18426 5948 18838
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5552 17734 5672 17762
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 4986 16144 5042 16153
rect 4986 16079 5042 16088
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4908 15348 4936 15574
rect 5000 15502 5028 16079
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4816 15320 4936 15348
rect 4816 14464 4844 15320
rect 5092 15280 5120 15846
rect 5184 15638 5212 16272
rect 5368 15706 5396 16594
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5354 15464 5410 15473
rect 5354 15399 5410 15408
rect 5368 15366 5396 15399
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 5092 14890 5120 15184
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5078 14648 5134 14657
rect 4988 14612 5040 14618
rect 5040 14592 5078 14600
rect 5184 14618 5212 15030
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 14618 5304 14826
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5040 14583 5134 14592
rect 5172 14612 5224 14618
rect 5040 14572 5120 14583
rect 4988 14554 5040 14560
rect 5172 14554 5224 14560
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 4816 14436 5028 14464
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4436 13942 4488 13948
rect 4534 13960 4568 13988
rect 4534 13818 4562 13960
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4534 13790 4568 13818
rect 4356 13484 4476 13512
rect 4448 13394 4476 13484
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4356 12782 4384 13330
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12986 4476 13126
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4540 12866 4568 13790
rect 4632 13433 4660 13874
rect 4618 13424 4674 13433
rect 4618 13359 4674 13368
rect 4724 13297 4752 14214
rect 4816 14006 4844 14282
rect 5000 14260 5028 14436
rect 4883 14232 5028 14260
rect 4883 14056 4911 14232
rect 5184 14192 5212 14554
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 4883 14028 5120 14056
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4986 13968 5042 13977
rect 4986 13903 5042 13912
rect 4896 13864 4948 13870
rect 4816 13824 4896 13852
rect 4710 13288 4766 13297
rect 4620 13252 4672 13258
rect 4710 13223 4766 13232
rect 4620 13194 4672 13200
rect 4448 12838 4568 12866
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 12096 4304 12102
rect 4356 12073 4384 12174
rect 4252 12038 4304 12044
rect 4342 12064 4398 12073
rect 4342 11999 4398 12008
rect 4342 11928 4398 11937
rect 4160 11892 4212 11898
rect 4342 11863 4398 11872
rect 4160 11834 4212 11840
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3896 10606 3924 11290
rect 4080 11286 4108 11562
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 10742 4016 10775
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3974 10568 4030 10577
rect 3974 10503 4030 10512
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10062 3924 10406
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3882 8800 3938 8809
rect 3882 8735 3938 8744
rect 3698 8599 3754 8608
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3698 8120 3754 8129
rect 3698 8055 3754 8064
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3712 5642 3740 8055
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 4593 3556 4626
rect 3514 4584 3570 4593
rect 3514 4519 3570 4528
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3332 4072 3384 4078
rect 3238 4040 3294 4049
rect 3332 4014 3384 4020
rect 3238 3975 3294 3984
rect 3252 3942 3280 3975
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3240 3732 3292 3738
rect 3344 3720 3372 3878
rect 3436 3738 3464 4111
rect 3292 3692 3372 3720
rect 3424 3732 3476 3738
rect 3240 3674 3292 3680
rect 3424 3674 3476 3680
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3146 1864 3202 1873
rect 3146 1799 3202 1808
rect 2318 1728 2374 1737
rect 2318 1663 2374 1672
rect 3344 1193 3372 2790
rect 3528 2514 3556 4519
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3620 2417 3648 5034
rect 3712 4010 3740 5578
rect 3804 4154 3832 8230
rect 3896 6866 3924 8735
rect 3988 7410 4016 10503
rect 4080 9994 4108 11222
rect 4172 10996 4200 11834
rect 4250 11792 4306 11801
rect 4250 11727 4306 11736
rect 4264 11150 4292 11727
rect 4356 11694 4384 11863
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4356 11354 4384 11630
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4172 10968 4292 10996
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4172 10266 4200 10746
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4172 9897 4200 10066
rect 4158 9888 4214 9897
rect 4158 9823 4214 9832
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4080 9602 4108 9658
rect 4172 9602 4200 9823
rect 4080 9574 4200 9602
rect 4158 9480 4214 9489
rect 4068 9444 4120 9450
rect 4158 9415 4214 9424
rect 4068 9386 4120 9392
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 7002 4016 7103
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3974 6760 4030 6769
rect 3974 6695 4030 6704
rect 3988 6662 4016 6695
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3896 6225 3924 6598
rect 3974 6488 4030 6497
rect 3974 6423 4030 6432
rect 3988 6390 4016 6423
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3882 6216 3938 6225
rect 3882 6151 3938 6160
rect 4080 5914 4108 9386
rect 4172 8362 4200 9415
rect 4264 8809 4292 10968
rect 4356 10810 4384 11154
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4356 10470 4384 10746
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4342 10296 4398 10305
rect 4342 10231 4398 10240
rect 4356 9738 4384 10231
rect 4448 9897 4476 12838
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11937 4568 12038
rect 4526 11928 4582 11937
rect 4526 11863 4582 11872
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4540 11082 4568 11698
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4526 10704 4582 10713
rect 4526 10639 4582 10648
rect 4540 10606 4568 10639
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4632 10266 4660 13194
rect 4712 13184 4764 13190
rect 4816 13172 4844 13824
rect 4896 13806 4948 13812
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4908 13172 4936 13398
rect 5000 13258 5028 13903
rect 5092 13802 5120 14028
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 4764 13144 4844 13172
rect 4883 13144 4936 13172
rect 5184 13172 5212 14096
rect 5368 13569 5396 14758
rect 5460 14550 5488 16594
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 13938 5488 14350
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5354 13560 5410 13569
rect 5354 13495 5410 13504
rect 5184 13144 5396 13172
rect 4712 13126 4764 13132
rect 4724 11150 4752 13126
rect 4883 12968 4911 13144
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 4883 12940 4936 12968
rect 4802 12880 4858 12889
rect 4802 12815 4858 12824
rect 4816 12714 4844 12815
rect 4908 12714 4936 12940
rect 4986 12744 5042 12753
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4896 12708 4948 12714
rect 4986 12679 5042 12688
rect 4896 12650 4948 12656
rect 4816 12306 4844 12650
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4908 12238 4936 12650
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4816 11558 4844 12106
rect 5000 12084 5028 12679
rect 4883 12056 5028 12084
rect 4883 11880 4911 12056
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 4883 11852 5028 11880
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4804 11552 4856 11558
rect 4908 11529 4936 11562
rect 4804 11494 4856 11500
rect 4894 11520 4950 11529
rect 4894 11455 4950 11464
rect 4908 11354 4936 11455
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4710 10568 4766 10577
rect 4710 10503 4766 10512
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4434 9888 4490 9897
rect 4434 9823 4490 9832
rect 4356 9722 4476 9738
rect 4356 9716 4488 9722
rect 4356 9710 4436 9716
rect 4436 9658 4488 9664
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4250 8800 4306 8809
rect 4250 8735 4306 8744
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4264 8362 4292 8434
rect 4356 8430 4384 9590
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4448 9450 4476 9522
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4448 9217 4476 9386
rect 4434 9208 4490 9217
rect 4434 9143 4436 9152
rect 4488 9143 4490 9152
rect 4436 9114 4488 9120
rect 4448 9083 4476 9114
rect 4434 8664 4490 8673
rect 4434 8599 4490 8608
rect 4448 8498 4476 8599
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7478 4200 7890
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4158 7168 4214 7177
rect 4158 7103 4214 7112
rect 4172 6662 4200 7103
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4158 6352 4214 6361
rect 4158 6287 4214 6296
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3882 5808 3938 5817
rect 3882 5743 3938 5752
rect 4068 5772 4120 5778
rect 3896 4758 3924 5743
rect 4068 5714 4120 5720
rect 4080 5681 4108 5714
rect 4066 5672 4122 5681
rect 3976 5636 4028 5642
rect 4066 5607 4122 5616
rect 3976 5578 4028 5584
rect 3988 5166 4016 5578
rect 4172 5522 4200 6287
rect 4080 5494 4200 5522
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3974 4720 4030 4729
rect 3974 4655 4030 4664
rect 3988 4622 4016 4655
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3804 4126 3924 4154
rect 3896 4078 3924 4126
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 4080 3602 4108 5494
rect 4158 5128 4214 5137
rect 4158 5063 4214 5072
rect 4172 4185 4200 5063
rect 4264 4554 4292 8191
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4356 6934 4384 7414
rect 4448 7206 4476 7686
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4448 6322 4476 7142
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4434 6216 4490 6225
rect 4356 6186 4434 6202
rect 4344 6180 4434 6186
rect 4396 6174 4434 6180
rect 4434 6151 4490 6160
rect 4344 6122 4396 6128
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5846 4476 6054
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4356 5030 4384 5782
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4356 4214 4384 4762
rect 4448 4729 4476 5102
rect 4434 4720 4490 4729
rect 4540 4690 4568 10134
rect 4632 9897 4660 10202
rect 4724 10169 4752 10503
rect 4816 10266 4844 11018
rect 5000 10996 5028 11852
rect 5262 11520 5318 11529
rect 5262 11455 5318 11464
rect 5276 11218 5304 11455
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 4883 10968 5028 10996
rect 4883 10792 4911 10968
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 4883 10764 4936 10792
rect 4908 10577 4936 10764
rect 5080 10600 5132 10606
rect 4894 10568 4950 10577
rect 5080 10542 5132 10548
rect 4894 10503 4950 10512
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4710 10160 4766 10169
rect 4710 10095 4766 10104
rect 4618 9888 4674 9897
rect 4816 9874 4844 10202
rect 4908 10033 4936 10503
rect 4894 10024 4950 10033
rect 5092 9994 5120 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10198 5212 10406
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5276 10062 5304 11018
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4894 9959 4950 9968
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4618 9823 4674 9832
rect 4770 9846 4844 9874
rect 4620 9716 4672 9722
rect 4770 9674 4798 9846
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 4620 9658 4672 9664
rect 4632 6118 4660 9658
rect 4724 9654 4798 9674
rect 4712 9648 4798 9654
rect 4764 9646 4798 9648
rect 5264 9648 5316 9654
rect 4712 9590 4764 9596
rect 4986 9616 5042 9625
rect 4986 9551 5042 9560
rect 5170 9616 5226 9625
rect 5264 9590 5316 9596
rect 5170 9551 5226 9560
rect 4894 9480 4950 9489
rect 4804 9444 4856 9450
rect 4894 9415 4950 9424
rect 4804 9386 4856 9392
rect 4816 8906 4844 9386
rect 4908 9110 4936 9415
rect 5000 9217 5028 9551
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4986 9208 5042 9217
rect 4986 9143 5042 9152
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 5000 8974 5028 9046
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 8566 4752 8774
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 6662 4752 8230
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4724 5710 4752 6598
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4710 5536 4766 5545
rect 4632 5098 4660 5510
rect 4710 5471 4766 5480
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4724 4978 4752 5471
rect 4816 5250 4844 8842
rect 5092 8752 5120 9454
rect 5184 8752 5212 9551
rect 5276 9081 5304 9590
rect 5262 9072 5318 9081
rect 5262 9007 5318 9016
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5092 8430 5120 8656
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4908 7732 4936 7958
rect 4883 7704 4936 7732
rect 4883 7528 4911 7704
rect 5092 7664 5120 8366
rect 5184 8294 5212 8656
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5368 7954 5396 13144
rect 5460 13025 5488 13670
rect 5446 13016 5502 13025
rect 5446 12951 5502 12960
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5460 11694 5488 12854
rect 5552 12238 5580 17734
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5644 13462 5672 17614
rect 5816 17604 5868 17610
rect 5816 17546 5868 17552
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5736 17134 5764 17478
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5736 16454 5764 17070
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 14006 5764 16390
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5644 12850 5672 13398
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5630 12744 5686 12753
rect 5736 12714 5764 13738
rect 5828 13161 5856 17546
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5920 14482 5948 17002
rect 6012 16697 6040 21286
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 6104 16833 6132 19994
rect 6196 19378 6224 20946
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6288 19145 6316 23582
rect 6458 23520 6514 23582
rect 8298 23610 8354 24000
rect 10138 23610 10194 24000
rect 11978 23610 12034 24000
rect 13818 23610 13874 24000
rect 15658 23610 15714 24000
rect 17498 23610 17554 24000
rect 8298 23582 8616 23610
rect 8298 23520 8354 23582
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 6642 22808 6698 22817
rect 6642 22743 6698 22752
rect 6656 21690 6684 22743
rect 7010 21720 7066 21729
rect 6644 21684 6696 21690
rect 7010 21655 7066 21664
rect 6644 21626 6696 21632
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6380 20330 6408 20946
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6550 20224 6606 20233
rect 6550 20159 6606 20168
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6380 19718 6408 19858
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6274 19136 6330 19145
rect 6274 19071 6330 19080
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6196 18698 6224 18770
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6196 18426 6224 18634
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6380 17762 6408 19450
rect 6472 19446 6500 19994
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6472 18465 6500 18702
rect 6564 18698 6592 20159
rect 6656 19310 6684 21626
rect 7024 21554 7052 21655
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6458 18456 6514 18465
rect 6458 18391 6514 18400
rect 6196 17734 6408 17762
rect 6196 17338 6224 17734
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6090 16824 6146 16833
rect 6090 16759 6146 16768
rect 6092 16720 6144 16726
rect 5998 16688 6054 16697
rect 6196 16697 6224 17138
rect 6092 16662 6144 16668
rect 6182 16688 6238 16697
rect 5998 16623 6054 16632
rect 6012 16250 6040 16623
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6104 16046 6132 16662
rect 6182 16623 6238 16632
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 6012 14822 6040 15574
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5814 13152 5870 13161
rect 5814 13087 5870 13096
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5630 12679 5686 12688
rect 5724 12708 5776 12714
rect 5644 12646 5672 12679
rect 5724 12650 5776 12656
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5630 12472 5686 12481
rect 5630 12407 5686 12416
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 10606 5488 11630
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10266 5488 10406
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5460 9178 5488 9998
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5354 7848 5410 7857
rect 5354 7783 5410 7792
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 4883 7500 5028 7528
rect 5000 7002 5028 7500
rect 5092 7392 5120 7568
rect 5368 7546 5396 7783
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5092 7364 5212 7392
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4988 6792 5040 6798
rect 4908 6769 4988 6780
rect 4894 6760 4988 6769
rect 4950 6752 4988 6760
rect 4988 6734 5040 6740
rect 5092 6730 5120 7210
rect 5184 6769 5212 7364
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5170 6760 5226 6769
rect 4894 6695 4950 6704
rect 5080 6724 5132 6730
rect 5170 6695 5226 6704
rect 5080 6666 5132 6672
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5092 5488 5120 6326
rect 5170 5808 5226 5817
rect 5170 5743 5226 5752
rect 5184 5710 5212 5743
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 5092 5302 5120 5392
rect 5080 5296 5132 5302
rect 4816 5222 4936 5250
rect 5080 5238 5132 5244
rect 5262 5264 5318 5273
rect 4632 4950 4752 4978
rect 4632 4758 4660 4950
rect 4710 4856 4766 4865
rect 4710 4791 4766 4800
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4434 4655 4490 4664
rect 4528 4684 4580 4690
rect 4448 4622 4476 4655
rect 4528 4626 4580 4632
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4344 4208 4396 4214
rect 4158 4176 4214 4185
rect 4448 4185 4476 4422
rect 4344 4150 4396 4156
rect 4434 4176 4490 4185
rect 4158 4111 4214 4120
rect 4434 4111 4490 4120
rect 4540 4078 4568 4422
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4158 3632 4214 3641
rect 4068 3596 4120 3602
rect 4158 3567 4214 3576
rect 4068 3538 4120 3544
rect 4172 3466 4200 3567
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3698 3088 3754 3097
rect 3698 3023 3754 3032
rect 3606 2408 3662 2417
rect 3606 2343 3662 2352
rect 3330 1184 3386 1193
rect 3330 1119 3386 1128
rect 1398 54 1808 82
rect 2410 128 2466 480
rect 2410 76 2412 128
rect 2464 76 2466 128
rect 1398 0 1454 54
rect 2410 0 2466 76
rect 3422 82 3478 480
rect 3712 82 3740 3023
rect 4540 2922 4568 3674
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 3988 2582 4016 2858
rect 4066 2680 4122 2689
rect 4066 2615 4122 2624
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 4080 2514 4108 2615
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 4264 1834 4292 2314
rect 4252 1828 4304 1834
rect 4252 1770 4304 1776
rect 3422 54 3740 82
rect 4434 82 4490 480
rect 4632 241 4660 4558
rect 4724 4486 4752 4791
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4816 3942 4844 4694
rect 4908 4672 4936 5222
rect 5262 5199 5318 5208
rect 5276 5098 5304 5199
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5368 4826 5396 6870
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5172 4684 5224 4690
rect 4908 4644 5172 4672
rect 5172 4626 5224 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3670 5304 3878
rect 5368 3738 5396 4626
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 4802 2544 4858 2553
rect 4802 2479 4858 2488
rect 4816 2038 4844 2479
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 5368 1970 5396 2790
rect 5460 2310 5488 8978
rect 5552 7274 5580 12038
rect 5644 9926 5672 12407
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5736 11200 5764 12174
rect 5828 11937 5856 12922
rect 5814 11928 5870 11937
rect 5814 11863 5870 11872
rect 5920 11558 5948 14282
rect 6012 13530 6040 14758
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12374 6040 12582
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 5736 11172 5856 11200
rect 5722 11112 5778 11121
rect 5722 11047 5778 11056
rect 5736 11014 5764 11047
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5828 10130 5856 11172
rect 5920 10810 5948 11222
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5906 10432 5962 10441
rect 5906 10367 5962 10376
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5722 9888 5778 9897
rect 5644 9586 5672 9862
rect 5722 9823 5778 9832
rect 5736 9722 5764 9823
rect 5814 9752 5870 9761
rect 5724 9716 5776 9722
rect 5814 9687 5870 9696
rect 5724 9658 5776 9664
rect 5632 9580 5684 9586
rect 5684 9540 5764 9568
rect 5632 9522 5684 9528
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5644 8362 5672 9114
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5630 7848 5686 7857
rect 5630 7783 5686 7792
rect 5644 7750 5672 7783
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5552 5846 5580 6938
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5644 6458 5672 6666
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5644 6254 5672 6394
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5552 4690 5580 5782
rect 5644 5302 5672 6054
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5644 4826 5672 5034
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5632 4616 5684 4622
rect 5736 4604 5764 9540
rect 5828 6390 5856 9687
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5814 6216 5870 6225
rect 5814 6151 5870 6160
rect 5684 4576 5764 4604
rect 5632 4558 5684 4564
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5538 4040 5594 4049
rect 5538 3975 5594 3984
rect 5552 2825 5580 3975
rect 5538 2816 5594 2825
rect 5538 2751 5594 2760
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 4712 1896 4764 1902
rect 4712 1838 4764 1844
rect 4618 232 4674 241
rect 4618 167 4674 176
rect 4724 82 4752 1838
rect 4434 54 4752 82
rect 5446 82 5502 480
rect 5552 82 5580 2246
rect 5644 785 5672 4422
rect 5722 3632 5778 3641
rect 5828 3602 5856 6151
rect 5920 4842 5948 10367
rect 6012 9042 6040 12310
rect 6104 10266 6132 15846
rect 6196 15570 6224 16390
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6288 15434 6316 17614
rect 6564 17456 6592 18634
rect 6656 18465 6684 19110
rect 6642 18456 6698 18465
rect 6642 18391 6698 18400
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6380 17428 6592 17456
rect 6380 16130 6408 17428
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6472 16658 6500 17274
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6550 16552 6606 16561
rect 6550 16487 6606 16496
rect 6564 16250 6592 16487
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6380 16102 6592 16130
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6196 14006 6224 15098
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14618 6316 14894
rect 6380 14634 6408 15914
rect 6564 15620 6592 16102
rect 6656 15881 6684 17818
rect 6642 15872 6698 15881
rect 6642 15807 6698 15816
rect 6472 15592 6592 15620
rect 6644 15632 6696 15638
rect 6472 15162 6500 15592
rect 6564 15580 6644 15586
rect 6564 15574 6696 15580
rect 6564 15558 6684 15574
rect 6564 15502 6592 15558
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6564 14890 6592 15302
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6564 14793 6592 14826
rect 6550 14784 6606 14793
rect 6550 14719 6606 14728
rect 6276 14612 6328 14618
rect 6380 14606 6592 14634
rect 6276 14554 6328 14560
rect 6564 14464 6592 14606
rect 6472 14436 6592 14464
rect 6368 14272 6420 14278
rect 6472 14260 6500 14436
rect 6420 14232 6500 14260
rect 6552 14272 6604 14278
rect 6368 14214 6420 14220
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6472 13814 6500 14232
rect 6550 14240 6552 14249
rect 6604 14240 6606 14249
rect 6550 14175 6606 14184
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6380 13786 6500 13814
rect 6182 12880 6238 12889
rect 6182 12815 6238 12824
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6090 10160 6146 10169
rect 6090 10095 6146 10104
rect 6104 9761 6132 10095
rect 6090 9752 6146 9761
rect 6090 9687 6146 9696
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5998 8936 6054 8945
rect 5998 8871 6054 8880
rect 6012 7818 6040 8871
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6104 7460 6132 9454
rect 6196 9110 6224 12815
rect 6288 12374 6316 13738
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 12073 6316 12174
rect 6274 12064 6330 12073
rect 6274 11999 6330 12008
rect 6380 11914 6408 13786
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 13326 6500 13670
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6564 12850 6592 14175
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6288 11898 6408 11914
rect 6276 11892 6408 11898
rect 6328 11886 6408 11892
rect 6276 11834 6328 11840
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 9518 6316 11494
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6288 8906 6316 9318
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6274 8800 6330 8809
rect 6274 8735 6330 8744
rect 6182 7984 6238 7993
rect 6182 7919 6238 7928
rect 6196 7585 6224 7919
rect 6288 7886 6316 8735
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6104 7432 6316 7460
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6092 7200 6144 7206
rect 5998 7168 6054 7177
rect 6092 7142 6144 7148
rect 5998 7103 6054 7112
rect 6012 6934 6040 7103
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6104 6662 6132 7142
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6012 5846 6040 6394
rect 6104 6118 6132 6598
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6012 5642 6040 5782
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 5001 6040 5034
rect 5998 4992 6054 5001
rect 5998 4927 6054 4936
rect 5920 4814 6040 4842
rect 5906 4448 5962 4457
rect 5906 4383 5962 4392
rect 5920 4078 5948 4383
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5920 3641 5948 3878
rect 5906 3632 5962 3641
rect 5722 3567 5778 3576
rect 5816 3596 5868 3602
rect 5736 3534 5764 3567
rect 5906 3567 5962 3576
rect 5816 3538 5868 3544
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 6012 2922 6040 4814
rect 6104 4468 6132 6054
rect 6196 5681 6224 7278
rect 6288 6458 6316 7432
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6274 6352 6330 6361
rect 6274 6287 6330 6296
rect 6288 5846 6316 6287
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6182 5672 6238 5681
rect 6182 5607 6238 5616
rect 6276 5636 6328 5642
rect 6196 4622 6224 5607
rect 6276 5578 6328 5584
rect 6288 4622 6316 5578
rect 6380 5574 6408 11766
rect 6472 11762 6500 12378
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6564 11286 6592 12582
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6380 4826 6408 5034
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6104 4440 6316 4468
rect 6090 4312 6146 4321
rect 6090 4247 6146 4256
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5736 2582 5764 2858
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 6104 2514 6132 4247
rect 6288 4154 6316 4440
rect 6288 4126 6408 4154
rect 6184 4072 6236 4078
rect 6380 4060 6408 4126
rect 6236 4032 6408 4060
rect 6184 4014 6236 4020
rect 6196 3652 6224 4014
rect 6368 3664 6420 3670
rect 6196 3624 6316 3652
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 5630 776 5686 785
rect 5630 711 5686 720
rect 5446 54 5580 82
rect 6196 82 6224 2586
rect 6288 2106 6316 3624
rect 6368 3606 6420 3612
rect 6380 3505 6408 3606
rect 6366 3496 6422 3505
rect 6472 3482 6500 9862
rect 6564 8022 6592 10202
rect 6656 10169 6684 15438
rect 6748 12102 6776 20878
rect 6840 20534 6868 21286
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 7010 20360 7066 20369
rect 6840 20058 6868 20334
rect 7010 20295 7066 20304
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6826 19680 6882 19689
rect 6932 19666 6960 20198
rect 6882 19638 6960 19666
rect 6826 19615 6882 19624
rect 7024 19446 7052 20295
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6932 18034 6960 19246
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18154 7052 18566
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6932 18006 7052 18034
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6840 17746 6868 17818
rect 7024 17785 7052 18006
rect 7010 17776 7066 17785
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6920 17740 6972 17746
rect 7010 17711 7066 17720
rect 6920 17682 6972 17688
rect 6840 17270 6868 17682
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6828 16992 6880 16998
rect 6932 16980 6960 17682
rect 7024 17202 7052 17711
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 6880 16952 6960 16980
rect 6828 16934 6880 16940
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16584 6880 16590
rect 6932 16561 6960 16662
rect 6828 16526 6880 16532
rect 6918 16552 6974 16561
rect 6840 16182 6868 16526
rect 6918 16487 6974 16496
rect 7024 16454 7052 17002
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16289 7052 16390
rect 7010 16280 7066 16289
rect 7010 16215 7066 16224
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6826 15736 6882 15745
rect 6826 15671 6882 15680
rect 6840 15094 6868 15671
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14278 6868 14758
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 12986 6868 14214
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11762 6776 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 10713 6776 11018
rect 6734 10704 6790 10713
rect 6734 10639 6790 10648
rect 6734 10432 6790 10441
rect 6734 10367 6790 10376
rect 6642 10160 6698 10169
rect 6642 10095 6698 10104
rect 6748 10112 6776 10367
rect 6840 10112 6868 12650
rect 6932 12238 6960 15846
rect 7024 14074 7052 15846
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7010 13968 7066 13977
rect 7010 13903 7066 13912
rect 7024 13802 7052 13903
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12918 7052 13330
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6932 10418 6960 11834
rect 7024 10538 7052 12310
rect 7116 11200 7144 21354
rect 7208 21078 7236 22986
rect 7654 22944 7710 22953
rect 7654 22879 7710 22888
rect 7838 22944 7894 22953
rect 7838 22879 7894 22888
rect 7668 22846 7696 22879
rect 7564 22840 7616 22846
rect 7564 22782 7616 22788
rect 7656 22840 7708 22846
rect 7656 22782 7708 22788
rect 7576 22681 7604 22782
rect 7378 22672 7434 22681
rect 7378 22607 7434 22616
rect 7562 22672 7618 22681
rect 7562 22607 7618 22616
rect 7392 22001 7420 22607
rect 7852 22370 7880 22879
rect 8206 22536 8262 22545
rect 8206 22471 8262 22480
rect 7840 22364 7892 22370
rect 7840 22306 7892 22312
rect 8024 22364 8076 22370
rect 8024 22306 8076 22312
rect 7378 21992 7434 22001
rect 7378 21927 7434 21936
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 7300 21486 7328 21558
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7208 19310 7236 20742
rect 7300 20602 7328 21422
rect 7654 21176 7710 21185
rect 7852 21146 7880 21422
rect 7654 21111 7710 21120
rect 7840 21140 7892 21146
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7378 20632 7434 20641
rect 7288 20596 7340 20602
rect 7378 20567 7434 20576
rect 7288 20538 7340 20544
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7300 19990 7328 20266
rect 7288 19984 7340 19990
rect 7288 19926 7340 19932
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 18834 7236 19110
rect 7300 18970 7328 19654
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7392 18612 7420 20567
rect 7484 19514 7512 20946
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 19990 7604 20878
rect 7668 20874 7696 21111
rect 7840 21082 7892 21088
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7852 20398 7880 21082
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 20097 7880 20334
rect 7944 20330 7972 20946
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 7838 20088 7894 20097
rect 7838 20023 7894 20032
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7300 18584 7420 18612
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7208 17649 7236 18158
rect 7194 17640 7250 17649
rect 7194 17575 7250 17584
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7208 11354 7236 16934
rect 7300 16726 7328 18584
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17785 7420 18226
rect 7484 17882 7512 19450
rect 7576 18902 7604 19926
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7668 18834 7696 19790
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 18426 7604 18702
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7576 18290 7604 18362
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7378 17776 7434 17785
rect 7378 17711 7434 17720
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 7286 16416 7342 16425
rect 7286 16351 7342 16360
rect 7300 15910 7328 16351
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 14521 7328 15302
rect 7286 14512 7342 14521
rect 7286 14447 7342 14456
rect 7392 14396 7420 17138
rect 7484 16969 7512 17206
rect 7470 16960 7526 16969
rect 7470 16895 7526 16904
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 15337 7512 16526
rect 7470 15328 7526 15337
rect 7470 15263 7526 15272
rect 7470 15192 7526 15201
rect 7470 15127 7526 15136
rect 7300 14368 7420 14396
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7116 11172 7236 11200
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6932 10390 7052 10418
rect 6748 10084 6868 10112
rect 6840 10010 6868 10084
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6656 9982 6868 10010
rect 6656 9926 6684 9982
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6656 8974 6684 9658
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6656 7936 6684 8774
rect 6564 7908 6684 7936
rect 6564 7857 6592 7908
rect 6748 7886 6776 9862
rect 6840 9110 6868 9982
rect 6932 9450 6960 10066
rect 7024 9926 7052 10390
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7116 9738 7144 10950
rect 7024 9710 7144 9738
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6828 9104 6880 9110
rect 7024 9058 7052 9710
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7116 9450 7144 9590
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 6828 9046 6880 9052
rect 6907 9030 7052 9058
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6907 8922 6935 9030
rect 6736 7880 6788 7886
rect 6550 7848 6606 7857
rect 6606 7806 6684 7834
rect 6736 7822 6788 7828
rect 6550 7783 6606 7792
rect 6564 7177 6592 7783
rect 6656 7478 6684 7806
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6550 7168 6606 7177
rect 6550 7103 6606 7112
rect 6656 6934 6684 7414
rect 6748 7410 6776 7822
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6840 7002 6868 8910
rect 6907 8894 6960 8922
rect 6932 8378 6960 8894
rect 6932 8350 7144 8378
rect 7116 8294 7144 8350
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6932 7818 6960 8026
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6644 6928 6696 6934
rect 6696 6888 6776 6916
rect 6644 6870 6696 6876
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6642 5808 6698 5817
rect 6564 4078 6592 5782
rect 6642 5743 6698 5752
rect 6656 5098 6684 5743
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6748 5030 6776 6888
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6642 4856 6698 4865
rect 6642 4791 6698 4800
rect 6656 4758 6684 4791
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6734 4312 6790 4321
rect 6734 4247 6790 4256
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6748 4010 6776 4247
rect 6840 4078 6868 6666
rect 6932 5896 6960 7482
rect 7024 7041 7052 8230
rect 7102 7984 7158 7993
rect 7102 7919 7158 7928
rect 7010 7032 7066 7041
rect 7010 6967 7066 6976
rect 7116 6458 7144 7919
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7208 6390 7236 11172
rect 7300 8090 7328 14368
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7392 13394 7420 13670
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7392 12850 7420 13330
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 10130 7420 12582
rect 7484 12306 7512 15127
rect 7576 13938 7604 18090
rect 7668 17542 7696 18770
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7668 14414 7696 16390
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7668 13814 7696 14350
rect 7760 13814 7788 19926
rect 7852 18902 7880 20023
rect 8036 19334 8064 22306
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8128 19854 8156 21286
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 7932 19304 7984 19310
rect 8036 19306 8156 19334
rect 8128 19258 8156 19306
rect 8220 19258 8248 22471
rect 8588 22420 8616 23582
rect 10138 23582 10456 23610
rect 10138 23520 10194 23582
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8680 22545 8708 22714
rect 8666 22536 8722 22545
rect 8666 22471 8722 22480
rect 9220 22432 9272 22438
rect 8588 22392 8708 22420
rect 8298 22128 8354 22137
rect 8298 22063 8354 22072
rect 8312 20534 8340 22063
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8390 20768 8446 20777
rect 8390 20703 8446 20712
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8312 20398 8340 20470
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8404 19922 8432 20703
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8312 19258 8340 19858
rect 7984 19252 8340 19258
rect 7932 19246 8340 19252
rect 7944 19230 8340 19246
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7838 18456 7894 18465
rect 7838 18391 7894 18400
rect 7852 18222 7880 18391
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7840 18080 7892 18086
rect 7838 18048 7840 18057
rect 7892 18048 7894 18057
rect 7838 17983 7894 17992
rect 7852 17134 7880 17983
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7852 15910 7880 16662
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7852 15026 7880 15438
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7852 14793 7880 14826
rect 7838 14784 7894 14793
rect 7838 14719 7894 14728
rect 7838 14648 7894 14657
rect 7838 14583 7894 14592
rect 7852 13938 7880 14583
rect 7944 14414 7972 18702
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7564 13796 7616 13802
rect 7668 13786 7880 13814
rect 7564 13738 7616 13744
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7484 9654 7512 12242
rect 7576 10674 7604 13738
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13190 7696 13670
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7668 10985 7696 12854
rect 7760 12714 7788 13786
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 12102 7788 12310
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11898 7788 12038
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7746 11792 7802 11801
rect 7746 11727 7802 11736
rect 7760 11354 7788 11727
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7852 11268 7880 13786
rect 7944 11830 7972 14214
rect 8036 13433 8064 19110
rect 8128 17338 8156 19230
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8128 15978 8156 16662
rect 8220 16289 8248 19230
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18154 8340 19110
rect 8404 18970 8432 19858
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 17882 8340 18090
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8298 17776 8354 17785
rect 8298 17711 8354 17720
rect 8312 17338 8340 17711
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8206 16280 8262 16289
rect 8206 16215 8262 16224
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 13569 8156 15302
rect 8220 14618 8248 16050
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 13734 8248 14350
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8114 13560 8170 13569
rect 8114 13495 8170 13504
rect 8022 13424 8078 13433
rect 8022 13359 8078 13368
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12442 8064 13126
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 8036 11336 8064 12378
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11898 8156 12174
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8036 11308 8156 11336
rect 7852 11240 8064 11268
rect 7748 11144 7800 11150
rect 7800 11104 7880 11132
rect 7748 11086 7800 11092
rect 7654 10976 7710 10985
rect 7654 10911 7710 10920
rect 7654 10840 7710 10849
rect 7654 10775 7710 10784
rect 7748 10804 7800 10810
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 9648 7524 9654
rect 7392 9608 7472 9636
rect 7392 8498 7420 9608
rect 7472 9590 7524 9596
rect 7576 9110 7604 10610
rect 7564 9104 7616 9110
rect 7470 9072 7526 9081
rect 7564 9046 7616 9052
rect 7470 9007 7526 9016
rect 7484 8906 7512 9007
rect 7562 8936 7618 8945
rect 7472 8900 7524 8906
rect 7562 8871 7618 8880
rect 7472 8842 7524 8848
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7392 7834 7420 8230
rect 7300 7806 7420 7834
rect 7300 7546 7328 7806
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 7300 7002 7328 7375
rect 7392 7274 7420 7686
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7288 6996 7340 7002
rect 7340 6956 7420 6984
rect 7288 6938 7340 6944
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 6932 5868 7144 5896
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3936 6696 3942
rect 6828 3936 6880 3942
rect 6644 3878 6696 3884
rect 6748 3884 6828 3890
rect 6748 3878 6880 3884
rect 6472 3454 6592 3482
rect 6366 3431 6422 3440
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 2990 6500 3295
rect 6564 3126 6592 3454
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6380 1057 6408 2926
rect 6472 2854 6500 2926
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6656 2417 6684 3878
rect 6748 3862 6868 3878
rect 6748 3466 6776 3862
rect 6932 3720 6960 5714
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7024 4049 7052 5034
rect 7116 4758 7144 5868
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7116 4282 7144 4694
rect 7208 4554 7236 6122
rect 7288 6112 7340 6118
rect 7286 6080 7288 6089
rect 7340 6080 7342 6089
rect 7286 6015 7342 6024
rect 7300 5778 7328 6015
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7392 4826 7420 6956
rect 7484 6118 7512 8842
rect 7576 7954 7604 8871
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7196 4072 7248 4078
rect 7010 4040 7066 4049
rect 7196 4014 7248 4020
rect 7010 3975 7066 3984
rect 7024 3738 7052 3975
rect 7208 3942 7236 4014
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 6840 3692 6960 3720
rect 7012 3732 7064 3738
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6734 3088 6790 3097
rect 6734 3023 6790 3032
rect 6642 2408 6698 2417
rect 6642 2343 6698 2352
rect 6748 2038 6776 3023
rect 6840 2938 6868 3692
rect 7012 3674 7064 3680
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7102 3496 7158 3505
rect 7024 3233 7052 3470
rect 7102 3431 7158 3440
rect 7010 3224 7066 3233
rect 7010 3159 7066 3168
rect 7116 3058 7144 3431
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7208 2990 7236 3878
rect 7300 3194 7328 4694
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7196 2984 7248 2990
rect 7010 2952 7066 2961
rect 6840 2910 6960 2938
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6366 1048 6422 1057
rect 6366 983 6422 992
rect 6458 82 6514 480
rect 6840 241 6868 2790
rect 6932 921 6960 2910
rect 7196 2926 7248 2932
rect 7010 2887 7066 2896
rect 7024 2854 7052 2887
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7010 2680 7066 2689
rect 7010 2615 7066 2624
rect 7024 2582 7052 2615
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6918 912 6974 921
rect 6918 847 6974 856
rect 6826 232 6882 241
rect 6826 167 6882 176
rect 6196 54 6514 82
rect 7392 82 7420 4150
rect 7484 3777 7512 5238
rect 7576 4758 7604 7414
rect 7668 7410 7696 10775
rect 7748 10746 7800 10752
rect 7760 10470 7788 10746
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 9024 7788 10406
rect 7852 10266 7880 11104
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7838 10160 7894 10169
rect 7838 10095 7894 10104
rect 7852 9489 7880 10095
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7760 8996 7880 9024
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 8022 7788 8842
rect 7852 8537 7880 8996
rect 7838 8528 7894 8537
rect 7838 8463 7894 8472
rect 7838 8256 7894 8265
rect 7838 8191 7894 8200
rect 7852 8022 7880 8191
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7760 7546 7788 7958
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 5778 7696 6870
rect 7944 6866 7972 11018
rect 8036 10062 8064 11240
rect 8128 11121 8156 11308
rect 8114 11112 8170 11121
rect 8114 11047 8170 11056
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10674 8156 10950
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8114 10568 8170 10577
rect 8114 10503 8170 10512
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9518 8064 9862
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 9178 8064 9318
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8128 9042 8156 10503
rect 8220 9761 8248 12650
rect 8312 9926 8340 16934
rect 8404 16182 8432 18566
rect 8496 17202 8524 20810
rect 8588 20233 8616 21422
rect 8574 20224 8630 20233
rect 8574 20159 8630 20168
rect 8574 19952 8630 19961
rect 8574 19887 8630 19896
rect 8588 19446 8616 19887
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8574 19136 8630 19145
rect 8574 19071 8630 19080
rect 8588 18970 8616 19071
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8496 16522 8524 17002
rect 8588 16726 8616 18702
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 15745 8432 15846
rect 8390 15736 8446 15745
rect 8390 15671 8446 15680
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8404 15094 8432 15574
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8404 14550 8432 15030
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8404 13530 8432 14350
rect 8496 13814 8524 15574
rect 8588 15094 8616 16662
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8588 14006 8616 14418
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8496 13786 8616 13814
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12617 8432 13126
rect 8390 12608 8446 12617
rect 8390 12543 8446 12552
rect 8390 12472 8446 12481
rect 8390 12407 8446 12416
rect 8404 12238 8432 12407
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8390 12064 8446 12073
rect 8390 11999 8446 12008
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8206 9752 8262 9761
rect 8206 9687 8262 9696
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8036 8634 8064 8978
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8036 8401 8064 8570
rect 8022 8392 8078 8401
rect 8022 8327 8078 8336
rect 8128 8276 8156 8978
rect 8220 8362 8248 9522
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8312 8809 8340 9386
rect 8298 8800 8354 8809
rect 8298 8735 8354 8744
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8036 8248 8156 8276
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6390 7880 6598
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7668 4672 7696 5714
rect 7576 4644 7696 4672
rect 7576 4321 7604 4644
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7562 4312 7618 4321
rect 7562 4247 7618 4256
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7470 3768 7526 3777
rect 7470 3703 7526 3712
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 2990 7512 3470
rect 7576 3194 7604 4014
rect 7668 3466 7696 4558
rect 7760 4554 7788 6326
rect 7852 6254 7880 6326
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7944 5778 7972 6802
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7838 5672 7894 5681
rect 7838 5607 7894 5616
rect 7852 5234 7880 5607
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7838 4992 7894 5001
rect 7838 4927 7894 4936
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7746 4312 7802 4321
rect 7746 4247 7802 4256
rect 7760 3942 7788 4247
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7760 3346 7788 3606
rect 7668 3318 7788 3346
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7576 2446 7604 2751
rect 7668 2582 7696 3318
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7470 82 7526 480
rect 7760 377 7788 2858
rect 7852 2514 7880 4927
rect 8036 4457 8064 8248
rect 8312 8242 8340 8735
rect 8404 8362 8432 11999
rect 8496 11558 8524 13670
rect 8588 13258 8616 13786
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8574 12744 8630 12753
rect 8574 12679 8630 12688
rect 8588 12646 8616 12679
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8482 11384 8538 11393
rect 8588 11354 8616 12378
rect 8482 11319 8538 11328
rect 8576 11348 8628 11354
rect 8496 10606 8524 11319
rect 8576 11290 8628 11296
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 10044 8524 10406
rect 8574 10296 8630 10305
rect 8574 10231 8630 10240
rect 8588 10198 8616 10231
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8496 10016 8616 10044
rect 8484 9920 8536 9926
rect 8588 9897 8616 10016
rect 8484 9862 8536 9868
rect 8574 9888 8630 9897
rect 8496 8537 8524 9862
rect 8574 9823 8630 9832
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8588 8820 8616 9454
rect 8680 9178 8708 22392
rect 9220 22374 9272 22380
rect 9232 21593 9260 22374
rect 8850 21584 8906 21593
rect 8850 21519 8906 21528
rect 9218 21584 9274 21593
rect 9600 21554 9628 23122
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9772 22296 9824 22302
rect 9678 22264 9734 22273
rect 9862 22264 9918 22273
rect 9824 22244 9862 22250
rect 9772 22238 9862 22244
rect 9784 22222 9862 22238
rect 9678 22199 9734 22208
rect 9862 22199 9918 22208
rect 9218 21519 9274 21528
rect 9588 21548 9640 21554
rect 8758 21312 8814 21321
rect 8758 21247 8814 21256
rect 8772 21146 8800 21247
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8864 21026 8892 21519
rect 9588 21490 9640 21496
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 8772 20998 8892 21026
rect 9220 21004 9272 21010
rect 8772 19825 8800 20998
rect 9220 20946 9272 20952
rect 8944 20800 8996 20806
rect 9232 20777 9260 20946
rect 8944 20742 8996 20748
rect 9034 20768 9090 20777
rect 8956 20346 8984 20742
rect 9034 20703 9090 20712
rect 9218 20768 9274 20777
rect 9218 20703 9274 20712
rect 9048 20398 9076 20703
rect 8864 20318 8984 20346
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 8758 19816 8814 19825
rect 8758 19751 8814 19760
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8772 18057 8800 19654
rect 8864 19281 8892 20318
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8956 19689 8984 19858
rect 8942 19680 8998 19689
rect 8942 19615 8998 19624
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 19281 9076 19314
rect 8850 19272 8906 19281
rect 8850 19207 8906 19216
rect 9034 19272 9090 19281
rect 9034 19207 9090 19216
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8852 18080 8904 18086
rect 8758 18048 8814 18057
rect 8956 18068 8984 18566
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8904 18040 8984 18068
rect 8852 18022 8904 18028
rect 9048 18000 9076 18158
rect 8758 17983 8814 17992
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8758 17912 8814 17921
rect 8956 17904 9252 17924
rect 8814 17882 8892 17898
rect 8814 17876 8904 17882
rect 8814 17870 8852 17876
rect 8758 17847 8814 17856
rect 8852 17818 8904 17824
rect 9048 17649 9076 17904
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9034 17640 9090 17649
rect 9034 17575 9090 17584
rect 8852 17536 8904 17542
rect 8758 17504 8814 17513
rect 8852 17478 8904 17484
rect 8758 17439 8814 17448
rect 8772 16454 8800 17439
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8772 15638 8800 16118
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8864 15473 8892 17478
rect 9232 17338 9260 17682
rect 9324 17649 9352 21354
rect 9310 17640 9366 17649
rect 9310 17575 9366 17584
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 8956 16425 8984 16662
rect 9324 16590 9352 17478
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9036 16448 9088 16454
rect 8942 16416 8998 16425
rect 9036 16390 9088 16396
rect 9126 16416 9182 16425
rect 8942 16351 8998 16360
rect 9048 16266 9076 16390
rect 9126 16351 9182 16360
rect 8956 16238 9076 16266
rect 8956 15824 8984 16238
rect 9140 15978 9168 16351
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9232 15824 9260 16458
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 8956 15804 9260 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 9252 15748 9260 15804
rect 8956 15728 9260 15748
rect 8850 15464 8906 15473
rect 8850 15399 8906 15408
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8772 14618 8800 14826
rect 8956 14736 8984 15728
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9140 14890 9168 15030
rect 9232 14940 9260 15728
rect 9324 15065 9352 16390
rect 9310 15056 9366 15065
rect 9310 14991 9366 15000
rect 9232 14912 9352 14940
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8772 14074 8800 14554
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8864 13920 8892 14554
rect 8956 14006 8984 14640
rect 9324 14600 9352 14912
rect 9048 14572 9352 14600
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8772 13892 8892 13920
rect 8772 13462 8800 13892
rect 8956 13814 8984 13942
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8950 13786 8984 13814
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8772 12986 8800 13398
rect 8864 13190 8892 13738
rect 8950 13648 8978 13786
rect 9048 13716 9076 14572
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9140 13870 9168 14418
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9048 13688 9168 13716
rect 9140 13648 9168 13688
rect 9232 13648 9260 14214
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9324 13977 9352 14010
rect 9310 13968 9366 13977
rect 9310 13903 9366 13912
rect 9324 13784 9352 13903
rect 9416 13802 9444 21354
rect 9692 21321 9720 22199
rect 9678 21312 9734 21321
rect 9678 21247 9734 21256
rect 9632 21176 9688 21185
rect 9508 21134 9632 21162
rect 9508 20913 9536 21134
rect 9632 21111 9688 21120
rect 9588 21072 9640 21078
rect 9588 21014 9640 21020
rect 9494 20904 9550 20913
rect 9494 20839 9550 20848
rect 9600 20534 9628 21014
rect 9968 21010 9996 22714
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10060 21486 10088 21626
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9692 20534 9720 20810
rect 9968 20602 9996 20946
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9508 19009 9536 19722
rect 9600 19514 9628 19858
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9494 19000 9550 19009
rect 9600 18952 9628 19450
rect 9692 18952 9720 20470
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 9550 18944 9720 18952
rect 9494 18935 9720 18944
rect 9508 18924 9720 18935
rect 9508 18426 9536 18924
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9494 18320 9550 18329
rect 9494 18255 9550 18264
rect 9508 17105 9536 18255
rect 9600 18170 9628 18924
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18426 9720 18770
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9600 18142 9720 18170
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17241 9628 18022
rect 9692 17746 9720 18142
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17338 9720 17682
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9586 17232 9642 17241
rect 9586 17167 9642 17176
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 9692 16572 9720 17138
rect 9784 16697 9812 20266
rect 10060 20262 10088 21422
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 18748 9904 19858
rect 10060 19786 10088 20198
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9968 19292 9996 19654
rect 10048 19304 10100 19310
rect 9968 19264 10048 19292
rect 10048 19246 10100 19252
rect 9956 18760 10008 18766
rect 9876 18720 9956 18748
rect 9956 18702 10008 18708
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9968 18222 9996 18362
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 10060 18154 10088 19246
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9864 16720 9916 16726
rect 9770 16688 9826 16697
rect 9864 16662 9916 16668
rect 9770 16623 9826 16632
rect 9772 16584 9824 16590
rect 9692 16544 9772 16572
rect 9772 16526 9824 16532
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9404 13796 9456 13802
rect 9324 13756 9404 13784
rect 9404 13738 9456 13744
rect 8950 13628 9260 13648
rect 8950 13572 8956 13628
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 9252 13572 9260 13628
rect 8950 13552 9260 13572
rect 8950 13512 8978 13552
rect 8950 13484 8984 13512
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8758 12064 8814 12073
rect 8758 11999 8814 12008
rect 8772 10810 8800 11999
rect 8864 11762 8892 13126
rect 8956 12889 8984 13484
rect 8942 12880 8998 12889
rect 8942 12815 8998 12824
rect 9140 12753 9168 13552
rect 9232 12986 9260 13552
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12918 9352 13126
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9126 12744 9182 12753
rect 9324 12714 9352 12854
rect 9416 12850 9444 13738
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9402 12744 9458 12753
rect 9126 12679 9182 12688
rect 9312 12708 9364 12714
rect 9402 12679 9458 12688
rect 9312 12650 9364 12656
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 9126 12336 9182 12345
rect 8944 12300 8996 12306
rect 9126 12271 9182 12280
rect 8944 12242 8996 12248
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8956 11642 8984 12242
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8864 11614 8984 11642
rect 8864 11336 8892 11614
rect 9048 11472 9076 12174
rect 9140 11472 9168 12271
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 8864 11308 8984 11336
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8758 10432 8814 10441
rect 8758 10367 8814 10376
rect 8772 10130 8800 10367
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8864 9364 8892 11154
rect 8956 10384 8984 11308
rect 9048 11286 9076 11376
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10742 9076 10950
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9140 10674 9168 11376
rect 9324 11354 9352 12038
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9232 10384 9260 11222
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 8956 10364 9260 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 9252 10308 9260 10364
rect 8956 10288 9260 10308
rect 8956 9364 8984 10288
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9722 9076 9862
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8758 9344 8814 9353
rect 8864 9336 8984 9364
rect 8864 9330 8892 9336
rect 8814 9302 8892 9330
rect 8758 9279 8814 9288
rect 8758 9208 8814 9217
rect 8668 9172 8720 9178
rect 8758 9143 8814 9152
rect 8668 9114 8720 9120
rect 8772 9042 8800 9143
rect 8864 9058 8892 9302
rect 9232 9296 9260 10288
rect 9324 10282 9352 10950
rect 9416 10810 9444 12679
rect 9508 11898 9536 16050
rect 9600 14482 9628 16458
rect 9876 16114 9904 16662
rect 9968 16182 9996 17478
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 14793 9720 15302
rect 9784 15094 9812 15438
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9678 14784 9734 14793
rect 9678 14719 9734 14728
rect 9678 14512 9734 14521
rect 9588 14476 9640 14482
rect 9678 14447 9734 14456
rect 9588 14418 9640 14424
rect 9600 14346 9628 14418
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9692 14260 9720 14447
rect 9784 14385 9812 15030
rect 9876 14890 9904 15574
rect 9968 14906 9996 15642
rect 10060 15434 10088 17546
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 9864 14884 9916 14890
rect 9968 14878 10088 14906
rect 9864 14826 9916 14832
rect 9876 14618 9904 14826
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9968 14414 9996 14758
rect 9956 14408 10008 14414
rect 9770 14376 9826 14385
rect 9956 14350 10008 14356
rect 9770 14311 9826 14320
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9692 14232 9812 14260
rect 9678 14104 9734 14113
rect 9678 14039 9734 14048
rect 9692 14006 9720 14039
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9600 13326 9628 13359
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9600 11608 9628 12922
rect 9508 11580 9628 11608
rect 9508 11014 9536 11580
rect 9586 11520 9642 11529
rect 9586 11455 9642 11464
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9416 10606 9444 10746
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9324 10254 9444 10282
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 8956 9276 9260 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 9252 9220 9260 9276
rect 8956 9200 9260 9220
rect 8760 9036 8812 9042
rect 8864 9030 8984 9058
rect 8760 8978 8812 8984
rect 8850 8936 8906 8945
rect 8680 8894 8850 8922
rect 8680 8820 8708 8894
rect 8850 8871 8906 8880
rect 8588 8809 8800 8820
rect 8574 8800 8800 8809
rect 8630 8792 8800 8800
rect 8574 8735 8630 8744
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8496 8362 8524 8463
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8482 8256 8538 8265
rect 8312 8214 8432 8242
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8128 7546 8156 7890
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 7426 8248 7686
rect 8128 7398 8248 7426
rect 8128 6633 8156 7398
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8220 7002 8248 7210
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8220 6866 8248 6938
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8114 6624 8170 6633
rect 8114 6559 8170 6568
rect 8220 6254 8248 6802
rect 8312 6730 8340 8026
rect 8404 7954 8432 8214
rect 8482 8191 8538 8200
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8390 7576 8446 7585
rect 8496 7546 8524 8191
rect 8588 7721 8616 8735
rect 8574 7712 8630 7721
rect 8574 7647 8630 7656
rect 8390 7511 8446 7520
rect 8484 7540 8536 7546
rect 8404 6934 8432 7511
rect 8484 7482 8536 7488
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8484 6792 8536 6798
rect 8390 6760 8446 6769
rect 8300 6724 8352 6730
rect 8484 6734 8536 6740
rect 8390 6695 8446 6704
rect 8300 6666 8352 6672
rect 8208 6248 8260 6254
rect 8128 6208 8208 6236
rect 8128 5030 8156 6208
rect 8208 6190 8260 6196
rect 8298 5944 8354 5953
rect 8208 5908 8260 5914
rect 8404 5914 8432 6695
rect 8298 5879 8354 5888
rect 8392 5908 8444 5914
rect 8208 5850 8260 5856
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8114 4856 8170 4865
rect 8114 4791 8170 4800
rect 8128 4758 8156 4791
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8022 4448 8078 4457
rect 8022 4383 8078 4392
rect 8022 4312 8078 4321
rect 8128 4282 8156 4694
rect 8022 4247 8078 4256
rect 8116 4276 8168 4282
rect 7930 4176 7986 4185
rect 7930 4111 7986 4120
rect 7944 3670 7972 4111
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 8036 2650 8064 4247
rect 8116 4218 8168 4224
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8128 3913 8156 3946
rect 8114 3904 8170 3913
rect 8114 3839 8170 3848
rect 8220 3777 8248 5850
rect 8312 5098 8340 5879
rect 8392 5850 8444 5856
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8404 5030 8432 5510
rect 8496 5148 8524 6734
rect 8588 5953 8616 7210
rect 8680 7206 8708 8792
rect 8772 8401 8800 8792
rect 8852 8492 8904 8498
rect 8956 8480 8984 9030
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8904 8452 8984 8480
rect 8852 8434 8904 8440
rect 8758 8392 8814 8401
rect 8758 8327 8814 8336
rect 8864 8242 8892 8434
rect 9140 8430 9168 8774
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9232 8276 9260 9200
rect 8772 8214 8892 8242
rect 8956 8248 9260 8276
rect 8772 7750 8800 8214
rect 8956 8208 8984 8248
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8574 5944 8630 5953
rect 8574 5879 8630 5888
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 5302 8616 5714
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8496 5120 8616 5148
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 3942 8340 4694
rect 8404 4593 8432 4966
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8390 4584 8446 4593
rect 8390 4519 8446 4528
rect 8496 4154 8524 4762
rect 8588 4622 8616 5120
rect 8680 5012 8708 6938
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8772 5166 8800 6870
rect 8864 5896 8892 7890
rect 8956 7120 8984 8112
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7585 9168 7686
rect 9126 7576 9182 7585
rect 9126 7511 9182 7520
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 8956 6168 8984 7024
rect 9324 6458 9352 10134
rect 9416 8090 9444 10254
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9508 7954 9536 10678
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9402 7576 9458 7585
rect 9402 7511 9458 7520
rect 9416 7342 9444 7511
rect 9404 7336 9456 7342
rect 9456 7296 9536 7324
rect 9404 7278 9456 7284
rect 9402 7168 9458 7177
rect 9402 7103 9458 7112
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9324 6186 9352 6394
rect 9416 6322 9444 7103
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9036 6180 9088 6186
rect 8956 6140 9036 6168
rect 9036 6122 9088 6128
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 9402 5944 9458 5953
rect 8864 5868 8984 5896
rect 9402 5879 9458 5888
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8680 4984 8800 5012
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8404 4126 8524 4154
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8206 3768 8262 3777
rect 8312 3738 8340 3878
rect 8206 3703 8262 3712
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8114 3632 8170 3641
rect 8114 3567 8170 3576
rect 8298 3632 8354 3641
rect 8298 3567 8354 3576
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8128 2582 8156 3567
rect 8312 3369 8340 3567
rect 8298 3360 8354 3369
rect 8298 3295 8354 3304
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8220 2922 8248 3130
rect 8404 3058 8432 4126
rect 8588 4060 8616 4422
rect 8496 4032 8616 4060
rect 8680 4049 8708 4694
rect 8666 4040 8722 4049
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8128 513 8156 2518
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8114 504 8170 513
rect 8114 439 8170 448
rect 7746 368 7802 377
rect 7746 303 7802 312
rect 7392 54 7526 82
rect 8404 82 8432 2314
rect 8496 1465 8524 4032
rect 8666 3975 8668 3984
rect 8720 3975 8722 3984
rect 8668 3946 8720 3952
rect 8680 3915 8708 3946
rect 8772 3754 8800 4984
rect 8864 4457 8892 5646
rect 8956 5137 8984 5868
rect 9034 5400 9090 5409
rect 9128 5364 9180 5370
rect 9090 5344 9128 5352
rect 9034 5335 9128 5344
rect 9048 5324 9128 5335
rect 9128 5306 9180 5312
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 8942 5128 8998 5137
rect 8942 5063 8998 5072
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 8850 4448 8906 4457
rect 8850 4383 8906 4392
rect 9324 4282 9352 5238
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 9218 4176 9274 4185
rect 8680 3726 8800 3754
rect 8574 3360 8630 3369
rect 8574 3295 8630 3304
rect 8588 3058 8616 3295
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8680 2825 8708 3726
rect 8864 3584 8892 4150
rect 9218 4111 9274 4120
rect 9232 4010 9260 4111
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8864 3556 8984 3584
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8666 2816 8722 2825
rect 8666 2751 8722 2760
rect 8482 1456 8538 1465
rect 8482 1391 8538 1400
rect 8772 785 8800 3334
rect 8850 2952 8906 2961
rect 8956 2922 8984 3556
rect 9048 2961 9076 3606
rect 9128 3596 9180 3602
rect 9180 3556 9352 3584
rect 9128 3538 9180 3544
rect 9218 3088 9274 3097
rect 9218 3023 9274 3032
rect 9034 2952 9090 2961
rect 8850 2887 8906 2896
rect 8944 2916 8996 2922
rect 8864 2582 8892 2887
rect 9232 2922 9260 3023
rect 9034 2887 9090 2896
rect 9220 2916 9272 2922
rect 8944 2858 8996 2864
rect 9220 2858 9272 2864
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 8956 2038 8984 2518
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 9324 1902 9352 3556
rect 9416 3058 9444 5879
rect 9508 5846 9536 7296
rect 9600 6798 9628 11455
rect 9692 10130 9720 13670
rect 9784 13025 9812 14232
rect 9770 13016 9826 13025
rect 9770 12951 9826 12960
rect 9876 12850 9904 14282
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9876 12374 9904 12786
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9862 12200 9918 12209
rect 9862 12135 9918 12144
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 10674 9812 11698
rect 9876 11354 9904 12135
rect 9968 12102 9996 13262
rect 10060 12345 10088 14878
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9954 11928 10010 11937
rect 9954 11863 10010 11872
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9772 10668 9824 10674
rect 9824 10628 9904 10656
rect 9772 10610 9824 10616
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9692 9722 9720 10066
rect 9784 9994 9812 10474
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9876 9926 9904 10628
rect 9968 10577 9996 11863
rect 10060 11014 10088 12174
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10606 10088 10950
rect 10048 10600 10100 10606
rect 9954 10568 10010 10577
rect 10048 10542 10100 10548
rect 9954 10503 10010 10512
rect 10048 10464 10100 10470
rect 10046 10432 10048 10441
rect 10100 10432 10102 10441
rect 10046 10367 10102 10376
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9508 5234 9536 5782
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9508 4690 9536 5170
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9494 4584 9550 4593
rect 9600 4554 9628 6734
rect 9692 6497 9720 9454
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9784 8974 9812 9007
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8498 9812 8910
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9876 8566 9904 8774
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9864 8356 9916 8362
rect 9784 7546 9812 8327
rect 9864 8298 9916 8304
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9678 6488 9734 6497
rect 9678 6423 9734 6432
rect 9772 6112 9824 6118
rect 9678 6080 9734 6089
rect 9772 6054 9824 6060
rect 9678 6015 9734 6024
rect 9692 5642 9720 6015
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5234 9720 5578
rect 9784 5234 9812 6054
rect 9876 5302 9904 8298
rect 9968 5710 9996 10202
rect 10060 9926 10088 10367
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 7478 10088 9318
rect 10152 9178 10180 19178
rect 10244 18358 10272 21558
rect 10428 21486 10456 23582
rect 11624 23582 12034 23610
rect 10600 22296 10652 22302
rect 10600 22238 10652 22244
rect 10506 21856 10562 21865
rect 10506 21791 10562 21800
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10336 18222 10364 18838
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10152 8498 10180 9114
rect 10244 9042 10272 18022
rect 10336 17921 10364 18158
rect 10322 17912 10378 17921
rect 10322 17847 10378 17856
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10336 16794 10364 17750
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10336 15026 10364 15370
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10336 14550 10364 14826
rect 10428 14618 10456 20266
rect 10520 16266 10548 21791
rect 10612 18465 10640 22238
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10874 21584 10930 21593
rect 10874 21519 10930 21528
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10598 18456 10654 18465
rect 10598 18391 10654 18400
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10612 17746 10640 18090
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10612 16436 10640 17682
rect 10704 17377 10732 20742
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10796 19718 10824 20334
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10690 17368 10746 17377
rect 10690 17303 10746 17312
rect 10692 16448 10744 16454
rect 10612 16408 10692 16436
rect 10692 16390 10744 16396
rect 10520 16238 10640 16266
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10520 15162 10548 15982
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10506 15056 10562 15065
rect 10506 14991 10562 15000
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10428 13938 10456 14554
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10428 13462 10456 13670
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10428 12646 10456 13398
rect 10520 12918 10548 14991
rect 10612 14074 10640 16238
rect 10704 16182 10732 16390
rect 10796 16250 10824 19654
rect 10888 17814 10916 21519
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 17202 10916 17546
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 14278 10732 15846
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10704 13705 10732 13738
rect 10690 13696 10746 13705
rect 10690 13631 10746 13640
rect 10796 13530 10824 14350
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12986 10640 13126
rect 10600 12980 10652 12986
rect 10888 12968 10916 16730
rect 10980 15638 11008 22102
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 20534 11100 21286
rect 11256 20788 11284 21354
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11348 20942 11376 21286
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11440 20806 11468 20946
rect 11428 20800 11480 20806
rect 11256 20760 11376 20788
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11242 20224 11298 20233
rect 11164 19990 11192 20198
rect 11242 20159 11298 20168
rect 11152 19984 11204 19990
rect 11152 19926 11204 19932
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11072 19174 11100 19858
rect 11152 19508 11204 19514
rect 11256 19496 11284 20159
rect 11204 19468 11284 19496
rect 11152 19450 11204 19456
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11060 19168 11112 19174
rect 11058 19136 11060 19145
rect 11112 19136 11114 19145
rect 11058 19071 11114 19080
rect 11072 18834 11100 19071
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11072 18426 11100 18770
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11164 18601 11192 18634
rect 11150 18592 11206 18601
rect 11150 18527 11206 18536
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11072 18086 11100 18362
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 15910 11100 16934
rect 11164 16833 11192 18362
rect 11256 17202 11284 19314
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11150 16824 11206 16833
rect 11150 16759 11206 16768
rect 11164 16658 11192 16759
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 16046 11192 16458
rect 11256 16250 11284 17138
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 11152 15632 11204 15638
rect 11204 15592 11284 15620
rect 11152 15574 11204 15580
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11072 14929 11100 15302
rect 11058 14920 11114 14929
rect 10968 14884 11020 14890
rect 11058 14855 11114 14864
rect 10968 14826 11020 14832
rect 10600 12922 10652 12928
rect 10704 12940 10916 12968
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10612 12646 10640 12922
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10428 11694 10456 12582
rect 10506 12200 10562 12209
rect 10704 12186 10732 12940
rect 10782 12880 10838 12889
rect 10782 12815 10838 12824
rect 10506 12135 10562 12144
rect 10612 12158 10732 12186
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10336 9178 10364 11562
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10674 10456 11154
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7546 10180 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10244 7324 10272 8774
rect 10060 7296 10272 7324
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9954 5536 10010 5545
rect 9954 5471 10010 5480
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9968 5080 9996 5471
rect 10060 5409 10088 7296
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10152 5914 10180 6666
rect 10244 6186 10272 6734
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10244 5914 10272 6122
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10152 5817 10180 5850
rect 10138 5808 10194 5817
rect 10138 5743 10194 5752
rect 10046 5400 10102 5409
rect 10046 5335 10102 5344
rect 10322 5400 10378 5409
rect 10322 5335 10378 5344
rect 10336 5234 10364 5335
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 9968 5052 10088 5080
rect 9862 4992 9918 5001
rect 9918 4950 9996 4978
rect 9862 4927 9918 4936
rect 9678 4856 9734 4865
rect 9678 4791 9734 4800
rect 9692 4604 9720 4791
rect 9772 4616 9824 4622
rect 9692 4576 9772 4604
rect 9772 4558 9824 4564
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9494 4519 9550 4528
rect 9588 4548 9640 4554
rect 9508 3602 9536 4519
rect 9588 4490 9640 4496
rect 9600 4214 9628 4490
rect 9770 4312 9826 4321
rect 9770 4247 9826 4256
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9586 4040 9642 4049
rect 9586 3975 9642 3984
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9600 3466 9628 3975
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9402 2952 9458 2961
rect 9402 2887 9458 2896
rect 9416 2009 9444 2887
rect 9508 2582 9536 3130
rect 9692 2854 9720 3538
rect 9784 3126 9812 4247
rect 9876 4185 9904 4558
rect 9862 4176 9918 4185
rect 9862 4111 9918 4120
rect 9968 3738 9996 4950
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9954 3632 10010 3641
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9402 2000 9458 2009
rect 9402 1935 9458 1944
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 8758 776 8814 785
rect 8758 711 8814 720
rect 8482 82 8538 480
rect 8404 54 8538 82
rect 3422 0 3478 54
rect 4434 0 4490 54
rect 5446 0 5502 54
rect 6458 0 6514 54
rect 7470 0 7526 54
rect 8482 0 8538 54
rect 9402 82 9458 480
rect 9692 82 9720 2790
rect 9876 2582 9904 3606
rect 9954 3567 10010 3576
rect 9968 3126 9996 3567
rect 10060 3126 10088 5052
rect 10138 4992 10194 5001
rect 10138 4927 10194 4936
rect 10152 4185 10180 4927
rect 10230 4584 10286 4593
rect 10230 4519 10286 4528
rect 10138 4176 10194 4185
rect 10244 4146 10272 4519
rect 10322 4176 10378 4185
rect 10138 4111 10194 4120
rect 10232 4140 10284 4146
rect 10322 4111 10378 4120
rect 10232 4082 10284 4088
rect 10336 4010 10364 4111
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10138 3904 10194 3913
rect 10138 3839 10194 3848
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10046 2680 10102 2689
rect 10046 2615 10102 2624
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 10060 2310 10088 2615
rect 10152 2582 10180 3839
rect 10322 3768 10378 3777
rect 10322 3703 10378 3712
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 2961 10272 3470
rect 10230 2952 10286 2961
rect 10336 2922 10364 3703
rect 10428 3058 10456 9998
rect 10520 9722 10548 12135
rect 10612 10266 10640 12158
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11558 10732 12038
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10690 10704 10746 10713
rect 10690 10639 10746 10648
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10704 10130 10732 10639
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 8498 10548 9318
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10520 8090 10548 8298
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7313 10548 7686
rect 10506 7304 10562 7313
rect 10506 7239 10562 7248
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 6866 10548 7142
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10612 5778 10640 9386
rect 10704 8809 10732 9862
rect 10690 8800 10746 8809
rect 10690 8735 10746 8744
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10704 6798 10732 8570
rect 10796 8129 10824 12815
rect 10876 12708 10928 12714
rect 10980 12696 11008 14826
rect 11164 14822 11192 15302
rect 11256 15162 11284 15592
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11256 14634 11284 14894
rect 11164 14606 11284 14634
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10928 12668 11008 12696
rect 10876 12650 10928 12656
rect 10888 12238 10916 12650
rect 10966 12608 11022 12617
rect 10966 12543 11022 12552
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10874 11928 10930 11937
rect 10874 11863 10930 11872
rect 10888 11694 10916 11863
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11354 10916 11630
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10888 10742 10916 11018
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10130 10916 10406
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9178 10916 10066
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10782 8120 10838 8129
rect 10782 8055 10838 8064
rect 10782 7712 10838 7721
rect 10782 7647 10838 7656
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6118 10732 6598
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10704 5846 10732 6054
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10230 2887 10286 2896
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10152 1834 10180 2518
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 9402 54 9720 82
rect 10414 82 10470 480
rect 10520 82 10548 5238
rect 10612 4865 10640 5510
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10598 4856 10654 4865
rect 10598 4791 10654 4800
rect 10598 4312 10654 4321
rect 10598 4247 10654 4256
rect 10612 2650 10640 4247
rect 10704 3738 10732 4966
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10704 3194 10732 3538
rect 10796 3534 10824 7647
rect 10888 7410 10916 8570
rect 10980 7886 11008 12543
rect 11072 12306 11100 13466
rect 11164 12345 11192 14606
rect 11348 14074 11376 20760
rect 11428 20742 11480 20748
rect 11440 19718 11468 20742
rect 11518 20496 11574 20505
rect 11518 20431 11574 20440
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11440 18290 11468 18770
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11440 17882 11468 18226
rect 11532 17882 11560 20431
rect 11624 19514 11652 23582
rect 11978 23520 12034 23582
rect 13740 23582 13874 23610
rect 13542 23080 13598 23089
rect 13542 23015 13598 23024
rect 13556 22001 13584 23015
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13542 21992 13598 22001
rect 13542 21927 13598 21936
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12806 21720 12862 21729
rect 12956 21712 13252 21732
rect 12806 21655 12862 21664
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 11888 21072 11940 21078
rect 11888 21014 11940 21020
rect 11900 20913 11928 21014
rect 11980 20936 12032 20942
rect 11886 20904 11942 20913
rect 11980 20878 12032 20884
rect 11886 20839 11942 20848
rect 11900 20398 11928 20839
rect 11992 20777 12020 20878
rect 11978 20768 12034 20777
rect 11978 20703 12034 20712
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11624 17270 11652 17682
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11624 16658 11652 17002
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11440 16114 11468 16594
rect 11624 16182 11652 16594
rect 11612 16176 11664 16182
rect 11612 16118 11664 16124
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11426 15736 11482 15745
rect 11426 15671 11482 15680
rect 11440 15502 11468 15671
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11440 15201 11468 15438
rect 11426 15192 11482 15201
rect 11426 15127 11482 15136
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11334 13968 11390 13977
rect 11334 13903 11390 13912
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11150 12336 11206 12345
rect 11060 12300 11112 12306
rect 11150 12271 11206 12280
rect 11060 12242 11112 12248
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11072 11286 11100 12038
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11072 10810 11100 11222
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11164 10198 11192 12038
rect 11256 11665 11284 13126
rect 11348 12170 11376 13903
rect 11440 13161 11468 14758
rect 11426 13152 11482 13161
rect 11426 13087 11482 13096
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 11242 11656 11298 11665
rect 11242 11591 11298 11600
rect 11440 11506 11468 12582
rect 11256 11478 11468 11506
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9489 11100 9522
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11072 8022 11100 8502
rect 11164 8090 11192 10134
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 7313 11008 7346
rect 10966 7304 11022 7313
rect 11072 7274 11100 7754
rect 10966 7239 11022 7248
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11164 6934 11192 7822
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 3913 10916 6598
rect 10980 6186 11008 6666
rect 11150 6488 11206 6497
rect 11150 6423 11206 6432
rect 11164 6186 11192 6423
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 4826 11100 6054
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11164 4758 11192 5510
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10966 4040 11022 4049
rect 10966 3975 11022 3984
rect 10874 3904 10930 3913
rect 10874 3839 10930 3848
rect 10874 3632 10930 3641
rect 10874 3567 10930 3576
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10690 3088 10746 3097
rect 10888 3058 10916 3567
rect 10980 3466 11008 3975
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3466 11100 3878
rect 11164 3602 11192 4082
rect 11256 4078 11284 11478
rect 11426 11112 11482 11121
rect 11336 11076 11388 11082
rect 11426 11047 11482 11056
rect 11336 11018 11388 11024
rect 11348 10713 11376 11018
rect 11334 10704 11390 10713
rect 11334 10639 11390 10648
rect 11334 10568 11390 10577
rect 11334 10503 11390 10512
rect 11348 8401 11376 10503
rect 11440 8498 11468 11047
rect 11532 10266 11560 15914
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11532 8634 11560 10202
rect 11624 8945 11652 14010
rect 11716 12918 11744 20266
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17241 11836 18022
rect 11794 17232 11850 17241
rect 11794 17167 11850 17176
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11702 12608 11758 12617
rect 11702 12543 11758 12552
rect 11716 12442 11744 12543
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11716 10810 11744 12242
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10169 11744 10406
rect 11702 10160 11758 10169
rect 11702 10095 11758 10104
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11610 8936 11666 8945
rect 11610 8871 11666 8880
rect 11610 8800 11666 8809
rect 11610 8735 11666 8744
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11520 8424 11572 8430
rect 11334 8392 11390 8401
rect 11520 8366 11572 8372
rect 11334 8327 11390 8336
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11348 4457 11376 7754
rect 11440 7206 11468 8230
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11532 6662 11560 8366
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11334 4448 11390 4457
rect 11334 4383 11390 4392
rect 11624 4264 11652 8735
rect 11716 8634 11744 9046
rect 11808 8650 11836 17070
rect 11900 13870 11928 19110
rect 11992 16425 12020 19790
rect 12084 19378 12112 19926
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 18902 12112 19314
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11978 16416 12034 16425
rect 11978 16351 12034 16360
rect 12084 16114 12112 18634
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11992 13462 12020 14214
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11900 12646 11928 13398
rect 12084 13258 12112 15438
rect 12176 14958 12204 21422
rect 12544 21418 12572 21558
rect 12532 21412 12584 21418
rect 12716 21412 12768 21418
rect 12532 21354 12584 21360
rect 12636 21372 12716 21400
rect 12636 20806 12664 21372
rect 12716 21354 12768 21360
rect 12820 21010 12848 21655
rect 12900 21616 12952 21622
rect 12900 21558 12952 21564
rect 12912 21418 12940 21558
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12268 19718 12296 19926
rect 12360 19854 12388 20470
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 20233 12480 20334
rect 12438 20224 12494 20233
rect 12438 20159 12494 20168
rect 12530 19952 12586 19961
rect 12530 19887 12586 19896
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12360 19292 12388 19790
rect 12544 19553 12572 19887
rect 12530 19544 12586 19553
rect 12530 19479 12586 19488
rect 12440 19304 12492 19310
rect 12360 19264 12440 19292
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12268 14414 12296 19110
rect 12360 18426 12388 19264
rect 12440 19246 12492 19252
rect 12636 18970 12664 20742
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 19718 12756 20334
rect 12820 20262 12848 20946
rect 13004 20874 13032 20946
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 12808 20256 12860 20262
rect 13544 20256 13596 20262
rect 12860 20216 12940 20244
rect 12808 20198 12860 20204
rect 12912 19922 12940 20216
rect 13544 20198 13596 20204
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12254 14240 12310 14249
rect 12176 13326 12204 14214
rect 12254 14175 12310 14184
rect 12268 13530 12296 14175
rect 12360 13814 12388 18022
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12452 14414 12480 17818
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12452 14074 12480 14350
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12360 13786 12480 13814
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 11898 11928 12582
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 9654 11928 11630
rect 11992 11354 12020 12854
rect 12084 11354 12112 12922
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12070 11248 12126 11257
rect 12070 11183 12126 11192
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11900 8809 11928 9415
rect 11992 8974 12020 10746
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11886 8800 11942 8809
rect 11886 8735 11942 8744
rect 11704 8628 11756 8634
rect 11808 8622 12020 8650
rect 11704 8570 11756 8576
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 6118 11744 7890
rect 11808 7546 11836 8502
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11900 6905 11928 7686
rect 11886 6896 11942 6905
rect 11992 6866 12020 8622
rect 11886 6831 11942 6840
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11808 5930 11836 6190
rect 11486 4236 11652 4264
rect 11716 5902 11836 5930
rect 11244 4072 11296 4078
rect 11486 4060 11514 4236
rect 11244 4014 11296 4020
rect 11348 4032 11514 4060
rect 11612 4072 11664 4078
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10690 3023 10746 3032
rect 10876 3052 10928 3058
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 10704 2446 10732 3023
rect 10876 2994 10928 3000
rect 11072 2854 11100 3402
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11060 2848 11112 2854
rect 11164 2825 11192 2858
rect 11256 2854 11284 3878
rect 11348 3058 11376 4032
rect 11612 4014 11664 4020
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11244 2848 11296 2854
rect 11060 2790 11112 2796
rect 11150 2816 11206 2825
rect 11244 2790 11296 2796
rect 11150 2751 11206 2760
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11440 1329 11468 3334
rect 11624 3233 11652 4014
rect 11716 3670 11744 5902
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 5545 11836 5578
rect 11794 5536 11850 5545
rect 11794 5471 11850 5480
rect 11808 4214 11836 5471
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11610 3224 11666 3233
rect 11610 3159 11666 3168
rect 11624 2446 11652 3159
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11426 1320 11482 1329
rect 11426 1255 11482 1264
rect 10414 54 10548 82
rect 11426 82 11482 480
rect 11532 82 11560 2042
rect 11716 1902 11744 3334
rect 11808 3126 11836 4150
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 2446 11836 2790
rect 11900 2689 11928 6598
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 4146 12020 6054
rect 12084 5302 12112 11183
rect 12176 9654 12204 13262
rect 12268 12986 12296 13262
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12360 12866 12388 13398
rect 12452 13394 12480 13786
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12268 12838 12388 12866
rect 12268 10062 12296 12838
rect 12346 12744 12402 12753
rect 12346 12679 12402 12688
rect 12360 12646 12388 12679
rect 12348 12640 12400 12646
rect 12452 12617 12480 13194
rect 12348 12582 12400 12588
rect 12438 12608 12494 12617
rect 12438 12543 12494 12552
rect 12438 12472 12494 12481
rect 12438 12407 12494 12416
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 12073 12388 12242
rect 12346 12064 12402 12073
rect 12346 11999 12402 12008
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12254 9888 12310 9897
rect 12254 9823 12310 9832
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12268 9489 12296 9823
rect 12254 9480 12310 9489
rect 12254 9415 12310 9424
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 9217 12204 9318
rect 12162 9208 12218 9217
rect 12162 9143 12218 9152
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8294 12204 8774
rect 12268 8430 12296 8910
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7857 12204 8230
rect 12360 8106 12388 11766
rect 12452 11558 12480 12407
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12452 10266 12480 10775
rect 12544 10713 12572 18702
rect 12636 17746 12664 18770
rect 12728 18154 12756 19654
rect 12820 18902 12848 19858
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13266 19272 13322 19281
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 13096 18834 13124 19246
rect 13176 19236 13228 19242
rect 13266 19207 13322 19216
rect 13176 19178 13228 19184
rect 13188 18970 13216 19178
rect 13280 19174 13308 19207
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18204 12848 18566
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12900 18216 12952 18222
rect 12820 18176 12900 18204
rect 12900 18158 12952 18164
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12912 17814 12940 18158
rect 13174 17912 13230 17921
rect 13174 17847 13230 17856
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12636 17542 12664 17682
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 17105 12664 17206
rect 12728 17134 12756 17750
rect 13188 17746 13216 17847
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12820 17241 12848 17614
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 12806 17232 12862 17241
rect 12806 17167 12862 17176
rect 12716 17128 12768 17134
rect 12622 17096 12678 17105
rect 12716 17070 12768 17076
rect 12622 17031 12678 17040
rect 12728 16794 12756 17070
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13188 16969 13216 17002
rect 12806 16960 12862 16969
rect 12806 16895 12862 16904
rect 13174 16960 13230 16969
rect 13174 16895 13230 16904
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12820 16658 12848 16895
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12636 16454 12664 16526
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12636 15638 12664 16390
rect 12820 15910 12848 16594
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12622 15328 12678 15337
rect 12622 15263 12678 15272
rect 12636 11286 12664 15263
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12530 10704 12586 10713
rect 12530 10639 12586 10648
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12268 8078 12388 8106
rect 12162 7848 12218 7857
rect 12162 7783 12218 7792
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 7002 12204 7142
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6322 12204 6938
rect 12268 6458 12296 8078
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12360 7342 12388 7958
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12176 5846 12204 6258
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12084 4049 12112 5034
rect 12268 4690 12296 6394
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12070 4040 12126 4049
rect 12070 3975 12126 3984
rect 12084 3618 12112 3975
rect 11992 3590 12112 3618
rect 11886 2680 11942 2689
rect 11886 2615 11942 2624
rect 11992 2582 12020 3590
rect 12070 3496 12126 3505
rect 12070 3431 12126 3440
rect 12084 3194 12112 3431
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12072 2984 12124 2990
rect 12176 2972 12204 4422
rect 12360 4264 12388 5578
rect 12268 4236 12388 4264
rect 12268 4078 12296 4236
rect 12452 4154 12480 9862
rect 12544 8090 12572 10474
rect 12636 10266 12664 11222
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 10130 12756 15846
rect 12912 15570 12940 15982
rect 13004 15881 13032 16050
rect 13176 15904 13228 15910
rect 12990 15872 13046 15881
rect 13176 15846 13228 15852
rect 12990 15807 13046 15816
rect 13188 15638 13216 15846
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 12900 15564 12952 15570
rect 12820 15524 12900 15552
rect 12820 15366 12848 15524
rect 12900 15506 12952 15512
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12820 15201 12848 15302
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12806 15192 12862 15201
rect 12956 15184 13252 15204
rect 12806 15127 12862 15136
rect 12820 15026 12848 15127
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12820 13734 12848 14554
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12912 13546 12940 13806
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12820 13518 12940 13546
rect 12820 11880 12848 13518
rect 13188 13462 13216 13670
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13280 13326 13308 18702
rect 13372 17270 13400 19858
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13358 16416 13414 16425
rect 13358 16351 13414 16360
rect 13372 14482 13400 16351
rect 13464 15706 13492 19790
rect 13556 19514 13584 20198
rect 13648 20074 13676 22510
rect 13740 20602 13768 23582
rect 13818 23520 13874 23582
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15396 23582 15714 23610
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14002 22944 14058 22953
rect 14002 22879 14058 22888
rect 14016 21146 14044 22879
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13648 20046 13768 20074
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13556 18193 13584 19450
rect 13542 18184 13598 18193
rect 13542 18119 13598 18128
rect 13648 17921 13676 19722
rect 13634 17912 13690 17921
rect 13634 17847 13690 17856
rect 13740 17762 13768 20046
rect 14016 19938 14044 20402
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 13924 19910 14044 19938
rect 13924 19514 13952 19910
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13832 19145 13860 19314
rect 13912 19236 13964 19242
rect 14016 19224 14044 19790
rect 14200 19786 14228 20198
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19514 14136 19654
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13964 19196 14044 19224
rect 13912 19178 13964 19184
rect 13818 19136 13874 19145
rect 13818 19071 13874 19080
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 13832 18086 13860 18634
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13648 17734 13768 17762
rect 13832 17746 13860 18022
rect 13820 17740 13872 17746
rect 13556 17338 13584 17682
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13556 17066 13584 17274
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13358 13968 13414 13977
rect 13358 13903 13414 13912
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 13174 12608 13230 12617
rect 13174 12543 13230 12552
rect 12990 12472 13046 12481
rect 12990 12407 13046 12416
rect 13004 12374 13032 12407
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 13188 12220 13216 12543
rect 13188 12192 13308 12220
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 13280 11880 13308 12192
rect 12820 11852 12940 11880
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 11665 12848 11698
rect 12806 11656 12862 11665
rect 12806 11591 12862 11600
rect 12912 11286 12940 11852
rect 13188 11852 13308 11880
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11354 13124 11562
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12820 10674 12848 11222
rect 13188 11082 13216 11852
rect 13372 11286 13400 13903
rect 13464 12442 13492 15438
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13464 11762 13492 12378
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13358 11112 13414 11121
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 12990 10704 13046 10713
rect 12808 10668 12860 10674
rect 12990 10639 13046 10648
rect 12808 10610 12860 10616
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12808 10192 12860 10198
rect 12912 10169 12940 10474
rect 12808 10134 12860 10140
rect 12898 10160 12954 10169
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12622 10024 12678 10033
rect 12622 9959 12678 9968
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12360 4126 12480 4154
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12124 2944 12204 2972
rect 12072 2926 12124 2932
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12084 2106 12112 2926
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12176 2650 12204 2790
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 11716 649 11744 1838
rect 11702 640 11758 649
rect 11702 575 11758 584
rect 11426 54 11560 82
rect 12268 82 12296 3878
rect 12360 2922 12388 4126
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12544 1873 12572 7754
rect 12636 6458 12664 9959
rect 12728 9722 12756 10066
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12716 9376 12768 9382
rect 12820 9364 12848 10134
rect 12898 10095 12954 10104
rect 12768 9336 12848 9364
rect 12716 9318 12768 9324
rect 12728 9178 12756 9318
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12912 9058 12940 10095
rect 13004 9994 13032 10639
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10266 13216 10474
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13188 9840 13216 10066
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 12728 9030 12940 9058
rect 12728 8498 12756 9030
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12728 5846 12756 8230
rect 12820 6769 12848 8910
rect 13188 8820 13216 9744
rect 13280 8974 13308 11086
rect 13358 11047 13414 11056
rect 13372 11014 13400 11047
rect 13360 11008 13412 11014
rect 13464 10985 13492 11290
rect 13360 10950 13412 10956
rect 13450 10976 13506 10985
rect 13450 10911 13506 10920
rect 13450 10840 13506 10849
rect 13360 10804 13412 10810
rect 13450 10775 13506 10784
rect 13360 10746 13412 10752
rect 13372 10305 13400 10746
rect 13464 10742 13492 10775
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13358 10296 13414 10305
rect 13358 10231 13414 10240
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13358 10160 13414 10169
rect 13358 10095 13414 10104
rect 13372 9178 13400 10095
rect 13464 10062 13492 10202
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13556 9874 13584 16526
rect 13648 14482 13676 17734
rect 13820 17682 13872 17688
rect 13728 17672 13780 17678
rect 13924 17626 13952 18838
rect 14016 18329 14044 19196
rect 14108 18873 14136 19450
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14200 18970 14228 19314
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14094 18864 14150 18873
rect 14094 18799 14150 18808
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18358 14136 18566
rect 14096 18352 14148 18358
rect 14002 18320 14058 18329
rect 14096 18294 14148 18300
rect 14002 18255 14058 18264
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14002 17912 14058 17921
rect 14002 17847 14058 17856
rect 13728 17614 13780 17620
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13740 12889 13768 17614
rect 13832 17598 13952 17626
rect 13832 16266 13860 17598
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13924 16454 13952 16662
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13832 16238 13952 16266
rect 13818 16144 13874 16153
rect 13818 16079 13874 16088
rect 13726 12880 13782 12889
rect 13636 12844 13688 12850
rect 13726 12815 13782 12824
rect 13636 12786 13688 12792
rect 13648 12170 13676 12786
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 10198 13676 11494
rect 13740 11354 13768 12242
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13832 10520 13860 16079
rect 13924 14618 13952 16238
rect 14016 16017 14044 17847
rect 14108 17785 14136 18022
rect 14094 17776 14150 17785
rect 14094 17711 14150 17720
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14002 16008 14058 16017
rect 14002 15943 14058 15952
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14016 14498 14044 14758
rect 13924 14470 14044 14498
rect 13924 13818 13952 14470
rect 13924 13790 14044 13818
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12986 13952 13330
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13924 12442 13952 12718
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13924 11801 13952 12106
rect 13910 11792 13966 11801
rect 13910 11727 13966 11736
rect 13910 11112 13966 11121
rect 13910 11047 13966 11056
rect 13924 10810 13952 11047
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14016 10713 14044 13790
rect 14108 13138 14136 16934
rect 14200 14890 14228 18634
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14200 14618 14228 14826
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14200 14074 14228 14554
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14186 13968 14242 13977
rect 14186 13903 14242 13912
rect 14200 13870 14228 13903
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14108 13110 14228 13138
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14108 12782 14136 12922
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12646 14136 12718
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14108 11626 14136 12582
rect 14200 11898 14228 13110
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14186 11656 14242 11665
rect 14096 11620 14148 11626
rect 14186 11591 14242 11600
rect 14096 11562 14148 11568
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14108 10810 14136 11154
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14002 10704 14058 10713
rect 14002 10639 14058 10648
rect 13832 10492 13952 10520
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13464 9846 13584 9874
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13188 8792 13308 8820
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 13082 8392 13138 8401
rect 13082 8327 13138 8336
rect 13176 8356 13228 8362
rect 13096 8022 13124 8327
rect 13176 8298 13228 8304
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13188 7954 13216 8298
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 12898 7440 12954 7449
rect 12898 7375 12954 7384
rect 12806 6760 12862 6769
rect 12806 6695 12862 6704
rect 12912 6644 12940 7375
rect 12820 6616 12940 6644
rect 12820 6168 12848 6616
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 12992 6180 13044 6186
rect 12820 6140 12992 6168
rect 12992 6122 13044 6128
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4758 12664 4966
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12636 4486 12664 4694
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12728 4154 12756 5782
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12820 5370 12848 5646
rect 13096 5642 13124 5714
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12820 5137 12848 5306
rect 12806 5128 12862 5137
rect 12806 5063 12862 5072
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 12900 5024 12952 5030
rect 12806 4992 12862 5001
rect 12900 4966 12952 4972
rect 12806 4927 12862 4936
rect 12820 4622 12848 4927
rect 12808 4616 12860 4622
rect 12912 4593 12940 4966
rect 13096 4690 13124 5034
rect 13280 4758 13308 8792
rect 13372 8634 13400 9114
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13358 8256 13414 8265
rect 13358 8191 13414 8200
rect 13372 8022 13400 8191
rect 13464 8090 13492 9846
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6186 13400 7142
rect 13464 6934 13492 7686
rect 13556 7002 13584 9687
rect 13648 9042 13676 9930
rect 13924 9722 13952 10492
rect 14002 10296 14058 10305
rect 14002 10231 14058 10240
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13740 9178 13768 9658
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13648 8634 13676 8842
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13740 8537 13768 8774
rect 13832 8634 13860 9279
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13726 8528 13782 8537
rect 13636 8492 13688 8498
rect 13726 8463 13782 8472
rect 13636 8434 13688 8440
rect 13648 8022 13676 8434
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13648 7546 13676 7958
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13556 6458 13584 6734
rect 13740 6662 13768 7346
rect 13820 7200 13872 7206
rect 13924 7188 13952 8978
rect 14016 8945 14044 10231
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14108 9081 14136 10134
rect 14094 9072 14150 9081
rect 14094 9007 14150 9016
rect 14002 8936 14058 8945
rect 14002 8871 14058 8880
rect 14094 8800 14150 8809
rect 14094 8735 14150 8744
rect 14108 8129 14136 8735
rect 14094 8120 14150 8129
rect 14004 8084 14056 8090
rect 14094 8055 14150 8064
rect 14004 8026 14056 8032
rect 13872 7160 13952 7188
rect 13820 7142 13872 7148
rect 13832 6934 13860 7142
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13910 6896 13966 6905
rect 13910 6831 13966 6840
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13464 6186 13492 6394
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12808 4558 12860 4564
rect 12898 4584 12954 4593
rect 12636 4126 12756 4154
rect 12820 4154 12848 4558
rect 12898 4519 12954 4528
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 13280 4214 13308 4694
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13268 4208 13320 4214
rect 12820 4126 12940 4154
rect 13268 4150 13320 4156
rect 13372 4146 13400 4422
rect 12636 3369 12664 4126
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 12728 3097 12756 4014
rect 12912 3738 12940 4126
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13174 3632 13230 3641
rect 13174 3567 13230 3576
rect 13188 3534 13216 3567
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 13280 3126 13308 3674
rect 13268 3120 13320 3126
rect 12714 3088 12770 3097
rect 13268 3062 13320 3068
rect 12714 3023 12770 3032
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12636 2553 12664 2926
rect 12622 2544 12678 2553
rect 12622 2479 12678 2488
rect 12728 2281 12756 3023
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12898 2544 12954 2553
rect 12714 2272 12770 2281
rect 12714 2207 12770 2216
rect 12530 1864 12586 1873
rect 12530 1799 12586 1808
rect 12820 1737 12848 2518
rect 13372 2514 13400 2926
rect 12898 2479 12954 2488
rect 13360 2508 13412 2514
rect 12912 2446 12940 2479
rect 13360 2450 13412 2456
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13464 2310 13492 5646
rect 13556 5409 13584 5850
rect 13542 5400 13598 5409
rect 13542 5335 13598 5344
rect 13648 5030 13676 6326
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5642 13768 5850
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13726 4720 13782 4729
rect 13726 4655 13782 4664
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13556 3720 13584 4490
rect 13648 4282 13676 4558
rect 13740 4486 13768 4655
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13648 3738 13676 3946
rect 13636 3732 13688 3738
rect 13556 3692 13636 3720
rect 13556 3058 13584 3692
rect 13636 3674 13688 3680
rect 13726 3632 13782 3641
rect 13726 3567 13782 3576
rect 13740 3534 13768 3567
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13556 2310 13584 2858
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 12806 1728 12862 1737
rect 12806 1663 12862 1672
rect 12438 82 12494 480
rect 12268 54 12494 82
rect 9402 0 9458 54
rect 10414 0 10470 54
rect 11426 0 11482 54
rect 12438 0 12494 54
rect 13450 82 13506 480
rect 13648 82 13676 3402
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13740 2922 13768 2994
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13832 2854 13860 6734
rect 13924 6322 13952 6831
rect 14016 6798 14044 8026
rect 14200 7970 14228 11591
rect 14292 8974 14320 22442
rect 14462 22128 14518 22137
rect 14462 22063 14518 22072
rect 14476 19394 14504 22063
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14568 20398 14596 21082
rect 14752 20806 14780 22986
rect 15016 21412 15068 21418
rect 14936 21372 15016 21400
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20398 14780 20742
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14568 19786 14596 20334
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14384 19366 14504 19394
rect 14384 13394 14412 19366
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14476 18222 14504 19178
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18290 14596 18566
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17746 14504 18158
rect 14752 18154 14780 19110
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14476 16794 14504 17070
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14370 13016 14426 13025
rect 14370 12951 14426 12960
rect 14384 12918 14412 12951
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14384 10033 14412 12718
rect 14370 10024 14426 10033
rect 14370 9959 14426 9968
rect 14476 9602 14504 16526
rect 14568 15745 14596 17478
rect 14660 17105 14688 17682
rect 14646 17096 14702 17105
rect 14646 17031 14702 17040
rect 14554 15736 14610 15745
rect 14554 15671 14610 15680
rect 14660 15570 14688 17031
rect 14844 16522 14872 20946
rect 14936 20942 14964 21372
rect 15016 21354 15068 21360
rect 15120 21350 15148 23530
rect 15396 21690 15424 23582
rect 15658 23520 15714 23582
rect 17328 23582 17554 23610
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 15660 22296 15712 22302
rect 15660 22238 15712 22244
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15108 21344 15160 21350
rect 15014 21312 15070 21321
rect 15108 21286 15160 21292
rect 15014 21247 15070 21256
rect 15028 21146 15056 21247
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14936 18902 14964 20878
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 15028 19281 15056 19858
rect 15014 19272 15070 19281
rect 15014 19207 15070 19216
rect 14924 18896 14976 18902
rect 14924 18838 14976 18844
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 15028 18329 15056 18770
rect 15014 18320 15070 18329
rect 15014 18255 15070 18264
rect 15028 18086 15056 18255
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15028 17921 15056 18022
rect 15014 17912 15070 17921
rect 15014 17847 15070 17856
rect 14924 17808 14976 17814
rect 15120 17785 15148 21286
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15212 20233 15240 20334
rect 15198 20224 15254 20233
rect 15198 20159 15254 20168
rect 15198 20088 15254 20097
rect 15198 20023 15254 20032
rect 15212 18834 15240 20023
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15212 18426 15240 18770
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 14924 17750 14976 17756
rect 15106 17776 15162 17785
rect 14936 17649 14964 17750
rect 15106 17711 15162 17720
rect 15108 17672 15160 17678
rect 14922 17640 14978 17649
rect 15108 17614 15160 17620
rect 14922 17575 14978 17584
rect 14922 17504 14978 17513
rect 14922 17439 14978 17448
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14738 15328 14794 15337
rect 14738 15263 14794 15272
rect 14752 14550 14780 15263
rect 14740 14544 14792 14550
rect 14660 14504 14740 14532
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 14074 14596 14418
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14568 13977 14596 14010
rect 14554 13968 14610 13977
rect 14554 13903 14610 13912
rect 14554 13560 14610 13569
rect 14554 13495 14610 13504
rect 14568 13274 14596 13495
rect 14660 13433 14688 14504
rect 14740 14486 14792 14492
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13734 14780 14214
rect 14844 14074 14872 15574
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14646 13424 14702 13433
rect 14646 13359 14702 13368
rect 14568 13246 14780 13274
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14568 10674 14596 13126
rect 14660 12102 14688 13126
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11558 14688 12038
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 10849 14688 11494
rect 14646 10840 14702 10849
rect 14646 10775 14702 10784
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14384 9574 14504 9602
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14108 7942 14228 7970
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13924 3602 13952 4218
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14016 2650 14044 6394
rect 14108 4826 14136 7942
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7721 14228 7822
rect 14186 7712 14242 7721
rect 14186 7647 14242 7656
rect 14292 7274 14320 8434
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14292 6390 14320 7210
rect 14384 6934 14412 9574
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9178 14504 9454
rect 14568 9178 14596 10610
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14660 10266 14688 10474
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14660 9722 14688 10202
rect 14752 10130 14780 13246
rect 14844 11762 14872 13806
rect 14936 12714 14964 17439
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 14890 15056 16934
rect 15120 16794 15148 17614
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16046 15148 16390
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15120 14958 15148 15506
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 15120 14793 15148 14894
rect 15106 14784 15162 14793
rect 15106 14719 15162 14728
rect 15212 14385 15240 18022
rect 15198 14376 15254 14385
rect 15198 14311 15254 14320
rect 15304 14074 15332 21082
rect 15488 21078 15516 21830
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15580 21418 15608 21626
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15580 21146 15608 21354
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15396 20058 15424 20266
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15488 19854 15516 21014
rect 15672 20262 15700 22238
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15764 20942 15792 21354
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 15934 21040 15990 21049
rect 15934 20975 15990 20984
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15396 16998 15424 19450
rect 15476 19168 15528 19174
rect 15580 19156 15608 19858
rect 15672 19174 15700 19926
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15856 19310 15884 19722
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15528 19128 15608 19156
rect 15660 19168 15712 19174
rect 15476 19110 15528 19116
rect 15660 19110 15712 19116
rect 15488 18426 15516 19110
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15488 17746 15516 18362
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15488 17066 15516 17682
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14922 12472 14978 12481
rect 14922 12407 14978 12416
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14936 11354 14964 12407
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15028 11665 15056 12310
rect 15014 11656 15070 11665
rect 15014 11591 15070 11600
rect 15028 11558 15056 11591
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 10198 14872 10610
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 15014 10160 15070 10169
rect 14740 10124 14792 10130
rect 15014 10095 15070 10104
rect 14740 10066 14792 10072
rect 14738 10024 14794 10033
rect 14738 9959 14794 9968
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14752 9654 14780 9959
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 8265 14504 8842
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14462 8256 14518 8265
rect 14462 8191 14518 8200
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14370 6488 14426 6497
rect 14370 6423 14426 6432
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14200 5574 14228 5782
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14108 4486 14136 4762
rect 14200 4758 14228 5510
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14094 4312 14150 4321
rect 14094 4247 14150 4256
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14108 241 14136 4247
rect 14292 4078 14320 6122
rect 14384 5409 14412 6423
rect 14476 6186 14504 7958
rect 14568 7410 14596 8502
rect 14660 8022 14688 8910
rect 14752 8090 14780 9590
rect 15028 9489 15056 10095
rect 15120 9926 15148 13874
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15014 9480 15070 9489
rect 15014 9415 15070 9424
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14844 7750 14872 9046
rect 15120 8974 15148 9386
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 7750 14964 8366
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14660 7478 14688 7686
rect 14738 7576 14794 7585
rect 14738 7511 14794 7520
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14568 5409 14596 7346
rect 14660 7274 14688 7414
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14370 5400 14426 5409
rect 14370 5335 14426 5344
rect 14554 5400 14610 5409
rect 14554 5335 14610 5344
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 4826 14412 5170
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14370 4584 14426 4593
rect 14370 4519 14426 4528
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14384 3942 14412 4519
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 3176 14320 3334
rect 14372 3188 14424 3194
rect 14292 3148 14372 3176
rect 14372 3130 14424 3136
rect 14476 2990 14504 4626
rect 14660 4282 14688 6326
rect 14752 5914 14780 7511
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14844 5642 14872 7686
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14844 4214 14872 4422
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14752 3738 14780 4082
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14752 3058 14780 3674
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14476 2553 14504 2926
rect 14752 2650 14780 2994
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14462 2544 14518 2553
rect 14462 2479 14518 2488
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14752 2310 14780 2450
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14476 2038 14504 2246
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 14752 1873 14780 2246
rect 14738 1864 14794 1873
rect 14738 1799 14794 1808
rect 14094 232 14150 241
rect 14094 167 14150 176
rect 13450 54 13676 82
rect 14462 60 14518 480
rect 14936 105 14964 7686
rect 15028 7449 15056 8774
rect 15120 8634 15148 8910
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15014 7440 15070 7449
rect 15014 7375 15070 7384
rect 15014 7304 15070 7313
rect 15014 7239 15070 7248
rect 15028 7002 15056 7239
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15028 6458 15056 6666
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15120 6254 15148 6870
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15028 5098 15056 5714
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 15028 4010 15056 5034
rect 15108 4276 15160 4282
rect 15212 4264 15240 13126
rect 15304 12782 15332 13126
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10985 15332 11086
rect 15290 10976 15346 10985
rect 15290 10911 15346 10920
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10441 15332 10542
rect 15290 10432 15346 10441
rect 15290 10367 15346 10376
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15304 6662 15332 9862
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15396 5574 15424 16730
rect 15580 16658 15608 17818
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 16250 15608 16594
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15488 14346 15516 16118
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 15570 15608 15914
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15580 15366 15608 15506
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 15162 15608 15302
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15580 13802 15608 14418
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 8634 15516 13670
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 12782 15608 13330
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15566 12472 15622 12481
rect 15566 12407 15622 12416
rect 15580 12374 15608 12407
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15580 10713 15608 11698
rect 15566 10704 15622 10713
rect 15566 10639 15622 10648
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15488 5386 15516 8434
rect 15580 7857 15608 9318
rect 15672 8090 15700 15438
rect 15764 14618 15792 19178
rect 15856 18970 15884 19246
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15856 17202 15884 17546
rect 15948 17202 15976 20975
rect 16040 19718 16068 21286
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16132 20398 16160 20742
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16040 18902 16068 19654
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16026 18728 16082 18737
rect 16026 18663 16082 18672
rect 16040 18630 16068 18663
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16026 17232 16082 17241
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15936 17196 15988 17202
rect 16026 17167 16082 17176
rect 15936 17138 15988 17144
rect 16040 17134 16068 17167
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 15948 16046 15976 17002
rect 16040 16658 16068 17070
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16040 16250 16068 16594
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15948 15366 15976 15982
rect 16040 15706 16068 16186
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15844 14952 15896 14958
rect 15948 14940 15976 15302
rect 15896 14912 15976 14940
rect 15844 14894 15896 14900
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 11218 15792 14418
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15764 10266 15792 11154
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15566 7848 15622 7857
rect 15566 7783 15622 7792
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 7313 15608 7346
rect 15566 7304 15622 7313
rect 15566 7239 15622 7248
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15396 5358 15516 5386
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15160 4236 15240 4264
rect 15108 4218 15160 4224
rect 15304 4185 15332 4558
rect 15290 4176 15346 4185
rect 15290 4111 15346 4120
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15028 3097 15056 3946
rect 15304 3126 15332 3946
rect 15292 3120 15344 3126
rect 15014 3088 15070 3097
rect 15292 3062 15344 3068
rect 15014 3023 15070 3032
rect 15028 2904 15056 3023
rect 15108 2916 15160 2922
rect 15028 2876 15108 2904
rect 15108 2858 15160 2864
rect 15396 1970 15424 5358
rect 15474 5128 15530 5137
rect 15474 5063 15530 5072
rect 15488 3738 15516 5063
rect 15580 5012 15608 7142
rect 15672 5930 15700 7890
rect 15764 7177 15792 8774
rect 15856 7954 15884 14758
rect 15948 14346 15976 14912
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 14249 15976 14282
rect 15934 14240 15990 14249
rect 15934 14175 15990 14184
rect 15934 14104 15990 14113
rect 15934 14039 15990 14048
rect 15948 13530 15976 14039
rect 16040 13870 16068 14486
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16026 13696 16082 13705
rect 16026 13631 16082 13640
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16040 13410 16068 13631
rect 15948 13382 16068 13410
rect 15948 12306 15976 13382
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12714 16068 13126
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16026 12608 16082 12617
rect 16026 12543 16082 12552
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15948 11150 15976 12242
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15948 9518 15976 10066
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 16040 8378 16068 12543
rect 16132 12442 16160 19994
rect 16224 15162 16252 22578
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 16960 21418 16988 22102
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 21185 16804 21286
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16762 21176 16818 21185
rect 16956 21168 17252 21188
rect 16762 21111 16818 21120
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16684 20262 16712 20878
rect 16776 20330 16804 21014
rect 16946 20904 17002 20913
rect 16946 20839 17002 20848
rect 16960 20534 16988 20839
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16316 17882 16344 18158
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16132 11762 16160 12378
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 11354 16160 11562
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16132 10810 16160 11290
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16132 10538 16160 10746
rect 16224 10674 16252 14894
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16224 10266 16252 10610
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16316 9874 16344 17002
rect 16408 16590 16436 18702
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16224 9846 16344 9874
rect 15948 8022 15976 8366
rect 16040 8350 16160 8378
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15856 7546 15884 7890
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15750 7168 15806 7177
rect 15750 7103 15806 7112
rect 15842 6216 15898 6225
rect 15842 6151 15898 6160
rect 15672 5902 15792 5930
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15672 5370 15700 5782
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15764 5302 15792 5902
rect 15752 5296 15804 5302
rect 15658 5264 15714 5273
rect 15752 5238 15804 5244
rect 15658 5199 15714 5208
rect 15672 5166 15700 5199
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15580 4984 15700 5012
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15580 3602 15608 4422
rect 15672 3777 15700 4984
rect 15750 3904 15806 3913
rect 15750 3839 15806 3848
rect 15658 3768 15714 3777
rect 15658 3703 15714 3712
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15580 2922 15608 3538
rect 15672 3369 15700 3703
rect 15764 3670 15792 3839
rect 15856 3777 15884 6151
rect 15948 4457 15976 7686
rect 16040 6866 16068 8230
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16040 5846 16068 6054
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 16132 5302 16160 8350
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16118 5128 16174 5137
rect 16118 5063 16174 5072
rect 16132 5030 16160 5063
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16118 4720 16174 4729
rect 16224 4690 16252 9846
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16408 9674 16436 15914
rect 16500 14550 16528 19314
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16592 14482 16620 19926
rect 16684 19718 16712 20198
rect 16776 19961 16804 20266
rect 16762 19952 16818 19961
rect 16868 19922 16896 20470
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16762 19887 16818 19896
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19514 16712 19654
rect 16868 19514 16896 19858
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 16960 18426 16988 18770
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 18080 16724 18086
rect 16776 18057 16804 18090
rect 16672 18022 16724 18028
rect 16762 18048 16818 18057
rect 16684 16046 16712 18022
rect 16762 17983 16818 17992
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 11898 16528 14214
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16592 13190 16620 13806
rect 16684 13569 16712 15302
rect 16776 14113 16804 17478
rect 16868 15366 16896 18294
rect 17236 18154 17264 18770
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 16960 16114 16988 16594
rect 17236 16250 17264 16594
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 16946 15464 17002 15473
rect 16946 15399 17002 15408
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16960 15162 16988 15399
rect 17052 15201 17080 15506
rect 17038 15192 17094 15201
rect 16948 15156 17000 15162
rect 17038 15127 17094 15136
rect 16948 15098 17000 15104
rect 16856 14816 16908 14822
rect 17052 14804 17080 15127
rect 16908 14776 17080 14804
rect 16856 14758 16908 14764
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 17328 14618 17356 23582
rect 17498 23520 17554 23582
rect 19338 23588 19394 24000
rect 21178 23610 21234 24000
rect 23018 23610 23074 24000
rect 19338 23536 19340 23588
rect 19392 23536 19394 23588
rect 19338 23520 19394 23536
rect 20916 23582 21234 23610
rect 19352 23499 19380 23520
rect 19156 22908 19208 22914
rect 19156 22850 19208 22856
rect 17590 22808 17646 22817
rect 17590 22743 17646 22752
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17420 19174 17448 19858
rect 17512 19310 17540 21286
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17420 18902 17448 19110
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16762 14104 16818 14113
rect 16762 14039 16818 14048
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16670 13560 16726 13569
rect 16670 13495 16726 13504
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16684 12646 16712 13398
rect 16776 12850 16804 13942
rect 16868 13734 16896 14486
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16960 13938 16988 14282
rect 17328 13938 17356 14350
rect 17420 14006 17448 18702
rect 17512 17746 17540 19246
rect 17604 17882 17632 22743
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17866 22536 17922 22545
rect 17866 22471 17922 22480
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17512 17338 17540 17682
rect 17696 17354 17724 20742
rect 17788 19446 17816 21422
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17604 17326 17724 17354
rect 17788 17338 17816 19382
rect 17880 18086 17908 22471
rect 17868 18080 17920 18086
rect 17866 18048 17868 18057
rect 17920 18048 17922 18057
rect 17866 17983 17922 17992
rect 17776 17332 17828 17338
rect 17604 16454 17632 17326
rect 17776 17274 17828 17280
rect 17788 17134 17816 17274
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17512 15570 17540 16186
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17512 15162 17540 15506
rect 17696 15502 17724 16050
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16868 13512 16896 13670
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 16868 13484 16988 13512
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16592 10656 16620 12582
rect 16684 11354 16712 12582
rect 16776 12374 16804 12786
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16762 11384 16818 11393
rect 16672 11348 16724 11354
rect 16762 11319 16818 11328
rect 16672 11290 16724 11296
rect 16592 10628 16712 10656
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 10266 16620 10474
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16316 9450 16344 9658
rect 16408 9646 16528 9674
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16316 9178 16344 9386
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16408 7546 16436 7958
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16408 6934 16436 7482
rect 16500 7154 16528 9646
rect 16592 9110 16620 10202
rect 16580 9104 16632 9110
rect 16684 9081 16712 10628
rect 16776 10266 16804 11319
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16868 10130 16896 13126
rect 16960 12986 16988 13484
rect 17328 13326 17356 13874
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 17512 12374 17540 14894
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17236 11801 17264 12242
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17222 11792 17278 11801
rect 17222 11727 17278 11736
rect 17236 11694 17264 11727
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 16960 10577 16988 10950
rect 16946 10568 17002 10577
rect 16946 10503 17002 10512
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 17130 10160 17186 10169
rect 16856 10124 16908 10130
rect 17130 10095 17186 10104
rect 16856 10066 16908 10072
rect 16946 10024 17002 10033
rect 16856 9988 16908 9994
rect 16946 9959 17002 9968
rect 16856 9930 16908 9936
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16580 9046 16632 9052
rect 16670 9072 16726 9081
rect 16592 8634 16620 9046
rect 16670 9007 16726 9016
rect 16670 8936 16726 8945
rect 16670 8871 16726 8880
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16592 8022 16620 8570
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16592 7274 16620 7822
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16500 7126 16620 7154
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16408 6458 16436 6870
rect 16500 6798 16528 6938
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16592 6458 16620 7126
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16408 6186 16436 6394
rect 16578 6216 16634 6225
rect 16396 6180 16448 6186
rect 16578 6151 16634 6160
rect 16396 6122 16448 6128
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16316 5545 16344 5714
rect 16302 5536 16358 5545
rect 16302 5471 16358 5480
rect 16408 5352 16436 6122
rect 16486 5944 16542 5953
rect 16592 5914 16620 6151
rect 16486 5879 16542 5888
rect 16580 5908 16632 5914
rect 16500 5778 16528 5879
rect 16580 5850 16632 5856
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16316 5324 16436 5352
rect 16316 4758 16344 5324
rect 16394 5264 16450 5273
rect 16394 5199 16450 5208
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16118 4655 16174 4664
rect 16212 4684 16264 4690
rect 15934 4448 15990 4457
rect 15934 4383 15990 4392
rect 15842 3768 15898 3777
rect 16132 3738 16160 4655
rect 16212 4626 16264 4632
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16224 4146 16252 4490
rect 16316 4282 16344 4694
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16304 4004 16356 4010
rect 16224 3964 16304 3992
rect 16224 3777 16252 3964
rect 16304 3946 16356 3952
rect 16210 3768 16266 3777
rect 15842 3703 15898 3712
rect 16120 3732 16172 3738
rect 16210 3703 16266 3712
rect 16120 3674 16172 3680
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 16224 3602 16252 3703
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 15750 3496 15806 3505
rect 15750 3431 15806 3440
rect 16026 3496 16082 3505
rect 16026 3431 16082 3440
rect 15764 3398 15792 3431
rect 15752 3392 15804 3398
rect 15658 3360 15714 3369
rect 15752 3334 15804 3340
rect 15658 3295 15714 3304
rect 15658 3224 15714 3233
rect 15658 3159 15714 3168
rect 15672 3126 15700 3159
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 15568 2372 15620 2378
rect 15672 2360 15700 3062
rect 15620 2332 15700 2360
rect 15568 2314 15620 2320
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 13450 0 13506 54
rect 14462 8 14464 60
rect 14516 8 14518 60
rect 14922 96 14978 105
rect 14922 31 14978 40
rect 15474 82 15530 480
rect 15764 82 15792 3062
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15856 2514 15884 2858
rect 16040 2825 16068 3431
rect 16132 3097 16160 3538
rect 16118 3088 16174 3097
rect 16118 3023 16174 3032
rect 16132 2990 16160 3023
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16120 2848 16172 2854
rect 16026 2816 16082 2825
rect 16120 2790 16172 2796
rect 16026 2751 16082 2760
rect 16132 2582 16160 2790
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 15474 54 15792 82
rect 16224 82 16252 2042
rect 16408 921 16436 5199
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16500 3942 16528 5034
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16592 3534 16620 5510
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16684 2582 16712 8871
rect 16776 5710 16804 9862
rect 16868 9042 16896 9930
rect 16960 9518 16988 9959
rect 17144 9722 17172 10095
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17328 9586 17356 10950
rect 17420 10418 17448 12174
rect 17512 11898 17540 12310
rect 17604 12238 17632 15438
rect 17788 15366 17816 16390
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17498 11656 17554 11665
rect 17604 11626 17632 12038
rect 17498 11591 17554 11600
rect 17592 11620 17644 11626
rect 17512 11200 17540 11591
rect 17592 11562 17644 11568
rect 17696 11268 17724 15302
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17788 13190 17816 14350
rect 17880 13870 17908 16662
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17880 13002 17908 13670
rect 17788 12974 17908 13002
rect 17788 12306 17816 12974
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17880 12102 17908 12650
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11354 17908 12038
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17776 11280 17828 11286
rect 17696 11240 17776 11268
rect 17776 11222 17828 11228
rect 17592 11212 17644 11218
rect 17512 11172 17592 11200
rect 17592 11154 17644 11160
rect 17604 10810 17632 11154
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17420 10390 17540 10418
rect 17406 10296 17462 10305
rect 17406 10231 17462 10240
rect 17420 10198 17448 10231
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 17222 9072 17278 9081
rect 16856 9036 16908 9042
rect 17222 9007 17278 9016
rect 16856 8978 16908 8984
rect 16868 8634 16896 8978
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 17236 8430 17264 9007
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17328 8362 17356 8774
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6361 16896 7142
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 16854 6352 16910 6361
rect 16854 6287 16910 6296
rect 16868 5914 16896 6287
rect 17328 6118 17356 7482
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17420 5710 17448 10134
rect 17512 5710 17540 10390
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9586 17632 10066
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17696 7002 17724 10678
rect 17972 10674 18000 22646
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18064 21078 18092 21558
rect 18156 21486 18184 21558
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18340 21418 18368 21898
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18616 21350 18644 21558
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 18512 21072 18564 21078
rect 18512 21014 18564 21020
rect 18524 20602 18552 21014
rect 18708 20806 18736 21286
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18420 20392 18472 20398
rect 18142 20360 18198 20369
rect 18142 20295 18198 20304
rect 18340 20352 18420 20380
rect 18156 20262 18184 20295
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18340 19786 18368 20352
rect 18420 20334 18472 20340
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18156 18970 18184 19178
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18248 18834 18276 19178
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18340 18222 18368 19722
rect 18524 19446 18552 20538
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18064 14618 18092 17818
rect 18156 15706 18184 18158
rect 18340 17882 18368 18158
rect 18432 18086 18460 18770
rect 18524 18358 18552 19382
rect 18616 19174 18644 19858
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18340 16794 18368 17818
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18248 15570 18276 15914
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18156 14890 18184 15370
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18156 14226 18184 14826
rect 18248 14278 18276 14826
rect 18064 14198 18184 14226
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18064 13988 18092 14198
rect 18248 14074 18276 14214
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18064 13960 18184 13988
rect 18050 13832 18106 13841
rect 18050 13767 18106 13776
rect 18064 13530 18092 13767
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18156 12442 18184 13960
rect 18248 13802 18276 14010
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18248 12918 18276 13398
rect 18340 13258 18368 13670
rect 18432 13297 18460 18022
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18524 15065 18552 17818
rect 18616 17746 18644 19110
rect 18604 17740 18656 17746
rect 18656 17700 18736 17728
rect 18604 17682 18656 17688
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18510 15056 18566 15065
rect 18510 14991 18566 15000
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18524 13530 18552 14486
rect 18616 13569 18644 17478
rect 18708 17338 18736 17700
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18708 16658 18736 17002
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18708 16250 18736 16594
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 14006 18736 15982
rect 18800 15337 18828 21490
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18892 16794 18920 20402
rect 18984 20262 19012 21014
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18984 16182 19012 20198
rect 19076 17814 19104 22034
rect 19064 17808 19116 17814
rect 19064 17750 19116 17756
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18786 15328 18842 15337
rect 18786 15263 18842 15272
rect 18892 14958 18920 15506
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 14414 18828 14826
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18602 13560 18658 13569
rect 18512 13524 18564 13530
rect 18602 13495 18658 13504
rect 18512 13466 18564 13472
rect 18512 13320 18564 13326
rect 18418 13288 18474 13297
rect 18328 13252 18380 13258
rect 18512 13262 18564 13268
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18418 13223 18474 13232
rect 18328 13194 18380 13200
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18340 12442 18368 13194
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18248 11626 18276 11834
rect 18432 11762 18460 13126
rect 18524 12170 18552 13262
rect 18616 13025 18644 13262
rect 18602 13016 18658 13025
rect 18602 12951 18658 12960
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10130 17816 10406
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17788 9722 17816 10066
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17880 9518 17908 10134
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17788 8294 17816 9114
rect 17880 8498 17908 9318
rect 17972 8974 18000 9862
rect 18064 9432 18092 10202
rect 18156 9722 18184 11562
rect 18616 11558 18644 12951
rect 18800 12850 18828 14350
rect 18878 13968 18934 13977
rect 18878 13903 18934 13912
rect 18892 13394 18920 13903
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 11014 18644 11086
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18248 10538 18276 10950
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18248 9926 18276 10474
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18248 9450 18276 9862
rect 18340 9761 18368 10746
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 18326 9752 18382 9761
rect 18326 9687 18382 9696
rect 18432 9568 18460 9959
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18340 9540 18460 9568
rect 18144 9444 18196 9450
rect 18064 9404 18144 9432
rect 18144 9386 18196 9392
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18050 9208 18106 9217
rect 18050 9143 18106 9152
rect 18064 9110 18092 9143
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 8090 17816 8230
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7200 17828 7206
rect 17880 7188 17908 7958
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17828 7160 17908 7188
rect 17960 7200 18012 7206
rect 17776 7142 17828 7148
rect 17960 7142 18012 7148
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 17788 6934 17816 7142
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17788 6458 17816 6734
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17590 6352 17646 6361
rect 17590 6287 17646 6296
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 5030 16896 5102
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16762 4856 16818 4865
rect 16868 4826 16896 4966
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 16762 4791 16818 4800
rect 16856 4820 16908 4826
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16394 912 16450 921
rect 16394 847 16450 856
rect 16486 82 16542 480
rect 16776 134 16804 4791
rect 16856 4762 16908 4768
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16868 3670 16896 4218
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16868 2854 16896 3606
rect 17328 3126 17356 5578
rect 17512 5302 17540 5646
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 17420 4298 17448 5238
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17512 5001 17540 5034
rect 17604 5030 17632 6287
rect 17682 5944 17738 5953
rect 17682 5879 17738 5888
rect 17696 5642 17724 5879
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17592 5024 17644 5030
rect 17498 4992 17554 5001
rect 17592 4966 17644 4972
rect 17498 4927 17554 4936
rect 17696 4706 17724 5102
rect 17788 4826 17816 5782
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17880 5681 17908 5714
rect 17866 5672 17922 5681
rect 17866 5607 17922 5616
rect 17866 5400 17922 5409
rect 17866 5335 17922 5344
rect 17880 5302 17908 5335
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17696 4678 17816 4706
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17604 4298 17632 4558
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17420 4270 17632 4298
rect 17420 4146 17448 4270
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17406 3904 17462 3913
rect 17406 3839 17462 3848
rect 17420 3738 17448 3839
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17512 2961 17540 2994
rect 17498 2952 17554 2961
rect 17498 2887 17554 2896
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2378 16896 2790
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 17406 2680 17462 2689
rect 17328 2650 17406 2666
rect 17316 2644 17406 2650
rect 17368 2638 17406 2644
rect 17696 2650 17724 4422
rect 17788 4154 17816 4678
rect 17880 4593 17908 4762
rect 17866 4584 17922 4593
rect 17866 4519 17922 4528
rect 17788 4126 17908 4154
rect 17880 3194 17908 4126
rect 17972 4010 18000 7142
rect 18064 7002 18092 7822
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18156 6905 18184 9386
rect 18340 8922 18368 9540
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18248 8894 18368 8922
rect 18142 6896 18198 6905
rect 18142 6831 18198 6840
rect 18248 6746 18276 8894
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18340 7585 18368 8774
rect 18432 8362 18460 9386
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18326 7576 18382 7585
rect 18326 7511 18382 7520
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 18340 7002 18368 7210
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18156 6718 18276 6746
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 18064 3738 18092 6054
rect 18156 4486 18184 6718
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6186 18276 6598
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18248 5914 18276 6122
rect 18432 6118 18460 8298
rect 18524 6458 18552 9862
rect 18616 9586 18644 10950
rect 18708 9994 18736 12582
rect 18800 11762 18828 12786
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18892 10810 18920 11222
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18800 10198 18828 10474
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18340 5817 18368 5850
rect 18326 5808 18382 5817
rect 18326 5743 18382 5752
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18340 5234 18368 5578
rect 18432 5273 18460 6054
rect 18418 5264 18474 5273
rect 18328 5228 18380 5234
rect 18418 5199 18474 5208
rect 18328 5170 18380 5176
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18524 4321 18552 6054
rect 18510 4312 18566 4321
rect 18510 4247 18566 4256
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18156 3913 18184 3946
rect 18142 3904 18198 3913
rect 18142 3839 18198 3848
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18064 3602 18092 3674
rect 18248 3670 18276 3946
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17880 2922 17908 3130
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17406 2615 17462 2624
rect 17684 2644 17736 2650
rect 17316 2586 17368 2592
rect 17684 2586 17736 2592
rect 17222 2544 17278 2553
rect 17222 2479 17278 2488
rect 17236 2446 17264 2479
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 18064 1465 18092 3334
rect 18156 2922 18184 3334
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18248 2514 18276 2858
rect 18340 2854 18368 3538
rect 18432 3108 18460 4082
rect 18616 3176 18644 9046
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18708 8514 18736 8842
rect 18800 8634 18828 9998
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18892 9450 18920 9930
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18892 8514 18920 8570
rect 18708 8486 18920 8514
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18708 5545 18736 6394
rect 18694 5536 18750 5545
rect 18694 5471 18750 5480
rect 18708 4154 18736 5471
rect 18800 4321 18828 7686
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18892 6390 18920 7278
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18984 6089 19012 15914
rect 19076 15745 19104 17274
rect 19168 16182 19196 22850
rect 19248 22840 19300 22846
rect 19248 22782 19300 22788
rect 19260 18426 19288 22782
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 19062 15736 19118 15745
rect 19062 15671 19118 15680
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 13814 19104 15438
rect 19168 14074 19196 15506
rect 19260 14385 19288 18022
rect 19352 17338 19380 22714
rect 20916 22234 20944 23582
rect 21178 23520 21234 23582
rect 22664 23582 23074 23610
rect 21730 22944 21786 22953
rect 21730 22879 21786 22888
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20444 22024 20496 22030
rect 20258 21992 20314 22001
rect 20444 21966 20496 21972
rect 20258 21927 20314 21936
rect 19798 21448 19854 21457
rect 19798 21383 19854 21392
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 20505 19472 21286
rect 19430 20496 19486 20505
rect 19430 20431 19486 20440
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19536 19174 19564 20266
rect 19616 20256 19668 20262
rect 19668 20233 19748 20244
rect 19668 20224 19762 20233
rect 19668 20216 19706 20224
rect 19616 20198 19668 20204
rect 19706 20159 19762 20168
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19444 17542 19472 18770
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19536 16998 19564 19110
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19352 15881 19380 15914
rect 19338 15872 19394 15881
rect 19338 15807 19394 15816
rect 19338 15736 19394 15745
rect 19444 15706 19472 16526
rect 19338 15671 19394 15680
rect 19432 15700 19484 15706
rect 19246 14376 19302 14385
rect 19246 14311 19302 14320
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19352 13814 19380 15671
rect 19432 15642 19484 15648
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 14550 19472 15302
rect 19536 14958 19564 16934
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19076 13786 19196 13814
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19076 9382 19104 10134
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9178 19104 9318
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 19076 8430 19104 8978
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19076 7478 19104 8366
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 19076 7274 19104 7414
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19076 6390 19104 6870
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 18970 6080 19026 6089
rect 18970 6015 19026 6024
rect 19076 5846 19104 6326
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 5166 19012 5510
rect 19076 5302 19104 5782
rect 19168 5574 19196 13786
rect 19260 13786 19380 13814
rect 19260 12714 19288 13786
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19260 8498 19288 9114
rect 19352 9110 19380 13670
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19444 12986 19472 13330
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19444 12306 19472 12922
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11898 19472 12242
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19444 8809 19472 9318
rect 19536 9042 19564 12038
rect 19628 11898 19656 18702
rect 19812 18465 19840 21383
rect 20076 20528 20128 20534
rect 20128 20488 20208 20516
rect 20076 20470 20128 20476
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19798 18456 19854 18465
rect 19708 18420 19760 18426
rect 19798 18391 19854 18400
rect 19708 18362 19760 18368
rect 19720 17762 19748 18362
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19812 17882 19840 18226
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19720 17734 19840 17762
rect 19812 16046 19840 17734
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19614 11520 19670 11529
rect 19614 11455 19670 11464
rect 19628 10810 19656 11455
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19628 9110 19656 10746
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19616 8968 19668 8974
rect 19536 8916 19616 8922
rect 19536 8910 19668 8916
rect 19536 8894 19656 8910
rect 19430 8800 19486 8809
rect 19430 8735 19486 8744
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 8090 19380 8230
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19260 7313 19288 7414
rect 19246 7304 19302 7313
rect 19246 7239 19302 7248
rect 19260 6254 19288 7239
rect 19352 6322 19380 7686
rect 19444 7342 19472 7890
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19536 6186 19564 8894
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19628 6730 19656 8774
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19260 5409 19288 6054
rect 19246 5400 19302 5409
rect 19246 5335 19302 5344
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18984 4554 19012 5102
rect 19076 4622 19104 5238
rect 19154 4856 19210 4865
rect 19154 4791 19210 4800
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18878 4448 18934 4457
rect 18878 4383 18934 4392
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18708 4146 18828 4154
rect 18708 4140 18840 4146
rect 18708 4126 18788 4140
rect 18788 4082 18840 4088
rect 18892 4049 18920 4383
rect 18970 4312 19026 4321
rect 19076 4282 19104 4558
rect 18970 4247 19026 4256
rect 19064 4276 19116 4282
rect 18984 4185 19012 4247
rect 19064 4218 19116 4224
rect 18970 4176 19026 4185
rect 19026 4134 19104 4162
rect 18970 4111 19026 4120
rect 18984 4078 19012 4111
rect 18972 4072 19024 4078
rect 18878 4040 18934 4049
rect 18788 4004 18840 4010
rect 19076 4049 19104 4134
rect 18972 4014 19024 4020
rect 19062 4040 19118 4049
rect 18878 3975 18934 3984
rect 19062 3975 19118 3984
rect 18788 3946 18840 3952
rect 18800 3890 18828 3946
rect 19076 3890 19104 3975
rect 18800 3862 19104 3890
rect 19168 3738 19196 4791
rect 19444 4758 19472 6054
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19536 4434 19564 5510
rect 19628 4729 19656 5646
rect 19614 4720 19670 4729
rect 19614 4655 19670 4664
rect 19444 4406 19564 4434
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19444 4154 19472 4406
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19260 4126 19472 4154
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18708 3369 18736 3538
rect 18694 3360 18750 3369
rect 18694 3295 18750 3304
rect 18616 3148 18828 3176
rect 18512 3120 18564 3126
rect 18432 3080 18512 3108
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18432 2582 18460 3080
rect 18512 3062 18564 3068
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18512 2576 18564 2582
rect 18512 2518 18564 2524
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18524 2378 18552 2518
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18050 1456 18106 1465
rect 18050 1391 18106 1400
rect 16224 54 16542 82
rect 16764 128 16816 134
rect 16764 70 16816 76
rect 17406 128 17462 480
rect 17406 76 17408 128
rect 17460 76 17462 128
rect 14462 0 14518 8
rect 15474 0 15530 54
rect 16486 0 16542 54
rect 17406 0 17462 76
rect 18418 82 18474 480
rect 18708 82 18736 2586
rect 18800 2310 18828 3148
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 18878 2680 18934 2689
rect 18878 2615 18934 2624
rect 18892 2582 18920 2615
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 19076 2514 19104 2994
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 19260 2378 19288 4126
rect 19536 4049 19564 4218
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 19628 3942 19656 4422
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19432 3528 19484 3534
rect 19536 3516 19564 3878
rect 19720 3738 19748 15846
rect 19904 15201 19932 20198
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19996 19310 20024 19858
rect 20074 19408 20130 19417
rect 20074 19343 20130 19352
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 20088 18426 20116 19343
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19996 15638 20024 17818
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19890 15192 19946 15201
rect 19890 15127 19946 15136
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19996 14550 20024 14894
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19812 13870 19840 14350
rect 19996 14328 20024 14486
rect 20088 14396 20116 17750
rect 20180 15570 20208 20488
rect 20272 18358 20300 21927
rect 20456 19310 20484 21966
rect 21454 21856 21510 21865
rect 20956 21788 21252 21808
rect 21454 21791 21510 21800
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20810 21720 20866 21729
rect 20956 21712 21252 21732
rect 20810 21655 20866 21664
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20272 16425 20300 17070
rect 20258 16416 20314 16425
rect 20258 16351 20314 16360
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20180 14929 20208 15302
rect 20166 14920 20222 14929
rect 20166 14855 20222 14864
rect 20272 14550 20300 16186
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 20088 14368 20300 14396
rect 19996 14300 20208 14328
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19812 12306 19840 13806
rect 19982 13152 20038 13161
rect 19982 13087 20038 13096
rect 19890 12336 19946 12345
rect 19800 12300 19852 12306
rect 19890 12271 19946 12280
rect 19800 12242 19852 12248
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19812 11626 19840 11766
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19812 11354 19840 11562
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19904 11286 19932 12271
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19890 10840 19946 10849
rect 19890 10775 19946 10784
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19812 9042 19840 9454
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19812 8634 19840 8978
rect 19904 8838 19932 10775
rect 19996 10130 20024 13087
rect 20180 12782 20208 14300
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20180 12442 20208 12718
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20180 11354 20208 11698
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20272 10810 20300 14368
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19996 10033 20024 10066
rect 19982 10024 20038 10033
rect 20168 9988 20220 9994
rect 19982 9959 20038 9968
rect 20088 9948 20168 9976
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19812 7886 19840 8298
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19798 7440 19854 7449
rect 19798 7375 19854 7384
rect 19812 5302 19840 7375
rect 19904 7274 19932 8502
rect 19996 8022 20024 9522
rect 19984 8016 20036 8022
rect 19984 7958 20036 7964
rect 19996 7410 20024 7958
rect 20088 7546 20116 9948
rect 20168 9930 20220 9936
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20166 9208 20222 9217
rect 20166 9143 20222 9152
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19892 7268 19944 7274
rect 19892 7210 19944 7216
rect 19904 7002 19932 7210
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20088 6390 20116 6598
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 19800 5296 19852 5302
rect 19852 5256 19932 5284
rect 19800 5238 19852 5244
rect 19904 4457 19932 5256
rect 20074 4720 20130 4729
rect 19996 4690 20074 4706
rect 19984 4684 20074 4690
rect 20036 4678 20074 4684
rect 20180 4690 20208 9143
rect 20272 7410 20300 9318
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20364 6458 20392 19110
rect 20442 18184 20498 18193
rect 20548 18154 20576 20266
rect 20640 19514 20668 21519
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20640 18154 20668 18702
rect 20732 18329 20760 21422
rect 20824 21078 20852 21655
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 20824 20602 20852 21014
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20824 19174 20852 19858
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20824 18358 20852 18838
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 20812 18352 20864 18358
rect 20718 18320 20774 18329
rect 20812 18294 20864 18300
rect 20718 18255 20774 18264
rect 20442 18119 20498 18128
rect 20536 18148 20588 18154
rect 20456 14346 20484 18119
rect 20536 18090 20588 18096
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 14521 20576 15302
rect 20640 15094 20668 18090
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20824 16998 20852 17682
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16114 20760 16662
rect 21284 16590 21312 20878
rect 21376 20330 21404 21014
rect 21468 20602 21496 21791
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21468 20398 21496 20538
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21364 19712 21416 19718
rect 21560 19700 21588 20810
rect 21638 20768 21694 20777
rect 21638 20703 21694 20712
rect 21652 20058 21680 20703
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21416 19672 21588 19700
rect 21364 19654 21416 19660
rect 21376 18766 21404 19654
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21546 18592 21602 18601
rect 21546 18527 21602 18536
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21468 17610 21496 17682
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21362 17504 21418 17513
rect 21362 17439 21418 17448
rect 21376 17338 21404 17439
rect 21468 17338 21496 17546
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20732 15609 20760 16050
rect 20824 15910 20852 16526
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 20718 15600 20774 15609
rect 20718 15535 20774 15544
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20824 15162 20852 15506
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20720 14544 20772 14550
rect 20534 14512 20590 14521
rect 20720 14486 20772 14492
rect 20534 14447 20590 14456
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20732 13530 20760 14486
rect 20824 14482 20852 15098
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 14074 20852 14418
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20824 13161 20852 13330
rect 20916 13297 20944 13466
rect 21008 13394 21036 13874
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 20902 13288 20958 13297
rect 20902 13223 20958 13232
rect 20810 13152 20866 13161
rect 20810 13087 20866 13096
rect 20824 12986 20852 13087
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20456 10742 20484 12378
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20548 10538 20576 12718
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20442 10432 20498 10441
rect 20442 10367 20498 10376
rect 20456 10266 20484 10367
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20456 8498 20484 10202
rect 20548 9654 20576 10202
rect 20640 9897 20668 11290
rect 20732 11200 20760 12650
rect 21284 12345 21312 14282
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 13870 21404 14214
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21270 12336 21326 12345
rect 20812 12300 20864 12306
rect 21270 12271 21326 12280
rect 20812 12242 20864 12248
rect 20824 11898 20852 12242
rect 21376 12152 21404 13806
rect 21468 12918 21496 15846
rect 21560 12986 21588 18527
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21456 12300 21508 12306
rect 21652 12288 21680 15982
rect 21744 15162 21772 22879
rect 22664 20534 22692 23582
rect 23018 23520 23074 23582
rect 22652 20528 22704 20534
rect 22652 20470 22704 20476
rect 21822 19816 21878 19825
rect 21822 19751 21878 19760
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21744 14958 21772 15098
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21836 14804 21864 19751
rect 23572 19304 23624 19310
rect 21914 19272 21970 19281
rect 23572 19246 23624 19252
rect 21914 19207 21970 19216
rect 21456 12242 21508 12248
rect 21560 12260 21680 12288
rect 21744 14776 21864 14804
rect 21284 12124 21404 12152
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20812 11212 20864 11218
rect 20732 11172 20812 11200
rect 20812 11154 20864 11160
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20626 9888 20682 9897
rect 20626 9823 20682 9832
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20442 8256 20498 8265
rect 20442 8191 20498 8200
rect 20456 7954 20484 8191
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20548 7342 20576 8774
rect 20732 8072 20760 10950
rect 20824 10810 20852 11154
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9722 20852 10066
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 21086 9480 21142 9489
rect 20996 9444 21048 9450
rect 21086 9415 21142 9424
rect 20996 9386 21048 9392
rect 21008 9110 21036 9386
rect 21100 9110 21128 9415
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21100 8820 21128 9046
rect 21284 8945 21312 12124
rect 21362 12064 21418 12073
rect 21362 11999 21418 12008
rect 21376 11898 21404 11999
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21468 11830 21496 12242
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21270 8936 21326 8945
rect 21270 8871 21326 8880
rect 20824 8792 21128 8820
rect 20824 8634 20852 8792
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 20640 8044 20760 8072
rect 20812 8084 20864 8090
rect 20640 7478 20668 8044
rect 20812 8026 20864 8032
rect 20718 7984 20774 7993
rect 20718 7919 20774 7928
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20732 6798 20760 7919
rect 20824 7546 20852 8026
rect 21008 8022 21036 8502
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 21284 7886 21312 8230
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20812 6928 20864 6934
rect 20812 6870 20864 6876
rect 20720 6792 20772 6798
rect 20626 6760 20682 6769
rect 20720 6734 20772 6740
rect 20626 6695 20682 6704
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20074 4655 20130 4664
rect 20168 4684 20220 4690
rect 19984 4626 20036 4632
rect 20168 4626 20220 4632
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19890 4448 19946 4457
rect 19890 4383 19946 4392
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19982 4176 20038 4185
rect 19812 4010 19840 4150
rect 19982 4111 20038 4120
rect 19800 4004 19852 4010
rect 19800 3946 19852 3952
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19536 3488 19656 3516
rect 19904 3505 19932 3878
rect 19432 3470 19484 3476
rect 19444 3058 19472 3470
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19536 2922 19564 3334
rect 19628 3097 19656 3488
rect 19890 3496 19946 3505
rect 19890 3431 19946 3440
rect 19614 3088 19670 3097
rect 19614 3023 19670 3032
rect 19892 3052 19944 3058
rect 19996 3040 20024 4111
rect 20088 3097 20116 4558
rect 19944 3012 20024 3040
rect 20074 3088 20130 3097
rect 20074 3023 20130 3032
rect 19892 2994 19944 3000
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 19352 1193 19380 2790
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 19800 2304 19852 2310
rect 19904 2281 19932 2994
rect 19800 2246 19852 2252
rect 19890 2272 19946 2281
rect 19338 1184 19394 1193
rect 19338 1119 19394 1128
rect 19720 513 19748 2246
rect 19706 504 19762 513
rect 18418 54 18736 82
rect 19430 82 19486 480
rect 19706 439 19762 448
rect 19812 82 19840 2246
rect 19890 2207 19946 2216
rect 19430 54 19840 82
rect 20088 82 20116 3023
rect 20272 2514 20300 5578
rect 20456 5030 20484 5782
rect 20640 5302 20668 6695
rect 20718 6488 20774 6497
rect 20718 6423 20774 6432
rect 20732 6254 20760 6423
rect 20824 6390 20852 6870
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20824 5370 20852 6326
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 20534 5128 20590 5137
rect 20534 5063 20590 5072
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 20364 4593 20392 4626
rect 20350 4584 20406 4593
rect 20350 4519 20406 4528
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20272 785 20300 2450
rect 20258 776 20314 785
rect 20258 711 20314 720
rect 20364 649 20392 4014
rect 20456 3670 20484 4966
rect 20548 3738 20576 5063
rect 20994 4992 21050 5001
rect 20994 4927 21050 4936
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20640 3738 20668 4626
rect 20824 4282 20852 4694
rect 21008 4622 21036 4927
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 21284 4154 21312 7686
rect 21376 5914 21404 11698
rect 21454 10024 21510 10033
rect 21454 9959 21510 9968
rect 21468 6458 21496 9959
rect 21560 9450 21588 12260
rect 21638 12200 21694 12209
rect 21638 12135 21694 12144
rect 21652 12102 21680 12135
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21744 11898 21772 14776
rect 21928 13814 21956 19207
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21836 13786 21956 13814
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21744 11694 21772 11834
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21744 10810 21772 11154
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21744 10130 21772 10746
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21744 9654 21772 10066
rect 21732 9648 21784 9654
rect 21732 9590 21784 9596
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21560 8566 21588 9386
rect 21730 9072 21786 9081
rect 21730 9007 21786 9016
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21548 8560 21600 8566
rect 21548 8502 21600 8508
rect 21652 7857 21680 8842
rect 21744 8430 21772 9007
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21638 7848 21694 7857
rect 21638 7783 21694 7792
rect 21652 7290 21680 7783
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21560 7262 21680 7290
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21560 6390 21588 7262
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21192 4126 21312 4154
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20732 1329 20760 3470
rect 20824 2854 20852 3606
rect 21192 3534 21220 4126
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 21376 2938 21404 5850
rect 21652 5846 21680 6666
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 21652 4758 21680 5782
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21652 4282 21680 4694
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21744 4185 21772 7686
rect 21730 4176 21786 4185
rect 21730 4111 21786 4120
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21284 2910 21404 2938
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 21284 2514 21312 2910
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20718 1320 20774 1329
rect 20718 1255 20774 1264
rect 20350 640 20406 649
rect 20350 575 20406 584
rect 20442 82 20498 480
rect 20088 54 20498 82
rect 21376 66 21404 2790
rect 21744 2417 21772 3878
rect 21836 2650 21864 13786
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 10577 21956 13126
rect 22020 11393 22048 14214
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22112 12986 22140 13330
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22006 11384 22062 11393
rect 22006 11319 22062 11328
rect 22006 10976 22062 10985
rect 22006 10911 22062 10920
rect 21914 10568 21970 10577
rect 21914 10503 21970 10512
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21928 9178 21956 9862
rect 22020 9722 22048 10911
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 9353 22048 9386
rect 22006 9344 22062 9353
rect 22006 9279 22062 9288
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21928 8634 21956 8774
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 22006 8528 22062 8537
rect 22006 8463 22062 8472
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21928 4622 21956 7142
rect 22020 6390 22048 8463
rect 22112 8362 22140 10406
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22100 6656 22152 6662
rect 22204 6633 22232 18158
rect 23584 16969 23612 19246
rect 23570 16960 23626 16969
rect 23492 16918 23570 16946
rect 22742 14240 22798 14249
rect 22742 14175 22798 14184
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22296 12753 22324 13126
rect 22282 12744 22338 12753
rect 22282 12679 22338 12688
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 11257 22324 12038
rect 22282 11248 22338 11257
rect 22282 11183 22338 11192
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 9897 22324 10950
rect 22374 10296 22430 10305
rect 22374 10231 22430 10240
rect 22282 9888 22338 9897
rect 22282 9823 22338 9832
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22100 6598 22152 6604
rect 22190 6624 22246 6633
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 22112 5710 22140 6598
rect 22190 6559 22246 6568
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22296 5137 22324 7686
rect 22282 5128 22338 5137
rect 22282 5063 22338 5072
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21928 3534 21956 4218
rect 22020 3641 22048 4966
rect 22006 3632 22062 3641
rect 22006 3567 22062 3576
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22112 2825 22140 2858
rect 22098 2816 22154 2825
rect 22098 2751 22154 2760
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21730 2408 21786 2417
rect 21730 2343 21786 2352
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 21744 2009 21772 2246
rect 22204 2038 22232 4966
rect 22388 4282 22416 10231
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22480 4729 22508 8230
rect 22466 4720 22522 4729
rect 22466 4655 22522 4664
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22192 2032 22244 2038
rect 21730 2000 21786 2009
rect 22192 1974 22244 1980
rect 21730 1935 21786 1944
rect 21454 96 21510 480
rect 22296 377 22324 3334
rect 22282 368 22338 377
rect 22282 303 22338 312
rect 18418 0 18474 54
rect 19430 0 19486 54
rect 20442 0 20498 54
rect 21364 60 21416 66
rect 21364 2 21416 8
rect 21454 0 21510 40
rect 22466 82 22522 480
rect 22572 82 22600 13194
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22664 5545 22692 12854
rect 22756 11801 22784 14175
rect 23492 14074 23520 16918
rect 23570 16895 23626 16904
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23584 13705 23612 13942
rect 23570 13696 23626 13705
rect 23570 13631 23626 13640
rect 22742 11792 22798 11801
rect 22742 11727 22798 11736
rect 22650 5536 22706 5545
rect 22650 5471 22706 5480
rect 22756 5166 22784 11727
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22466 54 22600 82
rect 23216 82 23244 7346
rect 23492 3890 23520 10678
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23584 7177 23612 7414
rect 23570 7168 23626 7177
rect 23570 7103 23626 7112
rect 23570 3904 23626 3913
rect 23492 3862 23570 3890
rect 23570 3839 23626 3848
rect 23478 82 23534 480
rect 23216 54 23534 82
rect 22466 0 22522 54
rect 23478 0 23534 54
<< via2 >>
rect 846 23160 902 23216
rect 386 21528 442 21584
rect 202 20576 258 20632
rect 18 20168 74 20224
rect 110 17040 166 17096
rect 110 16224 166 16280
rect 18 14592 74 14648
rect 18 12552 74 12608
rect 18 11872 74 11928
rect 18 11464 74 11520
rect 294 17312 350 17368
rect 110 7384 166 7440
rect 18 5072 74 5128
rect 478 19896 534 19952
rect 386 12824 442 12880
rect 754 22616 810 22672
rect 570 17448 626 17504
rect 662 17312 718 17368
rect 662 16632 718 16688
rect 662 16496 718 16552
rect 570 9832 626 9888
rect 938 18264 994 18320
rect 846 17992 902 18048
rect 846 16768 902 16824
rect 754 14456 810 14512
rect 1398 22888 1454 22944
rect 1306 22344 1362 22400
rect 1214 16904 1270 16960
rect 1122 13252 1178 13288
rect 1122 13232 1124 13252
rect 1124 13232 1176 13252
rect 1176 13232 1178 13252
rect 1674 22752 1730 22808
rect 1582 21256 1638 21312
rect 1490 18264 1546 18320
rect 1398 15000 1454 15056
rect 1214 12280 1270 12336
rect 1214 10920 1270 10976
rect 1214 9152 1270 9208
rect 1582 15136 1638 15192
rect 1582 14320 1638 14376
rect 1398 11056 1454 11112
rect 2318 21256 2374 21312
rect 2226 21120 2282 21176
rect 2134 20168 2190 20224
rect 2134 20032 2190 20088
rect 2226 19760 2282 19816
rect 2042 19080 2098 19136
rect 2042 16632 2098 16688
rect 2226 17448 2282 17504
rect 2226 17040 2282 17096
rect 2778 20712 2834 20768
rect 2502 19624 2558 19680
rect 2410 17176 2466 17232
rect 2226 16224 2282 16280
rect 1950 14184 2006 14240
rect 2318 16088 2374 16144
rect 2226 14864 2282 14920
rect 1582 10648 1638 10704
rect 1490 9288 1546 9344
rect 1214 8880 1270 8936
rect 1122 8336 1178 8392
rect 1398 8064 1454 8120
rect 1766 12552 1822 12608
rect 1766 8744 1822 8800
rect 1950 12008 2006 12064
rect 2134 12688 2190 12744
rect 2134 9832 2190 9888
rect 2134 9696 2190 9752
rect 2042 9152 2098 9208
rect 1950 8472 2006 8528
rect 1674 6568 1730 6624
rect 1582 6296 1638 6352
rect 1490 6024 1546 6080
rect 1398 3712 1454 3768
rect 2134 8608 2190 8664
rect 2134 7792 2190 7848
rect 1858 7384 1914 7440
rect 2042 6704 2098 6760
rect 2410 14048 2466 14104
rect 3698 23024 3754 23080
rect 3054 21392 3110 21448
rect 2962 19760 3018 19816
rect 2686 18400 2742 18456
rect 2686 17992 2742 18048
rect 2778 15136 2834 15192
rect 3238 19488 3294 19544
rect 3146 19080 3202 19136
rect 3238 15952 3294 16008
rect 3146 15816 3202 15872
rect 2594 11600 2650 11656
rect 2502 11192 2558 11248
rect 2778 13640 2834 13696
rect 2962 14184 3018 14240
rect 2686 10648 2742 10704
rect 2686 10240 2742 10296
rect 2870 10104 2926 10160
rect 2594 9424 2650 9480
rect 2594 8336 2650 8392
rect 2502 8064 2558 8120
rect 2410 7656 2466 7712
rect 2226 5888 2282 5944
rect 1674 3168 1730 3224
rect 2686 8200 2742 8256
rect 2686 6432 2742 6488
rect 2686 6024 2742 6080
rect 2962 9696 3018 9752
rect 3238 15136 3294 15192
rect 3330 14728 3386 14784
rect 3606 20576 3662 20632
rect 3974 20032 4030 20088
rect 3882 18944 3938 19000
rect 3514 13776 3570 13832
rect 3698 15408 3754 15464
rect 4894 22072 4950 22128
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4434 20984 4490 21040
rect 4710 20712 4766 20768
rect 4710 20032 4766 20088
rect 4526 19352 4582 19408
rect 5446 20848 5502 20904
rect 5354 20712 5410 20768
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4802 19352 4858 19408
rect 4066 17720 4122 17776
rect 3698 14184 3754 14240
rect 3146 12416 3202 12472
rect 3054 9016 3110 9072
rect 3238 9424 3294 9480
rect 3238 8880 3294 8936
rect 2962 7928 3018 7984
rect 3238 8200 3294 8256
rect 3146 7520 3202 7576
rect 2962 7112 3018 7168
rect 3054 6840 3110 6896
rect 2870 6160 2926 6216
rect 2686 4256 2742 4312
rect 2318 3984 2374 4040
rect 2410 3032 2466 3088
rect 2686 3576 2742 3632
rect 2594 3440 2650 3496
rect 2318 2896 2374 2952
rect 570 1536 626 1592
rect 294 40 350 96
rect 3422 12688 3478 12744
rect 3422 9152 3478 9208
rect 3422 7384 3478 7440
rect 3422 7112 3478 7168
rect 3698 8608 3754 8664
rect 3882 13504 3938 13560
rect 4342 18536 4398 18592
rect 4342 17720 4398 17776
rect 4250 16904 4306 16960
rect 4250 14864 4306 14920
rect 4158 12416 4214 12472
rect 4802 18944 4858 19000
rect 5354 19216 5410 19272
rect 4710 18400 4766 18456
rect 4434 15408 4490 15464
rect 4434 14048 4490 14104
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4894 16904 4950 16960
rect 5262 16904 5318 16960
rect 5814 18808 5870 18864
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4986 16088 5042 16144
rect 5354 15408 5410 15464
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 5078 14592 5134 14648
rect 4618 13368 4674 13424
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4986 13912 5042 13968
rect 4710 13232 4766 13288
rect 4342 12008 4398 12064
rect 4342 11872 4398 11928
rect 3974 10784 4030 10840
rect 3974 10512 4030 10568
rect 3882 8744 3938 8800
rect 3698 8064 3754 8120
rect 3514 4528 3570 4584
rect 3422 4120 3478 4176
rect 3238 3984 3294 4040
rect 3146 1808 3202 1864
rect 2318 1672 2374 1728
rect 4250 11736 4306 11792
rect 4158 9832 4214 9888
rect 4158 9424 4214 9480
rect 3974 7112 4030 7168
rect 3974 6704 4030 6760
rect 3974 6432 4030 6488
rect 3882 6160 3938 6216
rect 4342 10240 4398 10296
rect 4526 11872 4582 11928
rect 4526 10648 4582 10704
rect 5354 13504 5410 13560
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4802 12824 4858 12880
rect 4986 12688 5042 12744
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4894 11464 4950 11520
rect 4710 10512 4766 10568
rect 4434 9832 4490 9888
rect 4250 8744 4306 8800
rect 4434 9172 4490 9208
rect 4434 9152 4436 9172
rect 4436 9152 4488 9172
rect 4488 9152 4490 9172
rect 4434 8608 4490 8664
rect 4250 8200 4306 8256
rect 4158 7112 4214 7168
rect 4158 6296 4214 6352
rect 3882 5752 3938 5808
rect 4066 5616 4122 5672
rect 3974 4664 4030 4720
rect 4158 5072 4214 5128
rect 4434 6160 4490 6216
rect 4434 4664 4490 4720
rect 5262 11464 5318 11520
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4894 10512 4950 10568
rect 4710 10104 4766 10160
rect 4618 9832 4674 9888
rect 4894 9968 4950 10024
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4986 9560 5042 9616
rect 5170 9560 5226 9616
rect 4894 9424 4950 9480
rect 4986 9152 5042 9208
rect 4710 5480 4766 5536
rect 5262 9016 5318 9072
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 5446 12960 5502 13016
rect 5630 12688 5686 12744
rect 6642 22752 6698 22808
rect 7010 21664 7066 21720
rect 6550 20168 6606 20224
rect 6274 19080 6330 19136
rect 6458 18400 6514 18456
rect 6090 16768 6146 16824
rect 5998 16632 6054 16688
rect 6182 16632 6238 16688
rect 5814 13096 5870 13152
rect 5630 12416 5686 12472
rect 5354 7792 5410 7848
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4894 6704 4950 6760
rect 5170 6704 5226 6760
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 5170 5752 5226 5808
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4710 4800 4766 4856
rect 4158 4120 4214 4176
rect 4434 4120 4490 4176
rect 4158 3576 4214 3632
rect 3698 3032 3754 3088
rect 3606 2352 3662 2408
rect 3330 1128 3386 1184
rect 4066 2624 4122 2680
rect 5262 5208 5318 5264
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 4802 2488 4858 2544
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 5814 11872 5870 11928
rect 5722 11056 5778 11112
rect 5906 10376 5962 10432
rect 5722 9832 5778 9888
rect 5814 9696 5870 9752
rect 5630 7792 5686 7848
rect 5814 6160 5870 6216
rect 5538 3984 5594 4040
rect 5538 2760 5594 2816
rect 4618 176 4674 232
rect 5722 3576 5778 3632
rect 6642 18400 6698 18456
rect 6550 16496 6606 16552
rect 6642 15816 6698 15872
rect 6550 14728 6606 14784
rect 6550 14220 6552 14240
rect 6552 14220 6604 14240
rect 6604 14220 6606 14240
rect 6550 14184 6606 14220
rect 6182 12824 6238 12880
rect 6090 10104 6146 10160
rect 6090 9696 6146 9752
rect 5998 8880 6054 8936
rect 6274 12008 6330 12064
rect 6274 8744 6330 8800
rect 6182 7928 6238 7984
rect 6182 7520 6238 7576
rect 5998 7112 6054 7168
rect 5998 4936 6054 4992
rect 5906 4392 5962 4448
rect 5906 3576 5962 3632
rect 6274 6296 6330 6352
rect 6182 5616 6238 5672
rect 6090 4256 6146 4312
rect 5630 720 5686 776
rect 6366 3440 6422 3496
rect 7010 20304 7066 20360
rect 6826 19624 6882 19680
rect 7010 17720 7066 17776
rect 6918 16496 6974 16552
rect 7010 16224 7066 16280
rect 6826 15680 6882 15736
rect 6734 10648 6790 10704
rect 6734 10376 6790 10432
rect 6642 10104 6698 10160
rect 7010 13912 7066 13968
rect 7654 22888 7710 22944
rect 7838 22888 7894 22944
rect 7378 22616 7434 22672
rect 7562 22616 7618 22672
rect 8206 22480 8262 22536
rect 7378 21936 7434 21992
rect 7654 21120 7710 21176
rect 7378 20576 7434 20632
rect 7838 20032 7894 20088
rect 7194 17584 7250 17640
rect 7378 17720 7434 17776
rect 7286 16360 7342 16416
rect 7286 14456 7342 14512
rect 7470 16904 7526 16960
rect 7470 15272 7526 15328
rect 7470 15136 7526 15192
rect 6550 7792 6606 7848
rect 6550 7112 6606 7168
rect 6642 5752 6698 5808
rect 6642 4800 6698 4856
rect 6734 4256 6790 4312
rect 7102 7928 7158 7984
rect 7010 6976 7066 7032
rect 8666 22480 8722 22536
rect 8298 22072 8354 22128
rect 8390 20712 8446 20768
rect 7838 18400 7894 18456
rect 7838 18028 7840 18048
rect 7840 18028 7892 18048
rect 7892 18028 7894 18048
rect 7838 17992 7894 18028
rect 7838 14728 7894 14784
rect 7838 14592 7894 14648
rect 7746 11736 7802 11792
rect 8298 17720 8354 17776
rect 8206 16224 8262 16280
rect 8114 13504 8170 13560
rect 8022 13368 8078 13424
rect 7654 10920 7710 10976
rect 7654 10784 7710 10840
rect 7470 9016 7526 9072
rect 7562 8880 7618 8936
rect 7286 7384 7342 7440
rect 6458 3304 6514 3360
rect 7286 6060 7288 6080
rect 7288 6060 7340 6080
rect 7340 6060 7342 6080
rect 7286 6024 7342 6060
rect 7010 3984 7066 4040
rect 6734 3032 6790 3088
rect 6642 2352 6698 2408
rect 7102 3440 7158 3496
rect 7010 3168 7066 3224
rect 6366 992 6422 1048
rect 7010 2896 7066 2952
rect 7010 2624 7066 2680
rect 6918 856 6974 912
rect 6826 176 6882 232
rect 7838 10104 7894 10160
rect 7838 9424 7894 9480
rect 7838 8472 7894 8528
rect 7838 8200 7894 8256
rect 8114 11056 8170 11112
rect 8114 10512 8170 10568
rect 8574 20168 8630 20224
rect 8574 19896 8630 19952
rect 8574 19080 8630 19136
rect 8390 15680 8446 15736
rect 8390 12552 8446 12608
rect 8390 12416 8446 12472
rect 8390 12008 8446 12064
rect 8206 9696 8262 9752
rect 8022 8336 8078 8392
rect 8298 8744 8354 8800
rect 7562 4256 7618 4312
rect 7470 3712 7526 3768
rect 7838 5616 7894 5672
rect 7838 4936 7894 4992
rect 7746 4256 7802 4312
rect 7562 2760 7618 2816
rect 8574 12688 8630 12744
rect 8482 11328 8538 11384
rect 8574 10240 8630 10296
rect 8574 9832 8630 9888
rect 8850 21528 8906 21584
rect 9218 21528 9274 21584
rect 9678 22208 9734 22264
rect 9862 22208 9918 22264
rect 8758 21256 8814 21312
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 9034 20712 9090 20768
rect 9218 20712 9274 20768
rect 8758 19760 8814 19816
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8942 19624 8998 19680
rect 8850 19216 8906 19272
rect 9034 19216 9090 19272
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8758 17992 8814 18048
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 8758 17856 8814 17912
rect 9034 17584 9090 17640
rect 8758 17448 8814 17504
rect 9310 17584 9366 17640
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 8942 16360 8998 16416
rect 9126 16360 9182 16416
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8850 15408 8906 15464
rect 9310 15000 9366 15056
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 9310 13912 9366 13968
rect 9678 21256 9734 21312
rect 9632 21120 9688 21176
rect 9494 20848 9550 20904
rect 9494 18944 9550 19000
rect 9494 18264 9550 18320
rect 9586 17176 9642 17232
rect 9494 17040 9550 17096
rect 9770 16632 9826 16688
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 8758 12008 8814 12064
rect 8942 12824 8998 12880
rect 9126 12688 9182 12744
rect 9402 12688 9458 12744
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 9126 12280 9182 12336
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8758 10376 8814 10432
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8758 9288 8814 9344
rect 8758 9152 8814 9208
rect 9678 14728 9734 14784
rect 9678 14456 9734 14512
rect 9770 14320 9826 14376
rect 9678 14048 9734 14104
rect 9586 13368 9642 13424
rect 9586 11464 9642 11520
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 8850 8880 8906 8936
rect 8574 8744 8630 8800
rect 8482 8472 8538 8528
rect 8114 6568 8170 6624
rect 8482 8200 8538 8256
rect 8390 7520 8446 7576
rect 8574 7656 8630 7712
rect 8390 6704 8446 6760
rect 8298 5888 8354 5944
rect 8114 4800 8170 4856
rect 8022 4392 8078 4448
rect 8022 4256 8078 4312
rect 7930 4120 7986 4176
rect 8114 3848 8170 3904
rect 8758 8336 8814 8392
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 8574 5888 8630 5944
rect 8390 4528 8446 4584
rect 9126 7520 9182 7576
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 9402 7520 9458 7576
rect 9402 7112 9458 7168
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 9402 5888 9458 5944
rect 8206 3712 8262 3768
rect 8114 3576 8170 3632
rect 8298 3576 8354 3632
rect 8298 3304 8354 3360
rect 8114 448 8170 504
rect 7746 312 7802 368
rect 8666 4004 8722 4040
rect 8666 3984 8668 4004
rect 8668 3984 8720 4004
rect 8720 3984 8722 4004
rect 9034 5344 9090 5400
rect 8942 5072 8998 5128
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8850 4392 8906 4448
rect 8574 3304 8630 3360
rect 9218 4120 9274 4176
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 8666 2760 8722 2816
rect 8482 1400 8538 1456
rect 8850 2896 8906 2952
rect 9218 3032 9274 3088
rect 9034 2896 9090 2952
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 9770 12960 9826 13016
rect 9862 12144 9918 12200
rect 10046 12280 10102 12336
rect 9954 11872 10010 11928
rect 9954 10512 10010 10568
rect 10046 10412 10048 10432
rect 10048 10412 10100 10432
rect 10100 10412 10102 10432
rect 10046 10376 10102 10412
rect 9494 4528 9550 4584
rect 9770 9016 9826 9072
rect 9770 8336 9826 8392
rect 9678 6432 9734 6488
rect 9678 6024 9734 6080
rect 10506 21800 10562 21856
rect 10322 17856 10378 17912
rect 10874 21528 10930 21584
rect 10598 18400 10654 18456
rect 10690 17312 10746 17368
rect 10506 15000 10562 15056
rect 10690 13640 10746 13696
rect 11242 20168 11298 20224
rect 11058 19116 11060 19136
rect 11060 19116 11112 19136
rect 11112 19116 11114 19136
rect 11058 19080 11114 19116
rect 11150 18536 11206 18592
rect 11150 16768 11206 16824
rect 11058 14864 11114 14920
rect 10506 12144 10562 12200
rect 10782 12824 10838 12880
rect 9954 5480 10010 5536
rect 10138 5752 10194 5808
rect 10046 5344 10102 5400
rect 10322 5344 10378 5400
rect 9862 4936 9918 4992
rect 9678 4800 9734 4856
rect 9770 4256 9826 4312
rect 9586 3984 9642 4040
rect 9402 2896 9458 2952
rect 9862 4120 9918 4176
rect 9402 1944 9458 2000
rect 8758 720 8814 776
rect 9954 3576 10010 3632
rect 10138 4936 10194 4992
rect 10230 4528 10286 4584
rect 10138 4120 10194 4176
rect 10322 4120 10378 4176
rect 10138 3848 10194 3904
rect 10046 2624 10102 2680
rect 10322 3712 10378 3768
rect 10230 2896 10286 2952
rect 10690 10648 10746 10704
rect 10506 7248 10562 7304
rect 10690 8744 10746 8800
rect 10966 12552 11022 12608
rect 10874 11872 10930 11928
rect 10782 8064 10838 8120
rect 10782 7656 10838 7712
rect 10598 4800 10654 4856
rect 10598 4256 10654 4312
rect 11518 20440 11574 20496
rect 13542 23024 13598 23080
rect 13542 21936 13598 21992
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12806 21664 12862 21720
rect 11886 20848 11942 20904
rect 11978 20712 12034 20768
rect 11426 15680 11482 15736
rect 11426 15136 11482 15192
rect 11334 13912 11390 13968
rect 11150 12280 11206 12336
rect 11426 13096 11482 13152
rect 11242 11600 11298 11656
rect 11058 9424 11114 9480
rect 10966 7248 11022 7304
rect 11150 6432 11206 6488
rect 10966 3984 11022 4040
rect 10874 3848 10930 3904
rect 10874 3576 10930 3632
rect 10690 3032 10746 3088
rect 11426 11056 11482 11112
rect 11334 10648 11390 10704
rect 11334 10512 11390 10568
rect 11794 17176 11850 17232
rect 11702 12552 11758 12608
rect 11702 10104 11758 10160
rect 11610 8880 11666 8936
rect 11610 8744 11666 8800
rect 11334 8336 11390 8392
rect 11334 4392 11390 4448
rect 11978 16360 12034 16416
rect 12438 20168 12494 20224
rect 12530 19896 12586 19952
rect 12530 19488 12586 19544
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 12254 14184 12310 14240
rect 12070 11192 12126 11248
rect 11886 9424 11942 9480
rect 11886 8744 11942 8800
rect 11886 6840 11942 6896
rect 11150 2760 11206 2816
rect 11794 5480 11850 5536
rect 11610 3168 11666 3224
rect 11426 1264 11482 1320
rect 12346 12688 12402 12744
rect 12438 12552 12494 12608
rect 12438 12416 12494 12472
rect 12346 12008 12402 12064
rect 12254 9832 12310 9888
rect 12254 9424 12310 9480
rect 12162 9152 12218 9208
rect 12438 10784 12494 10840
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 13266 19216 13322 19272
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 13174 17856 13230 17912
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12806 17176 12862 17232
rect 12622 17040 12678 17096
rect 12806 16904 12862 16960
rect 13174 16904 13230 16960
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12622 15272 12678 15328
rect 12530 10648 12586 10704
rect 12162 7792 12218 7848
rect 12070 3984 12126 4040
rect 11886 2624 11942 2680
rect 12070 3440 12126 3496
rect 12990 15816 13046 15872
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 12806 15136 12862 15192
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 13358 16360 13414 16416
rect 14002 22888 14058 22944
rect 13542 18128 13598 18184
rect 13634 17856 13690 17912
rect 13818 19080 13874 19136
rect 13358 13912 13414 13968
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 13174 12552 13230 12608
rect 12990 12416 13046 12472
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 12806 11600 12862 11656
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 12990 10648 13046 10704
rect 12622 9968 12678 10024
rect 11702 584 11758 640
rect 12898 10104 12954 10160
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 13358 11056 13414 11112
rect 13450 10920 13506 10976
rect 13450 10784 13506 10840
rect 13358 10240 13414 10296
rect 13358 10104 13414 10160
rect 14094 18808 14150 18864
rect 14002 18264 14058 18320
rect 14002 17856 14058 17912
rect 13818 16088 13874 16144
rect 13726 12824 13782 12880
rect 14094 17720 14150 17776
rect 14002 15952 14058 16008
rect 13910 11736 13966 11792
rect 13910 11056 13966 11112
rect 14186 13912 14242 13968
rect 14186 11600 14242 11656
rect 14002 10648 14058 10704
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 13082 8336 13138 8392
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 12898 7384 12954 7440
rect 12806 6704 12862 6760
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 12806 5072 12862 5128
rect 12806 4936 12862 4992
rect 13358 8200 13414 8256
rect 13542 9696 13598 9752
rect 14002 10240 14058 10296
rect 13818 9288 13874 9344
rect 13726 8472 13782 8528
rect 14094 9016 14150 9072
rect 14002 8880 14058 8936
rect 14094 8744 14150 8800
rect 14094 8064 14150 8120
rect 13910 6840 13966 6896
rect 12898 4528 12954 4584
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 12622 3304 12678 3360
rect 13174 3576 13230 3632
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 12714 3032 12770 3088
rect 12622 2488 12678 2544
rect 12714 2216 12770 2272
rect 12530 1808 12586 1864
rect 12898 2488 12954 2544
rect 13542 5344 13598 5400
rect 13726 4664 13782 4720
rect 13726 3576 13782 3632
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 12806 1672 12862 1728
rect 14462 22072 14518 22128
rect 14370 12960 14426 13016
rect 14370 9968 14426 10024
rect 14646 17040 14702 17096
rect 14554 15680 14610 15736
rect 15014 21256 15070 21312
rect 15014 19216 15070 19272
rect 15014 18264 15070 18320
rect 15014 17856 15070 17912
rect 15198 20168 15254 20224
rect 15198 20032 15254 20088
rect 15106 17720 15162 17776
rect 14922 17584 14978 17640
rect 14922 17448 14978 17504
rect 14738 15272 14794 15328
rect 14554 13912 14610 13968
rect 14554 13504 14610 13560
rect 14646 13368 14702 13424
rect 14646 10784 14702 10840
rect 14186 7656 14242 7712
rect 15106 14728 15162 14784
rect 15198 14320 15254 14376
rect 15934 20984 15990 21040
rect 14922 12416 14978 12472
rect 15014 11600 15070 11656
rect 15014 10104 15070 10160
rect 14738 9968 14794 10024
rect 14462 8200 14518 8256
rect 14370 6432 14426 6488
rect 14094 4256 14150 4312
rect 15014 9424 15070 9480
rect 14738 7520 14794 7576
rect 14370 5344 14426 5400
rect 14554 5344 14610 5400
rect 14370 4528 14426 4584
rect 14462 2488 14518 2544
rect 14738 1808 14794 1864
rect 14094 176 14150 232
rect 15014 7384 15070 7440
rect 15014 7248 15070 7304
rect 15290 10920 15346 10976
rect 15290 10376 15346 10432
rect 15566 12416 15622 12472
rect 15566 10648 15622 10704
rect 16026 18672 16082 18728
rect 16026 17176 16082 17232
rect 15566 7792 15622 7848
rect 15566 7248 15622 7304
rect 15290 4120 15346 4176
rect 15014 3032 15070 3088
rect 15474 5072 15530 5128
rect 15934 14184 15990 14240
rect 15934 14048 15990 14104
rect 16026 13640 16082 13696
rect 16026 12552 16082 12608
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16762 21120 16818 21176
rect 16946 20848 17002 20904
rect 15750 7112 15806 7168
rect 15842 6160 15898 6216
rect 15658 5208 15714 5264
rect 15750 3848 15806 3904
rect 15658 3712 15714 3768
rect 16118 5072 16174 5128
rect 16118 4664 16174 4720
rect 16762 19896 16818 19952
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16762 17992 16818 18048
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16946 15408 17002 15464
rect 17038 15136 17094 15192
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 17590 22752 17646 22808
rect 16762 14048 16818 14104
rect 16670 13504 16726 13560
rect 17866 22480 17922 22536
rect 17866 18028 17868 18048
rect 17868 18028 17920 18048
rect 17920 18028 17922 18048
rect 17866 17992 17922 18028
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16762 11328 16818 11384
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 17222 11736 17278 11792
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16946 10512 17002 10568
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 17130 10104 17186 10160
rect 16946 9968 17002 10024
rect 16670 9016 16726 9072
rect 16670 8880 16726 8936
rect 16578 6160 16634 6216
rect 16302 5480 16358 5536
rect 16486 5888 16542 5944
rect 16394 5208 16450 5264
rect 15934 4392 15990 4448
rect 15842 3712 15898 3768
rect 16210 3712 16266 3768
rect 15750 3440 15806 3496
rect 16026 3440 16082 3496
rect 15658 3304 15714 3360
rect 15658 3168 15714 3224
rect 14922 40 14978 96
rect 16118 3032 16174 3088
rect 16026 2760 16082 2816
rect 17498 11600 17554 11656
rect 17406 10240 17462 10296
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 17222 9016 17278 9072
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16854 6296 16910 6352
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 18142 20304 18198 20360
rect 18050 13776 18106 13832
rect 18510 15000 18566 15056
rect 18786 15272 18842 15328
rect 18602 13504 18658 13560
rect 18418 13232 18474 13288
rect 18602 12960 18658 13016
rect 18878 13912 18934 13968
rect 18418 9968 18474 10024
rect 18326 9696 18382 9752
rect 18050 9152 18106 9208
rect 17590 6296 17646 6352
rect 16762 4800 16818 4856
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16394 856 16450 912
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 17682 5888 17738 5944
rect 17498 4936 17554 4992
rect 17866 5616 17922 5672
rect 17866 5344 17922 5400
rect 17406 3848 17462 3904
rect 17498 2896 17554 2952
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 17406 2624 17462 2680
rect 17866 4528 17922 4584
rect 18142 6840 18198 6896
rect 18326 7520 18382 7576
rect 18326 5752 18382 5808
rect 18418 5208 18474 5264
rect 18510 4256 18566 4312
rect 18142 3848 18198 3904
rect 17222 2488 17278 2544
rect 18694 5480 18750 5536
rect 19062 15680 19118 15736
rect 21730 22888 21786 22944
rect 20258 21936 20314 21992
rect 19798 21392 19854 21448
rect 19430 20440 19486 20496
rect 19706 20168 19762 20224
rect 19338 15816 19394 15872
rect 19338 15680 19394 15736
rect 19246 14320 19302 14376
rect 18970 6024 19026 6080
rect 19798 18400 19854 18456
rect 19614 11464 19670 11520
rect 19430 8744 19486 8800
rect 19246 7248 19302 7304
rect 19246 5344 19302 5400
rect 19154 4800 19210 4856
rect 18878 4392 18934 4448
rect 18786 4256 18842 4312
rect 18970 4256 19026 4312
rect 18970 4120 19026 4176
rect 18878 3984 18934 4040
rect 19062 3984 19118 4040
rect 19614 4664 19670 4720
rect 18694 3304 18750 3360
rect 18050 1400 18106 1456
rect 18878 2624 18934 2680
rect 19522 3984 19578 4040
rect 20074 19352 20130 19408
rect 19890 15136 19946 15192
rect 21454 21800 21510 21856
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 20810 21664 20866 21720
rect 20626 21528 20682 21584
rect 20258 16360 20314 16416
rect 20166 14864 20222 14920
rect 19982 13096 20038 13152
rect 19890 12280 19946 12336
rect 19890 10784 19946 10840
rect 19982 9968 20038 10024
rect 19798 7384 19854 7440
rect 20166 9152 20222 9208
rect 20074 4664 20130 4720
rect 20442 18128 20498 18184
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20718 18264 20774 18320
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 21638 20712 21694 20768
rect 21546 18536 21602 18592
rect 21362 17448 21418 17504
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 20718 15544 20774 15600
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 20534 14456 20590 14512
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20902 13232 20958 13288
rect 20810 13096 20866 13152
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20442 10376 20498 10432
rect 21270 12280 21326 12336
rect 21822 19760 21878 19816
rect 21914 19216 21970 19272
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20626 9832 20682 9888
rect 20442 8200 20498 8256
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21086 9424 21142 9480
rect 21362 12008 21418 12064
rect 21270 8880 21326 8936
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20718 7928 20774 7984
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20626 6704 20682 6760
rect 19890 4392 19946 4448
rect 19982 4120 20038 4176
rect 19890 3440 19946 3496
rect 19614 3032 19670 3088
rect 20074 3032 20130 3088
rect 19338 1128 19394 1184
rect 19706 448 19762 504
rect 19890 2216 19946 2272
rect 20718 6432 20774 6488
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20534 5072 20590 5128
rect 20350 4528 20406 4584
rect 20258 720 20314 776
rect 20994 4936 21050 4992
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 21454 9968 21510 10024
rect 21638 12144 21694 12200
rect 21730 9016 21786 9072
rect 21638 7792 21694 7848
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 21730 4120 21786 4176
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 20718 1264 20774 1320
rect 20350 584 20406 640
rect 22006 11328 22062 11384
rect 22006 10920 22062 10976
rect 21914 10512 21970 10568
rect 22006 9288 22062 9344
rect 22006 8472 22062 8528
rect 22742 14184 22798 14240
rect 22282 12688 22338 12744
rect 22282 11192 22338 11248
rect 22374 10240 22430 10296
rect 22282 9832 22338 9888
rect 22190 6568 22246 6624
rect 22282 5072 22338 5128
rect 22006 3576 22062 3632
rect 22098 2760 22154 2816
rect 21730 2352 21786 2408
rect 22466 4664 22522 4720
rect 21730 1944 21786 2000
rect 22282 312 22338 368
rect 21454 40 21510 96
rect 23570 16904 23626 16960
rect 23570 13640 23626 13696
rect 22742 11736 22798 11792
rect 22650 5480 22706 5536
rect 23570 7112 23626 7168
rect 23570 3848 23626 3904
<< metal3 >>
rect 0 23400 480 23520
rect 23520 23400 24000 23520
rect 62 22946 122 23400
rect 841 23218 907 23221
rect 841 23216 3940 23218
rect 841 23160 846 23216
rect 902 23160 3940 23216
rect 841 23158 3940 23160
rect 841 23155 907 23158
rect 3550 23020 3556 23084
rect 3620 23082 3626 23084
rect 3693 23082 3759 23085
rect 3620 23080 3759 23082
rect 3620 23024 3698 23080
rect 3754 23024 3759 23080
rect 3620 23022 3759 23024
rect 3880 23082 3940 23158
rect 13537 23082 13603 23085
rect 3880 23080 13603 23082
rect 3880 23024 13542 23080
rect 13598 23024 13603 23080
rect 3880 23022 13603 23024
rect 3620 23020 3626 23022
rect 3693 23019 3759 23022
rect 13537 23019 13603 23022
rect 1393 22946 1459 22949
rect 62 22944 1459 22946
rect 62 22888 1398 22944
rect 1454 22888 1459 22944
rect 62 22886 1459 22888
rect 1393 22883 1459 22886
rect 2814 22884 2820 22948
rect 2884 22946 2890 22948
rect 7649 22946 7715 22949
rect 2884 22944 7715 22946
rect 2884 22888 7654 22944
rect 7710 22888 7715 22944
rect 2884 22886 7715 22888
rect 2884 22884 2890 22886
rect 7649 22883 7715 22886
rect 7833 22946 7899 22949
rect 13997 22946 14063 22949
rect 7833 22944 14063 22946
rect 7833 22888 7838 22944
rect 7894 22888 14002 22944
rect 14058 22888 14063 22944
rect 7833 22886 14063 22888
rect 7833 22883 7899 22886
rect 13997 22883 14063 22886
rect 21725 22946 21791 22949
rect 23614 22946 23674 23400
rect 21725 22944 23674 22946
rect 21725 22888 21730 22944
rect 21786 22888 23674 22944
rect 21725 22886 23674 22888
rect 21725 22883 21791 22886
rect 1669 22810 1735 22813
rect 6637 22810 6703 22813
rect 1669 22808 6703 22810
rect 1669 22752 1674 22808
rect 1730 22752 6642 22808
rect 6698 22752 6703 22808
rect 1669 22750 6703 22752
rect 1669 22747 1735 22750
rect 6637 22747 6703 22750
rect 7966 22748 7972 22812
rect 8036 22810 8042 22812
rect 17585 22810 17651 22813
rect 8036 22808 17651 22810
rect 8036 22752 17590 22808
rect 17646 22752 17651 22808
rect 8036 22750 17651 22752
rect 8036 22748 8042 22750
rect 17585 22747 17651 22750
rect 0 22584 480 22704
rect 749 22674 815 22677
rect 7373 22674 7439 22677
rect 749 22672 7439 22674
rect 749 22616 754 22672
rect 810 22616 7378 22672
rect 7434 22616 7439 22672
rect 749 22614 7439 22616
rect 749 22611 815 22614
rect 7373 22611 7439 22614
rect 7557 22674 7623 22677
rect 17902 22674 17908 22676
rect 7557 22672 17908 22674
rect 7557 22616 7562 22672
rect 7618 22616 17908 22672
rect 7557 22614 17908 22616
rect 7557 22611 7623 22614
rect 17902 22612 17908 22614
rect 17972 22612 17978 22676
rect 62 22130 122 22584
rect 3918 22476 3924 22540
rect 3988 22538 3994 22540
rect 8201 22538 8267 22541
rect 3988 22536 8267 22538
rect 3988 22480 8206 22536
rect 8262 22480 8267 22536
rect 3988 22478 8267 22480
rect 3988 22476 3994 22478
rect 8201 22475 8267 22478
rect 8661 22538 8727 22541
rect 17861 22538 17927 22541
rect 8661 22536 17927 22538
rect 8661 22480 8666 22536
rect 8722 22480 17866 22536
rect 17922 22480 17927 22536
rect 8661 22478 17927 22480
rect 8661 22475 8727 22478
rect 17861 22475 17927 22478
rect 1301 22402 1367 22405
rect 15694 22402 15700 22404
rect 1301 22400 15700 22402
rect 1301 22344 1306 22400
rect 1362 22344 15700 22400
rect 1301 22342 15700 22344
rect 1301 22339 1367 22342
rect 15694 22340 15700 22342
rect 15764 22340 15770 22404
rect 23520 22312 24000 22432
rect 1894 22204 1900 22268
rect 1964 22266 1970 22268
rect 9673 22266 9739 22269
rect 1964 22264 9739 22266
rect 1964 22208 9678 22264
rect 9734 22208 9739 22264
rect 1964 22206 9739 22208
rect 1964 22204 1970 22206
rect 9673 22203 9739 22206
rect 9857 22266 9923 22269
rect 12382 22266 12388 22268
rect 9857 22264 12388 22266
rect 9857 22208 9862 22264
rect 9918 22208 12388 22264
rect 9857 22206 12388 22208
rect 9857 22203 9923 22206
rect 12382 22204 12388 22206
rect 12452 22204 12458 22268
rect 62 22070 4170 22130
rect 4110 21994 4170 22070
rect 4654 22068 4660 22132
rect 4724 22130 4730 22132
rect 4889 22130 4955 22133
rect 8293 22130 8359 22133
rect 14457 22130 14523 22133
rect 4724 22128 14523 22130
rect 4724 22072 4894 22128
rect 4950 22072 8298 22128
rect 8354 22072 14462 22128
rect 14518 22072 14523 22128
rect 4724 22070 14523 22072
rect 4724 22068 4730 22070
rect 4889 22067 4955 22070
rect 8293 22067 8359 22070
rect 14457 22067 14523 22070
rect 7373 21994 7439 21997
rect 13537 21994 13603 21997
rect 20253 21994 20319 21997
rect 4110 21934 5642 21994
rect 0 21768 480 21888
rect 5582 21858 5642 21934
rect 7373 21992 13416 21994
rect 7373 21936 7378 21992
rect 7434 21936 13416 21992
rect 7373 21934 13416 21936
rect 7373 21931 7439 21934
rect 10501 21858 10567 21861
rect 5582 21856 10567 21858
rect 5582 21800 10506 21856
rect 10562 21800 10567 21856
rect 5582 21798 10567 21800
rect 10501 21795 10567 21798
rect 4944 21792 5264 21793
rect 62 21314 122 21768
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 7005 21722 7071 21725
rect 12801 21722 12867 21725
rect 7005 21720 12867 21722
rect 7005 21664 7010 21720
rect 7066 21664 12806 21720
rect 12862 21664 12867 21720
rect 7005 21662 12867 21664
rect 13356 21722 13416 21934
rect 13537 21992 20319 21994
rect 13537 21936 13542 21992
rect 13598 21936 20258 21992
rect 20314 21936 20319 21992
rect 13537 21934 20319 21936
rect 13537 21931 13603 21934
rect 20253 21931 20319 21934
rect 21449 21858 21515 21861
rect 23614 21858 23674 22312
rect 21449 21856 23674 21858
rect 21449 21800 21454 21856
rect 21510 21800 23674 21856
rect 21449 21798 23674 21800
rect 21449 21795 21515 21798
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 20805 21722 20871 21725
rect 13356 21720 20871 21722
rect 13356 21664 20810 21720
rect 20866 21664 20871 21720
rect 13356 21662 20871 21664
rect 7005 21659 7071 21662
rect 12801 21659 12867 21662
rect 20805 21659 20871 21662
rect 381 21586 447 21589
rect 8845 21586 8911 21589
rect 381 21584 8911 21586
rect 381 21528 386 21584
rect 442 21528 8850 21584
rect 8906 21528 8911 21584
rect 381 21526 8911 21528
rect 381 21523 447 21526
rect 8845 21523 8911 21526
rect 9213 21586 9279 21589
rect 10542 21586 10548 21588
rect 9213 21584 10548 21586
rect 9213 21528 9218 21584
rect 9274 21528 10548 21584
rect 9213 21526 10548 21528
rect 9213 21523 9279 21526
rect 10542 21524 10548 21526
rect 10612 21524 10618 21588
rect 10869 21586 10935 21589
rect 20621 21586 20687 21589
rect 10869 21584 20687 21586
rect 10869 21528 10874 21584
rect 10930 21528 20626 21584
rect 20682 21528 20687 21584
rect 10869 21526 20687 21528
rect 10869 21523 10935 21526
rect 20621 21523 20687 21526
rect 3049 21450 3115 21453
rect 19793 21450 19859 21453
rect 3049 21448 19859 21450
rect 3049 21392 3054 21448
rect 3110 21392 19798 21448
rect 19854 21392 19859 21448
rect 3049 21390 19859 21392
rect 3049 21387 3115 21390
rect 19793 21387 19859 21390
rect 1577 21314 1643 21317
rect 62 21312 1643 21314
rect 62 21256 1582 21312
rect 1638 21256 1643 21312
rect 62 21254 1643 21256
rect 1577 21251 1643 21254
rect 2313 21314 2379 21317
rect 8753 21314 8819 21317
rect 2313 21312 8819 21314
rect 2313 21256 2318 21312
rect 2374 21256 8758 21312
rect 8814 21256 8819 21312
rect 2313 21254 8819 21256
rect 2313 21251 2379 21254
rect 8753 21251 8819 21254
rect 9673 21314 9739 21317
rect 15009 21314 15075 21317
rect 9673 21312 15075 21314
rect 9673 21256 9678 21312
rect 9734 21256 15014 21312
rect 15070 21256 15075 21312
rect 9673 21254 15075 21256
rect 9673 21251 9739 21254
rect 15009 21251 15075 21254
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 23520 21224 24000 21344
rect 16944 21183 17264 21184
rect 2221 21178 2287 21181
rect 7649 21178 7715 21181
rect 2221 21176 7715 21178
rect 2221 21120 2226 21176
rect 2282 21120 7654 21176
rect 7710 21120 7715 21176
rect 2221 21118 7715 21120
rect 2221 21115 2287 21118
rect 7649 21115 7715 21118
rect 9627 21178 9693 21181
rect 16757 21178 16823 21181
rect 9627 21176 16823 21178
rect 9627 21120 9632 21176
rect 9688 21120 16762 21176
rect 16818 21120 16823 21176
rect 9627 21118 16823 21120
rect 9627 21115 9693 21118
rect 16757 21115 16823 21118
rect 0 20952 480 21072
rect 3182 20980 3188 21044
rect 3252 21042 3258 21044
rect 4102 21042 4108 21044
rect 3252 20982 4108 21042
rect 3252 20980 3258 20982
rect 4102 20980 4108 20982
rect 4172 20980 4178 21044
rect 4429 21042 4495 21045
rect 4429 21040 9322 21042
rect 4429 20984 4434 21040
rect 4490 20984 9322 21040
rect 4429 20982 9322 20984
rect 4429 20979 4495 20982
rect 62 20498 122 20952
rect 9262 20940 9322 20982
rect 9806 20980 9812 21044
rect 9876 21042 9882 21044
rect 15929 21042 15995 21045
rect 9876 21040 15995 21042
rect 9876 20984 15934 21040
rect 15990 20984 15995 21040
rect 9876 20982 15995 20984
rect 9876 20980 9882 20982
rect 15929 20979 15995 20982
rect 9622 20940 9628 20942
rect 5441 20906 5507 20909
rect 9262 20906 9628 20940
rect 2408 20904 9628 20906
rect 2408 20848 5446 20904
rect 5502 20848 9494 20904
rect 9550 20880 9628 20904
rect 9550 20848 9555 20880
rect 9622 20878 9628 20880
rect 9692 20878 9698 20942
rect 11881 20906 11947 20909
rect 16941 20906 17007 20909
rect 11881 20904 17007 20906
rect 2408 20846 9555 20848
rect 238 20708 244 20772
rect 308 20770 314 20772
rect 2408 20770 2468 20846
rect 5441 20843 5507 20846
rect 9489 20843 9555 20846
rect 11881 20848 11886 20904
rect 11942 20848 16946 20904
rect 17002 20848 17007 20904
rect 11881 20846 17007 20848
rect 11881 20843 11947 20846
rect 16941 20843 17007 20846
rect 308 20710 2468 20770
rect 2773 20770 2839 20773
rect 4705 20770 4771 20773
rect 2773 20768 4771 20770
rect 2773 20712 2778 20768
rect 2834 20712 4710 20768
rect 4766 20712 4771 20768
rect 2773 20710 4771 20712
rect 308 20708 314 20710
rect 2773 20707 2839 20710
rect 4705 20707 4771 20710
rect 5349 20770 5415 20773
rect 8385 20770 8451 20773
rect 9029 20770 9095 20773
rect 5349 20768 9095 20770
rect 5349 20712 5354 20768
rect 5410 20712 8390 20768
rect 8446 20712 9034 20768
rect 9090 20712 9095 20768
rect 5349 20710 9095 20712
rect 5349 20707 5415 20710
rect 8385 20707 8451 20710
rect 9029 20707 9095 20710
rect 9213 20770 9279 20773
rect 10174 20770 10180 20772
rect 9213 20768 10180 20770
rect 9213 20712 9218 20768
rect 9274 20712 10180 20768
rect 9213 20710 10180 20712
rect 9213 20707 9279 20710
rect 10174 20708 10180 20710
rect 10244 20708 10250 20772
rect 11973 20770 12039 20773
rect 12750 20770 12756 20772
rect 11973 20768 12756 20770
rect 11973 20712 11978 20768
rect 12034 20712 12756 20768
rect 11973 20710 12756 20712
rect 11973 20707 12039 20710
rect 12750 20708 12756 20710
rect 12820 20708 12826 20772
rect 21633 20770 21699 20773
rect 23614 20770 23674 21224
rect 21633 20768 23674 20770
rect 21633 20712 21638 20768
rect 21694 20712 23674 20768
rect 21633 20710 23674 20712
rect 21633 20707 21699 20710
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 197 20634 263 20637
rect 3601 20634 3667 20637
rect 197 20632 3667 20634
rect 197 20576 202 20632
rect 258 20576 3606 20632
rect 3662 20576 3667 20632
rect 197 20574 3667 20576
rect 197 20571 263 20574
rect 3601 20571 3667 20574
rect 7373 20634 7439 20637
rect 7373 20632 11714 20634
rect 7373 20576 7378 20632
rect 7434 20576 11714 20632
rect 7373 20574 11714 20576
rect 7373 20571 7439 20574
rect 62 20438 3296 20498
rect 3236 20362 3296 20438
rect 3366 20436 3372 20500
rect 3436 20498 3442 20500
rect 11513 20498 11579 20501
rect 3436 20496 11579 20498
rect 3436 20440 11518 20496
rect 11574 20440 11579 20496
rect 3436 20438 11579 20440
rect 11654 20498 11714 20574
rect 19425 20498 19491 20501
rect 11654 20496 19491 20498
rect 11654 20440 19430 20496
rect 19486 20440 19491 20496
rect 11654 20438 19491 20440
rect 3436 20436 3442 20438
rect 11513 20435 11579 20438
rect 19425 20435 19491 20438
rect 7005 20362 7071 20365
rect 3236 20360 7071 20362
rect 3236 20304 7010 20360
rect 7066 20304 7071 20360
rect 3236 20302 7071 20304
rect 7005 20299 7071 20302
rect 8702 20300 8708 20364
rect 8772 20362 8778 20364
rect 18137 20362 18203 20365
rect 8772 20360 18203 20362
rect 8772 20304 18142 20360
rect 18198 20304 18203 20360
rect 8772 20302 18203 20304
rect 8772 20300 8778 20302
rect 18137 20299 18203 20302
rect 0 20224 480 20256
rect 0 20168 18 20224
rect 74 20168 480 20224
rect 0 20136 480 20168
rect 2129 20226 2195 20229
rect 6545 20226 6611 20229
rect 2129 20224 6611 20226
rect 2129 20168 2134 20224
rect 2190 20168 6550 20224
rect 6606 20168 6611 20224
rect 2129 20166 6611 20168
rect 2129 20163 2195 20166
rect 6545 20163 6611 20166
rect 7046 20164 7052 20228
rect 7116 20226 7122 20228
rect 8569 20226 8635 20229
rect 7116 20224 8635 20226
rect 7116 20168 8574 20224
rect 8630 20168 8635 20224
rect 7116 20166 8635 20168
rect 7116 20164 7122 20166
rect 8569 20163 8635 20166
rect 11237 20226 11303 20229
rect 12433 20226 12499 20229
rect 15193 20226 15259 20229
rect 11237 20224 15259 20226
rect 11237 20168 11242 20224
rect 11298 20168 12438 20224
rect 12494 20168 15198 20224
rect 15254 20168 15259 20224
rect 11237 20166 15259 20168
rect 11237 20163 11303 20166
rect 12433 20163 12499 20166
rect 15193 20163 15259 20166
rect 19558 20164 19564 20228
rect 19628 20226 19634 20228
rect 19701 20226 19767 20229
rect 23520 20228 24000 20256
rect 23520 20226 23612 20228
rect 19628 20224 19767 20226
rect 19628 20168 19706 20224
rect 19762 20168 19767 20224
rect 19628 20166 19767 20168
rect 23484 20166 23612 20226
rect 19628 20164 19634 20166
rect 19701 20163 19767 20166
rect 23520 20164 23612 20166
rect 23676 20164 24000 20228
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 23520 20136 24000 20164
rect 16944 20095 17264 20096
rect 2129 20090 2195 20093
rect 3969 20090 4035 20093
rect 2129 20088 4035 20090
rect 2129 20032 2134 20088
rect 2190 20032 3974 20088
rect 4030 20032 4035 20088
rect 2129 20030 4035 20032
rect 2129 20027 2195 20030
rect 3969 20027 4035 20030
rect 4705 20090 4771 20093
rect 7833 20090 7899 20093
rect 4705 20088 7899 20090
rect 4705 20032 4710 20088
rect 4766 20032 7838 20088
rect 7894 20032 7899 20088
rect 4705 20030 7899 20032
rect 4705 20027 4771 20030
rect 7833 20027 7899 20030
rect 9438 20028 9444 20092
rect 9508 20090 9514 20092
rect 15193 20090 15259 20093
rect 9508 20088 15259 20090
rect 9508 20032 15198 20088
rect 15254 20032 15259 20088
rect 9508 20030 15259 20032
rect 9508 20028 9514 20030
rect 15193 20027 15259 20030
rect 473 19954 539 19957
rect 8569 19954 8635 19957
rect 473 19952 8635 19954
rect 473 19896 478 19952
rect 534 19896 8574 19952
rect 8630 19896 8635 19952
rect 473 19894 8635 19896
rect 473 19891 539 19894
rect 8569 19891 8635 19894
rect 12525 19954 12591 19957
rect 16757 19954 16823 19957
rect 12525 19952 16823 19954
rect 12525 19896 12530 19952
rect 12586 19896 16762 19952
rect 16818 19896 16823 19952
rect 12525 19894 16823 19896
rect 12525 19891 12591 19894
rect 16757 19891 16823 19894
rect 238 19756 244 19820
rect 308 19818 314 19820
rect 2221 19818 2287 19821
rect 308 19816 2287 19818
rect 308 19760 2226 19816
rect 2282 19760 2287 19816
rect 308 19758 2287 19760
rect 308 19756 314 19758
rect 2221 19755 2287 19758
rect 2957 19818 3023 19821
rect 7414 19818 7420 19820
rect 2957 19816 7420 19818
rect 2957 19760 2962 19816
rect 3018 19760 7420 19816
rect 2957 19758 7420 19760
rect 2957 19755 3023 19758
rect 7414 19756 7420 19758
rect 7484 19756 7490 19820
rect 8753 19818 8819 19821
rect 21817 19818 21883 19821
rect 8753 19816 21883 19818
rect 8753 19760 8758 19816
rect 8814 19760 21822 19816
rect 21878 19760 21883 19816
rect 8753 19758 21883 19760
rect 8753 19755 8819 19758
rect 21817 19755 21883 19758
rect 2497 19682 2563 19685
rect 2497 19680 4170 19682
rect 2497 19624 2502 19680
rect 2558 19624 4170 19680
rect 2497 19622 4170 19624
rect 2497 19619 2563 19622
rect 2078 19484 2084 19548
rect 2148 19546 2154 19548
rect 3233 19546 3299 19549
rect 2148 19544 3299 19546
rect 2148 19488 3238 19544
rect 3294 19488 3299 19544
rect 2148 19486 3299 19488
rect 2148 19484 2154 19486
rect 3233 19483 3299 19486
rect 0 19350 480 19440
rect 0 19320 674 19350
rect 62 19290 674 19320
rect 614 19274 674 19290
rect 3550 19274 3556 19276
rect 614 19214 3556 19274
rect 3550 19212 3556 19214
rect 3620 19212 3626 19276
rect 4110 19274 4170 19622
rect 5758 19620 5764 19684
rect 5828 19682 5834 19684
rect 6821 19682 6887 19685
rect 5828 19680 6887 19682
rect 5828 19624 6826 19680
rect 6882 19624 6887 19680
rect 5828 19622 6887 19624
rect 5828 19620 5834 19622
rect 6821 19619 6887 19622
rect 8150 19620 8156 19684
rect 8220 19682 8226 19684
rect 8937 19682 9003 19685
rect 8220 19680 9003 19682
rect 8220 19624 8942 19680
rect 8998 19624 9003 19680
rect 8220 19622 9003 19624
rect 8220 19620 8226 19622
rect 8937 19619 9003 19622
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 5390 19484 5396 19548
rect 5460 19546 5466 19548
rect 12525 19546 12591 19549
rect 17350 19546 17356 19548
rect 5460 19544 12591 19546
rect 5460 19488 12530 19544
rect 12586 19488 12591 19544
rect 5460 19486 12591 19488
rect 5460 19484 5466 19486
rect 12525 19483 12591 19486
rect 13356 19486 17356 19546
rect 4521 19410 4587 19413
rect 4797 19410 4863 19413
rect 4521 19408 4863 19410
rect 4521 19352 4526 19408
rect 4582 19352 4802 19408
rect 4858 19352 4863 19408
rect 4521 19350 4863 19352
rect 4521 19347 4587 19350
rect 4797 19347 4863 19350
rect 6862 19348 6868 19412
rect 6932 19410 6938 19412
rect 13356 19410 13416 19486
rect 17350 19484 17356 19486
rect 17420 19484 17426 19548
rect 6932 19350 13416 19410
rect 6932 19348 6938 19350
rect 13670 19348 13676 19412
rect 13740 19410 13746 19412
rect 20069 19410 20135 19413
rect 13740 19408 20135 19410
rect 13740 19352 20074 19408
rect 20130 19352 20135 19408
rect 13740 19350 20135 19352
rect 13740 19348 13746 19350
rect 20069 19347 20135 19350
rect 5349 19274 5415 19277
rect 8845 19274 8911 19277
rect 4110 19272 8911 19274
rect 4110 19216 5354 19272
rect 5410 19216 8850 19272
rect 8906 19216 8911 19272
rect 4110 19214 8911 19216
rect 5349 19211 5415 19214
rect 8845 19211 8911 19214
rect 9029 19274 9095 19277
rect 13261 19274 13327 19277
rect 9029 19272 13327 19274
rect 9029 19216 9034 19272
rect 9090 19216 13266 19272
rect 13322 19216 13327 19272
rect 9029 19214 13327 19216
rect 9029 19211 9095 19214
rect 13261 19211 13327 19214
rect 15009 19274 15075 19277
rect 21909 19274 21975 19277
rect 15009 19272 21975 19274
rect 15009 19216 15014 19272
rect 15070 19216 21914 19272
rect 21970 19216 21975 19272
rect 15009 19214 21975 19216
rect 15009 19211 15075 19214
rect 21909 19211 21975 19214
rect 1158 19076 1164 19140
rect 1228 19138 1234 19140
rect 2037 19138 2103 19141
rect 1228 19136 2103 19138
rect 1228 19080 2042 19136
rect 2098 19080 2103 19136
rect 1228 19078 2103 19080
rect 1228 19076 1234 19078
rect 2037 19075 2103 19078
rect 3141 19138 3207 19141
rect 6269 19138 6335 19141
rect 8569 19138 8635 19141
rect 3141 19136 8635 19138
rect 3141 19080 3146 19136
rect 3202 19080 6274 19136
rect 6330 19080 8574 19136
rect 8630 19080 8635 19136
rect 3141 19078 8635 19080
rect 3141 19075 3207 19078
rect 6269 19075 6335 19078
rect 8569 19075 8635 19078
rect 11053 19138 11119 19141
rect 13813 19138 13879 19141
rect 11053 19136 13879 19138
rect 11053 19080 11058 19136
rect 11114 19080 13818 19136
rect 13874 19080 13879 19136
rect 11053 19078 13879 19080
rect 11053 19075 11119 19078
rect 13813 19075 13879 19078
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 23520 19048 24000 19168
rect 16944 19007 17264 19008
rect 3877 19002 3943 19005
rect 4797 19002 4863 19005
rect 7598 19002 7604 19004
rect 3877 19000 7604 19002
rect 3877 18944 3882 19000
rect 3938 18944 4802 19000
rect 4858 18944 7604 19000
rect 3877 18942 7604 18944
rect 3877 18939 3943 18942
rect 4797 18939 4863 18942
rect 7598 18940 7604 18942
rect 7668 18940 7674 19004
rect 9489 19002 9555 19005
rect 14038 19002 14044 19004
rect 9489 19000 14044 19002
rect 9489 18944 9494 19000
rect 9550 18944 14044 19000
rect 9489 18942 14044 18944
rect 9489 18939 9555 18942
rect 14038 18940 14044 18942
rect 14108 18940 14114 19004
rect 4102 18804 4108 18868
rect 4172 18866 4178 18868
rect 5809 18866 5875 18869
rect 14089 18866 14155 18869
rect 4172 18806 5412 18866
rect 4172 18804 4178 18806
rect 0 18504 480 18624
rect 1526 18532 1532 18596
rect 1596 18594 1602 18596
rect 4337 18594 4403 18597
rect 1596 18592 4403 18594
rect 1596 18536 4342 18592
rect 4398 18536 4403 18592
rect 1596 18534 4403 18536
rect 5352 18594 5412 18806
rect 5809 18864 14155 18866
rect 5809 18808 5814 18864
rect 5870 18808 14094 18864
rect 14150 18808 14155 18864
rect 5809 18806 14155 18808
rect 5809 18803 5875 18806
rect 14089 18803 14155 18806
rect 6494 18668 6500 18732
rect 6564 18730 6570 18732
rect 14590 18730 14596 18732
rect 6564 18670 14596 18730
rect 6564 18668 6570 18670
rect 14590 18668 14596 18670
rect 14660 18730 14666 18732
rect 16021 18730 16087 18733
rect 14660 18728 16087 18730
rect 14660 18672 16026 18728
rect 16082 18672 16087 18728
rect 14660 18670 16087 18672
rect 14660 18668 14666 18670
rect 16021 18667 16087 18670
rect 10174 18594 10180 18596
rect 5352 18534 10180 18594
rect 1596 18532 1602 18534
rect 4337 18531 4403 18534
rect 10174 18532 10180 18534
rect 10244 18532 10250 18596
rect 11145 18594 11211 18597
rect 12750 18594 12756 18596
rect 11145 18592 12756 18594
rect 11145 18536 11150 18592
rect 11206 18536 12756 18592
rect 11145 18534 12756 18536
rect 11145 18531 11211 18534
rect 12750 18532 12756 18534
rect 12820 18532 12826 18596
rect 21541 18594 21607 18597
rect 23614 18594 23674 19048
rect 21541 18592 23674 18594
rect 21541 18536 21546 18592
rect 21602 18536 23674 18592
rect 21541 18534 23674 18536
rect 21541 18531 21607 18534
rect 4944 18528 5264 18529
rect 62 18458 122 18504
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 2681 18458 2747 18461
rect 4705 18458 4771 18461
rect 62 18456 4771 18458
rect 62 18400 2686 18456
rect 2742 18400 4710 18456
rect 4766 18400 4771 18456
rect 62 18398 4771 18400
rect 2681 18395 2747 18398
rect 4705 18395 4771 18398
rect 6310 18396 6316 18460
rect 6380 18458 6386 18460
rect 6453 18458 6519 18461
rect 6380 18456 6519 18458
rect 6380 18400 6458 18456
rect 6514 18400 6519 18456
rect 6380 18398 6519 18400
rect 6380 18396 6386 18398
rect 6453 18395 6519 18398
rect 6637 18458 6703 18461
rect 7833 18458 7899 18461
rect 6637 18456 7899 18458
rect 6637 18400 6642 18456
rect 6698 18400 7838 18456
rect 7894 18400 7899 18456
rect 6637 18398 7899 18400
rect 6637 18395 6703 18398
rect 7833 18395 7899 18398
rect 8334 18396 8340 18460
rect 8404 18458 8410 18460
rect 10593 18458 10659 18461
rect 8404 18456 10659 18458
rect 8404 18400 10598 18456
rect 10654 18400 10659 18456
rect 8404 18398 10659 18400
rect 8404 18396 8410 18398
rect 10593 18395 10659 18398
rect 19793 18458 19859 18461
rect 19926 18458 19932 18460
rect 19793 18456 19932 18458
rect 19793 18400 19798 18456
rect 19854 18400 19932 18456
rect 19793 18398 19932 18400
rect 19793 18395 19859 18398
rect 19926 18396 19932 18398
rect 19996 18396 20002 18460
rect 606 18260 612 18324
rect 676 18322 682 18324
rect 933 18322 999 18325
rect 676 18320 999 18322
rect 676 18264 938 18320
rect 994 18264 999 18320
rect 676 18262 999 18264
rect 676 18260 682 18262
rect 933 18259 999 18262
rect 1485 18322 1551 18325
rect 8702 18322 8708 18324
rect 1485 18320 8708 18322
rect 1485 18264 1490 18320
rect 1546 18264 8708 18320
rect 1485 18262 8708 18264
rect 1485 18259 1551 18262
rect 8702 18260 8708 18262
rect 8772 18260 8778 18324
rect 9489 18322 9555 18325
rect 13997 18322 14063 18325
rect 9489 18320 14063 18322
rect 9489 18264 9494 18320
rect 9550 18264 14002 18320
rect 14058 18264 14063 18320
rect 9489 18262 14063 18264
rect 9489 18259 9555 18262
rect 13997 18259 14063 18262
rect 15009 18322 15075 18325
rect 20713 18322 20779 18325
rect 15009 18320 20779 18322
rect 15009 18264 15014 18320
rect 15070 18264 20718 18320
rect 20774 18264 20779 18320
rect 15009 18262 20779 18264
rect 15009 18259 15075 18262
rect 20713 18259 20779 18262
rect 3734 18124 3740 18188
rect 3804 18186 3810 18188
rect 13537 18186 13603 18189
rect 20437 18186 20503 18189
rect 3804 18126 9460 18186
rect 3804 18124 3810 18126
rect 841 18050 907 18053
rect 974 18050 980 18052
rect 841 18048 980 18050
rect 841 17992 846 18048
rect 902 17992 980 18048
rect 841 17990 980 17992
rect 841 17987 907 17990
rect 974 17988 980 17990
rect 1044 17988 1050 18052
rect 2681 18050 2747 18053
rect 7833 18050 7899 18053
rect 2681 18048 7899 18050
rect 2681 17992 2686 18048
rect 2742 17992 7838 18048
rect 7894 17992 7899 18048
rect 2681 17990 7899 17992
rect 2681 17987 2747 17990
rect 7833 17987 7899 17990
rect 8518 17988 8524 18052
rect 8588 18050 8594 18052
rect 8753 18050 8819 18053
rect 8588 18048 8819 18050
rect 8588 17992 8758 18048
rect 8814 17992 8819 18048
rect 8588 17990 8819 17992
rect 9400 18050 9460 18126
rect 13537 18184 20503 18186
rect 13537 18128 13542 18184
rect 13598 18128 20442 18184
rect 20498 18128 20503 18184
rect 13537 18126 20503 18128
rect 13537 18123 13603 18126
rect 20437 18123 20503 18126
rect 15326 18050 15332 18052
rect 9400 17990 15332 18050
rect 8588 17988 8594 17990
rect 8753 17987 8819 17990
rect 15326 17988 15332 17990
rect 15396 17988 15402 18052
rect 15878 17988 15884 18052
rect 15948 18050 15954 18052
rect 16757 18050 16823 18053
rect 15948 18048 16823 18050
rect 15948 17992 16762 18048
rect 16818 17992 16823 18048
rect 15948 17990 16823 17992
rect 15948 17988 15954 17990
rect 16757 17987 16823 17990
rect 17534 17988 17540 18052
rect 17604 18050 17610 18052
rect 17861 18050 17927 18053
rect 17604 18048 17927 18050
rect 17604 17992 17866 18048
rect 17922 17992 17927 18048
rect 17604 17990 17927 17992
rect 17604 17988 17610 17990
rect 17861 17987 17927 17990
rect 8944 17984 9264 17985
rect 0 17916 480 17944
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 23520 17960 24000 18080
rect 16944 17919 17264 17920
rect 0 17852 60 17916
rect 124 17852 480 17916
rect 1342 17852 1348 17916
rect 1412 17914 1418 17916
rect 8753 17914 8819 17917
rect 1412 17912 8819 17914
rect 1412 17856 8758 17912
rect 8814 17856 8819 17912
rect 1412 17854 8819 17856
rect 1412 17852 1418 17854
rect 0 17824 480 17852
rect 8753 17851 8819 17854
rect 10317 17914 10383 17917
rect 13169 17914 13235 17917
rect 10317 17912 13235 17914
rect 10317 17856 10322 17912
rect 10378 17856 13174 17912
rect 13230 17856 13235 17912
rect 10317 17854 13235 17856
rect 10317 17851 10383 17854
rect 13169 17851 13235 17854
rect 13629 17914 13695 17917
rect 13997 17914 14063 17917
rect 13629 17912 14063 17914
rect 13629 17856 13634 17912
rect 13690 17856 14002 17912
rect 14058 17856 14063 17912
rect 13629 17854 14063 17856
rect 13629 17851 13695 17854
rect 13997 17851 14063 17854
rect 14222 17852 14228 17916
rect 14292 17914 14298 17916
rect 15009 17914 15075 17917
rect 14292 17912 15075 17914
rect 14292 17856 15014 17912
rect 15070 17856 15075 17912
rect 14292 17854 15075 17856
rect 14292 17852 14298 17854
rect 15009 17851 15075 17854
rect 62 17370 122 17824
rect 2814 17716 2820 17780
rect 2884 17778 2890 17780
rect 4061 17778 4127 17781
rect 2884 17776 4127 17778
rect 2884 17720 4066 17776
rect 4122 17720 4127 17776
rect 2884 17718 4127 17720
rect 2884 17716 2890 17718
rect 4061 17715 4127 17718
rect 4337 17778 4403 17781
rect 7005 17778 7071 17781
rect 4337 17776 7071 17778
rect 4337 17720 4342 17776
rect 4398 17720 7010 17776
rect 7066 17720 7071 17776
rect 4337 17718 7071 17720
rect 4337 17715 4403 17718
rect 7005 17715 7071 17718
rect 7373 17778 7439 17781
rect 8293 17778 8359 17781
rect 7373 17776 8359 17778
rect 7373 17720 7378 17776
rect 7434 17720 8298 17776
rect 8354 17720 8359 17776
rect 7373 17718 8359 17720
rect 7373 17715 7439 17718
rect 8293 17715 8359 17718
rect 8702 17716 8708 17780
rect 8772 17778 8778 17780
rect 14089 17778 14155 17781
rect 8772 17776 14155 17778
rect 8772 17720 14094 17776
rect 14150 17720 14155 17776
rect 8772 17718 14155 17720
rect 8772 17716 8778 17718
rect 14089 17715 14155 17718
rect 15101 17776 15167 17781
rect 15101 17720 15106 17776
rect 15162 17720 15167 17776
rect 15101 17715 15167 17720
rect 2998 17580 3004 17644
rect 3068 17642 3074 17644
rect 4654 17642 4660 17644
rect 3068 17582 4660 17642
rect 3068 17580 3074 17582
rect 4654 17580 4660 17582
rect 4724 17580 4730 17644
rect 7189 17642 7255 17645
rect 9029 17642 9095 17645
rect 7189 17640 9095 17642
rect 7189 17584 7194 17640
rect 7250 17584 9034 17640
rect 9090 17584 9095 17640
rect 7189 17582 9095 17584
rect 7189 17579 7255 17582
rect 9029 17579 9095 17582
rect 9305 17642 9371 17645
rect 9622 17642 9628 17644
rect 9305 17640 9628 17642
rect 9305 17584 9310 17640
rect 9366 17584 9628 17640
rect 9305 17582 9628 17584
rect 9305 17579 9371 17582
rect 9622 17580 9628 17582
rect 9692 17580 9698 17644
rect 14917 17642 14983 17645
rect 9768 17640 14983 17642
rect 9768 17584 14922 17640
rect 14978 17584 14983 17640
rect 9768 17582 14983 17584
rect 565 17506 631 17509
rect 790 17506 796 17508
rect 565 17504 796 17506
rect 565 17448 570 17504
rect 626 17448 796 17504
rect 565 17446 796 17448
rect 565 17443 631 17446
rect 790 17444 796 17446
rect 860 17444 866 17508
rect 2221 17506 2287 17509
rect 2221 17504 4170 17506
rect 2221 17448 2226 17504
rect 2282 17448 4170 17504
rect 2221 17446 4170 17448
rect 2221 17443 2287 17446
rect 289 17370 355 17373
rect 62 17368 355 17370
rect 62 17312 294 17368
rect 350 17312 355 17368
rect 62 17310 355 17312
rect 289 17307 355 17310
rect 657 17370 723 17373
rect 790 17370 796 17372
rect 657 17368 796 17370
rect 657 17312 662 17368
rect 718 17312 796 17368
rect 657 17310 796 17312
rect 657 17307 723 17310
rect 790 17308 796 17310
rect 860 17308 866 17372
rect 2405 17232 2471 17237
rect 2405 17176 2410 17232
rect 2466 17176 2471 17232
rect 2405 17171 2471 17176
rect 4110 17234 4170 17446
rect 5758 17444 5764 17508
rect 5828 17506 5834 17508
rect 8753 17506 8819 17509
rect 9768 17506 9828 17582
rect 14917 17579 14983 17582
rect 5828 17504 8819 17506
rect 5828 17448 8758 17504
rect 8814 17448 8819 17504
rect 5828 17446 8819 17448
rect 5828 17444 5834 17446
rect 8753 17443 8819 17446
rect 8894 17446 9828 17506
rect 14917 17506 14983 17509
rect 15104 17506 15164 17715
rect 14917 17504 15164 17506
rect 14917 17448 14922 17504
rect 14978 17448 15164 17504
rect 14917 17446 15164 17448
rect 21357 17506 21423 17509
rect 23614 17506 23674 17960
rect 21357 17504 23674 17506
rect 21357 17448 21362 17504
rect 21418 17448 23674 17504
rect 21357 17446 23674 17448
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 5352 17310 7436 17370
rect 5352 17234 5412 17310
rect 4110 17174 5412 17234
rect 7376 17234 7436 17310
rect 7598 17308 7604 17372
rect 7668 17370 7674 17372
rect 8894 17370 8954 17446
rect 14917 17443 14983 17446
rect 21357 17443 21423 17446
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 7668 17310 8954 17370
rect 7668 17308 7674 17310
rect 9438 17308 9444 17372
rect 9508 17370 9514 17372
rect 10685 17370 10751 17373
rect 9508 17368 10751 17370
rect 9508 17312 10690 17368
rect 10746 17312 10751 17368
rect 9508 17310 10751 17312
rect 9508 17308 9514 17310
rect 10685 17307 10751 17310
rect 9581 17234 9647 17237
rect 11646 17234 11652 17236
rect 7376 17232 11652 17234
rect 7376 17176 9586 17232
rect 9642 17176 11652 17232
rect 7376 17174 11652 17176
rect 9581 17171 9647 17174
rect 11646 17172 11652 17174
rect 11716 17172 11722 17236
rect 11789 17234 11855 17237
rect 12801 17234 12867 17237
rect 16021 17234 16087 17237
rect 11789 17232 11898 17234
rect 11789 17176 11794 17232
rect 11850 17176 11898 17232
rect 11789 17171 11898 17176
rect 12801 17232 16087 17234
rect 12801 17176 12806 17232
rect 12862 17176 16026 17232
rect 16082 17176 16087 17232
rect 12801 17174 16087 17176
rect 12801 17171 12867 17174
rect 16021 17171 16087 17174
rect 0 17096 480 17128
rect 0 17040 110 17096
rect 166 17040 480 17096
rect 0 17008 480 17040
rect 2221 17098 2287 17101
rect 2408 17098 2468 17171
rect 9489 17098 9555 17101
rect 2221 17096 9555 17098
rect 2221 17040 2226 17096
rect 2282 17040 9494 17096
rect 9550 17040 9555 17096
rect 2221 17038 9555 17040
rect 2221 17035 2287 17038
rect 9489 17035 9555 17038
rect 1209 16962 1275 16965
rect 1710 16962 1716 16964
rect 1209 16960 1716 16962
rect 1209 16904 1214 16960
rect 1270 16904 1716 16960
rect 1209 16902 1716 16904
rect 1209 16899 1275 16902
rect 1710 16900 1716 16902
rect 1780 16900 1786 16964
rect 3550 16900 3556 16964
rect 3620 16962 3626 16964
rect 4245 16962 4311 16965
rect 3620 16960 4311 16962
rect 3620 16904 4250 16960
rect 4306 16904 4311 16960
rect 3620 16902 4311 16904
rect 3620 16900 3626 16902
rect 4245 16899 4311 16902
rect 4470 16900 4476 16964
rect 4540 16962 4546 16964
rect 4889 16962 4955 16965
rect 4540 16960 4955 16962
rect 4540 16904 4894 16960
rect 4950 16904 4955 16960
rect 4540 16902 4955 16904
rect 4540 16900 4546 16902
rect 4889 16899 4955 16902
rect 5257 16962 5323 16965
rect 5390 16962 5396 16964
rect 5257 16960 5396 16962
rect 5257 16904 5262 16960
rect 5318 16904 5396 16960
rect 5257 16902 5396 16904
rect 5257 16899 5323 16902
rect 5390 16900 5396 16902
rect 5460 16900 5466 16964
rect 7230 16900 7236 16964
rect 7300 16962 7306 16964
rect 7465 16962 7531 16965
rect 7300 16960 7531 16962
rect 7300 16904 7470 16960
rect 7526 16904 7531 16960
rect 7300 16902 7531 16904
rect 11838 16962 11898 17171
rect 12617 17098 12683 17101
rect 14641 17098 14707 17101
rect 12617 17096 14707 17098
rect 12617 17040 12622 17096
rect 12678 17040 14646 17096
rect 14702 17040 14707 17096
rect 12617 17038 14707 17040
rect 12617 17035 12683 17038
rect 14641 17035 14707 17038
rect 12801 16962 12867 16965
rect 11838 16960 12867 16962
rect 11838 16904 12806 16960
rect 12862 16904 12867 16960
rect 11838 16902 12867 16904
rect 7300 16900 7306 16902
rect 7465 16899 7531 16902
rect 12801 16899 12867 16902
rect 13169 16962 13235 16965
rect 14958 16962 14964 16964
rect 13169 16960 14964 16962
rect 13169 16904 13174 16960
rect 13230 16904 14964 16960
rect 13169 16902 14964 16904
rect 13169 16899 13235 16902
rect 14958 16900 14964 16902
rect 15028 16900 15034 16964
rect 23520 16962 24000 16992
rect 23484 16960 24000 16962
rect 23484 16904 23570 16960
rect 23626 16904 24000 16960
rect 23484 16902 24000 16904
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 23520 16872 24000 16902
rect 16944 16831 17264 16832
rect 841 16826 907 16829
rect 841 16824 4170 16826
rect 841 16768 846 16824
rect 902 16768 4170 16824
rect 841 16766 4170 16768
rect 841 16763 907 16766
rect 54 16628 60 16692
rect 124 16690 130 16692
rect 657 16690 723 16693
rect 2037 16690 2103 16693
rect 124 16688 2103 16690
rect 124 16632 662 16688
rect 718 16632 2042 16688
rect 2098 16632 2103 16688
rect 124 16630 2103 16632
rect 4110 16690 4170 16766
rect 4286 16764 4292 16828
rect 4356 16826 4362 16828
rect 6085 16826 6151 16829
rect 11145 16826 11211 16829
rect 4356 16824 6151 16826
rect 4356 16768 6090 16824
rect 6146 16768 6151 16824
rect 4356 16766 6151 16768
rect 4356 16764 4362 16766
rect 6085 16763 6151 16766
rect 9630 16824 11211 16826
rect 9630 16768 11150 16824
rect 11206 16768 11211 16824
rect 9630 16766 11211 16768
rect 5993 16690 6059 16693
rect 4110 16688 6059 16690
rect 4110 16632 5998 16688
rect 6054 16632 6059 16688
rect 4110 16630 6059 16632
rect 124 16628 130 16630
rect 657 16627 723 16630
rect 2037 16627 2103 16630
rect 5993 16627 6059 16630
rect 6177 16690 6243 16693
rect 9630 16690 9690 16766
rect 11145 16763 11211 16766
rect 6177 16688 9690 16690
rect 6177 16632 6182 16688
rect 6238 16632 9690 16688
rect 6177 16630 9690 16632
rect 9765 16690 9831 16693
rect 11830 16690 11836 16692
rect 9765 16688 11836 16690
rect 9765 16632 9770 16688
rect 9826 16632 11836 16688
rect 9765 16630 11836 16632
rect 6177 16627 6243 16630
rect 9765 16627 9831 16630
rect 11830 16628 11836 16630
rect 11900 16628 11906 16692
rect 657 16554 723 16557
rect 6545 16554 6611 16557
rect 657 16552 6611 16554
rect 657 16496 662 16552
rect 718 16496 6550 16552
rect 6606 16496 6611 16552
rect 657 16494 6611 16496
rect 657 16491 723 16494
rect 6545 16491 6611 16494
rect 6678 16492 6684 16556
rect 6748 16554 6754 16556
rect 6913 16554 6979 16557
rect 6748 16552 6979 16554
rect 6748 16496 6918 16552
rect 6974 16496 6979 16552
rect 6748 16494 6979 16496
rect 6748 16492 6754 16494
rect 6913 16491 6979 16494
rect 7782 16492 7788 16556
rect 7852 16554 7858 16556
rect 13670 16554 13676 16556
rect 7852 16494 13676 16554
rect 7852 16492 7858 16494
rect 13670 16492 13676 16494
rect 13740 16492 13746 16556
rect 7281 16418 7347 16421
rect 8937 16418 9003 16421
rect 7281 16416 9003 16418
rect 7281 16360 7286 16416
rect 7342 16360 8942 16416
rect 8998 16360 9003 16416
rect 7281 16358 9003 16360
rect 7281 16355 7347 16358
rect 8937 16355 9003 16358
rect 9121 16418 9187 16421
rect 11973 16418 12039 16421
rect 9121 16416 12039 16418
rect 9121 16360 9126 16416
rect 9182 16360 11978 16416
rect 12034 16360 12039 16416
rect 9121 16358 12039 16360
rect 9121 16355 9187 16358
rect 11973 16355 12039 16358
rect 13353 16418 13419 16421
rect 20253 16418 20319 16421
rect 13353 16416 20319 16418
rect 13353 16360 13358 16416
rect 13414 16360 20258 16416
rect 20314 16360 20319 16416
rect 13353 16358 20319 16360
rect 13353 16355 13419 16358
rect 20253 16355 20319 16358
rect 4944 16352 5264 16353
rect 0 16280 480 16312
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 0 16224 110 16280
rect 166 16224 480 16280
rect 0 16192 480 16224
rect 2221 16282 2287 16285
rect 3918 16282 3924 16284
rect 2221 16280 3924 16282
rect 2221 16224 2226 16280
rect 2282 16224 3924 16280
rect 2221 16222 3924 16224
rect 2221 16219 2287 16222
rect 3918 16220 3924 16222
rect 3988 16220 3994 16284
rect 7005 16282 7071 16285
rect 7598 16282 7604 16284
rect 7005 16280 7604 16282
rect 7005 16224 7010 16280
rect 7066 16224 7604 16280
rect 7005 16222 7604 16224
rect 7005 16219 7071 16222
rect 7598 16220 7604 16222
rect 7668 16220 7674 16284
rect 8201 16282 8267 16285
rect 11462 16282 11468 16284
rect 8201 16280 11468 16282
rect 8201 16224 8206 16280
rect 8262 16224 11468 16280
rect 8201 16222 11468 16224
rect 8201 16219 8267 16222
rect 11462 16220 11468 16222
rect 11532 16220 11538 16284
rect 2313 16146 2379 16149
rect 4981 16146 5047 16149
rect 13813 16146 13879 16149
rect 2313 16144 5047 16146
rect 2313 16088 2318 16144
rect 2374 16088 4986 16144
rect 5042 16088 5047 16144
rect 2313 16086 5047 16088
rect 2313 16083 2379 16086
rect 4981 16083 5047 16086
rect 7284 16144 13879 16146
rect 7284 16088 13818 16144
rect 13874 16088 13879 16144
rect 7284 16086 13879 16088
rect 3233 16010 3299 16013
rect 7284 16010 7344 16086
rect 13813 16083 13879 16086
rect 13997 16010 14063 16013
rect 14406 16010 14412 16012
rect 3233 16008 7344 16010
rect 3233 15952 3238 16008
rect 3294 15952 7344 16008
rect 3233 15950 7344 15952
rect 8756 16008 14412 16010
rect 8756 15952 14002 16008
rect 14058 15952 14412 16008
rect 8756 15950 14412 15952
rect 3233 15947 3299 15950
rect 3141 15874 3207 15877
rect 4102 15874 4108 15876
rect 3141 15872 4108 15874
rect 3141 15816 3146 15872
rect 3202 15816 4108 15872
rect 3141 15814 4108 15816
rect 3141 15811 3207 15814
rect 4102 15812 4108 15814
rect 4172 15812 4178 15876
rect 5942 15812 5948 15876
rect 6012 15874 6018 15876
rect 6637 15874 6703 15877
rect 6012 15872 6703 15874
rect 6012 15816 6642 15872
rect 6698 15816 6703 15872
rect 6012 15814 6703 15816
rect 6012 15812 6018 15814
rect 6637 15811 6703 15814
rect 6821 15738 6887 15741
rect 8385 15738 8451 15741
rect 6821 15736 8451 15738
rect 6821 15680 6826 15736
rect 6882 15680 8390 15736
rect 8446 15680 8451 15736
rect 6821 15678 8451 15680
rect 6821 15675 6887 15678
rect 8385 15675 8451 15678
rect 2262 15540 2268 15604
rect 2332 15602 2338 15604
rect 8756 15602 8816 15950
rect 13997 15947 14063 15950
rect 14406 15948 14412 15950
rect 14476 15948 14482 16012
rect 12750 15812 12756 15876
rect 12820 15874 12826 15876
rect 12985 15874 13051 15877
rect 12820 15872 13051 15874
rect 12820 15816 12990 15872
rect 13046 15816 13051 15872
rect 12820 15814 13051 15816
rect 12820 15812 12826 15814
rect 12985 15811 13051 15814
rect 17350 15812 17356 15876
rect 17420 15874 17426 15876
rect 19333 15874 19399 15877
rect 17420 15872 19399 15874
rect 17420 15816 19338 15872
rect 19394 15816 19399 15872
rect 17420 15814 19399 15816
rect 17420 15812 17426 15814
rect 19333 15811 19399 15814
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 23520 15784 24000 15904
rect 16944 15743 17264 15744
rect 11421 15738 11487 15741
rect 14549 15738 14615 15741
rect 11421 15736 14615 15738
rect 11421 15680 11426 15736
rect 11482 15680 14554 15736
rect 14610 15680 14615 15736
rect 11421 15678 14615 15680
rect 11421 15675 11487 15678
rect 14549 15675 14615 15678
rect 19057 15738 19123 15741
rect 19333 15738 19399 15741
rect 19057 15736 19399 15738
rect 19057 15680 19062 15736
rect 19118 15680 19338 15736
rect 19394 15680 19399 15736
rect 19057 15678 19399 15680
rect 19057 15675 19123 15678
rect 19333 15675 19399 15678
rect 2332 15542 8816 15602
rect 2332 15540 2338 15542
rect 11094 15540 11100 15604
rect 11164 15602 11170 15604
rect 20713 15602 20779 15605
rect 11164 15600 20779 15602
rect 11164 15544 20718 15600
rect 20774 15544 20779 15600
rect 11164 15542 20779 15544
rect 11164 15540 11170 15542
rect 20713 15539 20779 15542
rect 0 15376 480 15496
rect 3693 15466 3759 15469
rect 3918 15466 3924 15468
rect 3693 15464 3924 15466
rect 3693 15408 3698 15464
rect 3754 15408 3924 15464
rect 3693 15406 3924 15408
rect 3693 15403 3759 15406
rect 3918 15404 3924 15406
rect 3988 15466 3994 15468
rect 4429 15466 4495 15469
rect 3988 15464 4495 15466
rect 3988 15408 4434 15464
rect 4490 15408 4495 15464
rect 3988 15406 4495 15408
rect 3988 15404 3994 15406
rect 4429 15403 4495 15406
rect 5349 15466 5415 15469
rect 7782 15466 7788 15468
rect 5349 15464 7788 15466
rect 5349 15408 5354 15464
rect 5410 15408 7788 15464
rect 5349 15406 7788 15408
rect 5349 15403 5415 15406
rect 7782 15404 7788 15406
rect 7852 15404 7858 15468
rect 8845 15466 8911 15469
rect 11278 15466 11284 15468
rect 8845 15464 11284 15466
rect 8845 15408 8850 15464
rect 8906 15408 11284 15464
rect 8845 15406 11284 15408
rect 8845 15403 8911 15406
rect 11278 15404 11284 15406
rect 11348 15404 11354 15468
rect 16941 15466 17007 15469
rect 18454 15466 18460 15468
rect 16941 15464 18460 15466
rect 16941 15408 16946 15464
rect 17002 15408 18460 15464
rect 16941 15406 18460 15408
rect 16941 15403 17007 15406
rect 18454 15404 18460 15406
rect 18524 15404 18530 15468
rect 19926 15404 19932 15468
rect 19996 15466 20002 15468
rect 23614 15466 23674 15784
rect 19996 15406 23674 15466
rect 19996 15404 20002 15406
rect 62 15194 122 15376
rect 7465 15330 7531 15333
rect 12617 15330 12683 15333
rect 7465 15328 12683 15330
rect 7465 15272 7470 15328
rect 7526 15272 12622 15328
rect 12678 15272 12683 15328
rect 7465 15270 12683 15272
rect 7465 15267 7531 15270
rect 12617 15267 12683 15270
rect 14733 15330 14799 15333
rect 18781 15330 18847 15333
rect 14733 15328 18847 15330
rect 14733 15272 14738 15328
rect 14794 15272 18786 15328
rect 18842 15272 18847 15328
rect 14733 15270 18847 15272
rect 14733 15267 14799 15270
rect 18781 15267 18847 15270
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 1577 15194 1643 15197
rect 62 15192 1643 15194
rect 62 15136 1582 15192
rect 1638 15136 1643 15192
rect 62 15134 1643 15136
rect 1577 15131 1643 15134
rect 2078 15132 2084 15196
rect 2148 15194 2154 15196
rect 2773 15194 2839 15197
rect 2148 15192 2839 15194
rect 2148 15136 2778 15192
rect 2834 15136 2839 15192
rect 2148 15134 2839 15136
rect 2148 15132 2154 15134
rect 2773 15131 2839 15134
rect 3233 15194 3299 15197
rect 3366 15194 3372 15196
rect 3233 15192 3372 15194
rect 3233 15136 3238 15192
rect 3294 15136 3372 15192
rect 3233 15134 3372 15136
rect 3233 15131 3299 15134
rect 3366 15132 3372 15134
rect 3436 15132 3442 15196
rect 7465 15194 7531 15197
rect 11421 15194 11487 15197
rect 7465 15192 11487 15194
rect 7465 15136 7470 15192
rect 7526 15136 11426 15192
rect 11482 15136 11487 15192
rect 7465 15134 11487 15136
rect 7465 15131 7531 15134
rect 11421 15131 11487 15134
rect 12566 15132 12572 15196
rect 12636 15194 12642 15196
rect 12801 15194 12867 15197
rect 12636 15192 12867 15194
rect 12636 15136 12806 15192
rect 12862 15136 12867 15192
rect 12636 15134 12867 15136
rect 12636 15132 12642 15134
rect 12801 15131 12867 15134
rect 16062 15132 16068 15196
rect 16132 15194 16138 15196
rect 17033 15194 17099 15197
rect 16132 15192 17099 15194
rect 16132 15136 17038 15192
rect 17094 15136 17099 15192
rect 16132 15134 17099 15136
rect 16132 15132 16138 15134
rect 17033 15131 17099 15134
rect 17718 15132 17724 15196
rect 17788 15194 17794 15196
rect 19885 15194 19951 15197
rect 17788 15192 19951 15194
rect 17788 15136 19890 15192
rect 19946 15136 19951 15192
rect 17788 15134 19951 15136
rect 17788 15132 17794 15134
rect 19885 15131 19951 15134
rect 1393 15058 1459 15061
rect 9305 15058 9371 15061
rect 10501 15058 10567 15061
rect 1393 15056 10567 15058
rect 1393 15000 1398 15056
rect 1454 15000 9310 15056
rect 9366 15000 10506 15056
rect 10562 15000 10567 15056
rect 1393 14998 10567 15000
rect 1393 14995 1459 14998
rect 9305 14995 9371 14998
rect 10501 14995 10567 14998
rect 10726 14996 10732 15060
rect 10796 15058 10802 15060
rect 18505 15058 18571 15061
rect 10796 15056 18571 15058
rect 10796 15000 18510 15056
rect 18566 15000 18571 15056
rect 10796 14998 18571 15000
rect 10796 14996 10802 14998
rect 18505 14995 18571 14998
rect 2078 14860 2084 14924
rect 2148 14922 2154 14924
rect 2221 14922 2287 14925
rect 2148 14920 2287 14922
rect 2148 14864 2226 14920
rect 2282 14864 2287 14920
rect 2148 14862 2287 14864
rect 2148 14860 2154 14862
rect 2221 14859 2287 14862
rect 4245 14922 4311 14925
rect 11053 14922 11119 14925
rect 4245 14920 11119 14922
rect 4245 14864 4250 14920
rect 4306 14864 11058 14920
rect 11114 14864 11119 14920
rect 4245 14862 11119 14864
rect 4245 14859 4311 14862
rect 11053 14859 11119 14862
rect 12014 14860 12020 14924
rect 12084 14922 12090 14924
rect 20161 14922 20227 14925
rect 12084 14920 20227 14922
rect 12084 14864 20166 14920
rect 20222 14864 20227 14920
rect 12084 14862 20227 14864
rect 12084 14860 12090 14862
rect 20161 14859 20227 14862
rect 3325 14788 3391 14789
rect 3325 14786 3372 14788
rect 3244 14784 3372 14786
rect 3436 14786 3442 14788
rect 6545 14786 6611 14789
rect 7833 14786 7899 14789
rect 3436 14784 6611 14786
rect 3244 14728 3330 14784
rect 3436 14728 6550 14784
rect 6606 14728 6611 14784
rect 3244 14726 3372 14728
rect 3325 14724 3372 14726
rect 3436 14726 6611 14728
rect 3436 14724 3442 14726
rect 3325 14723 3391 14724
rect 6545 14723 6611 14726
rect 7652 14784 7899 14786
rect 7652 14728 7838 14784
rect 7894 14728 7899 14784
rect 7652 14726 7899 14728
rect 0 14648 480 14680
rect 0 14592 18 14648
rect 74 14592 480 14648
rect 0 14560 480 14592
rect 5073 14650 5139 14653
rect 6126 14650 6132 14652
rect 5073 14648 6132 14650
rect 5073 14592 5078 14648
rect 5134 14592 6132 14648
rect 5073 14590 6132 14592
rect 5073 14587 5139 14590
rect 6126 14588 6132 14590
rect 6196 14650 6202 14652
rect 7652 14650 7712 14726
rect 7833 14723 7899 14726
rect 9673 14786 9739 14789
rect 13486 14786 13492 14788
rect 9673 14784 13492 14786
rect 9673 14728 9678 14784
rect 9734 14728 13492 14784
rect 9673 14726 13492 14728
rect 9673 14723 9739 14726
rect 13486 14724 13492 14726
rect 13556 14724 13562 14788
rect 15101 14786 15167 14789
rect 15510 14786 15516 14788
rect 15101 14784 15516 14786
rect 15101 14728 15106 14784
rect 15162 14728 15516 14784
rect 15101 14726 15516 14728
rect 15101 14723 15167 14726
rect 15510 14724 15516 14726
rect 15580 14724 15586 14788
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 23520 14696 24000 14816
rect 16944 14655 17264 14656
rect 6196 14590 7712 14650
rect 7833 14650 7899 14653
rect 8334 14650 8340 14652
rect 7833 14648 8340 14650
rect 7833 14592 7838 14648
rect 7894 14592 8340 14648
rect 7833 14590 8340 14592
rect 6196 14588 6202 14590
rect 7833 14587 7899 14590
rect 8334 14588 8340 14590
rect 8404 14588 8410 14652
rect 749 14514 815 14517
rect 7281 14514 7347 14517
rect 749 14512 7347 14514
rect 749 14456 754 14512
rect 810 14456 7286 14512
rect 7342 14456 7347 14512
rect 749 14454 7347 14456
rect 749 14451 815 14454
rect 7281 14451 7347 14454
rect 7414 14452 7420 14516
rect 7484 14514 7490 14516
rect 9673 14514 9739 14517
rect 7484 14512 9739 14514
rect 7484 14456 9678 14512
rect 9734 14456 9739 14512
rect 7484 14454 9739 14456
rect 7484 14452 7490 14454
rect 9673 14451 9739 14454
rect 15142 14452 15148 14516
rect 15212 14514 15218 14516
rect 20529 14514 20595 14517
rect 15212 14512 20595 14514
rect 15212 14456 20534 14512
rect 20590 14456 20595 14512
rect 15212 14454 20595 14456
rect 15212 14452 15218 14454
rect 20529 14451 20595 14454
rect 1577 14378 1643 14381
rect 9765 14378 9831 14381
rect 15193 14378 15259 14381
rect 19241 14378 19307 14381
rect 1577 14376 9831 14378
rect 1577 14320 1582 14376
rect 1638 14320 9770 14376
rect 9826 14320 9831 14376
rect 1577 14318 9831 14320
rect 1577 14315 1643 14318
rect 9765 14315 9831 14318
rect 9952 14376 15259 14378
rect 9952 14320 15198 14376
rect 15254 14320 15259 14376
rect 9952 14318 15259 14320
rect 1945 14242 2011 14245
rect 2446 14242 2452 14244
rect 1945 14240 2452 14242
rect 1945 14184 1950 14240
rect 2006 14184 2452 14240
rect 1945 14182 2452 14184
rect 1945 14179 2011 14182
rect 2446 14180 2452 14182
rect 2516 14180 2522 14244
rect 2957 14242 3023 14245
rect 3182 14242 3188 14244
rect 2957 14240 3188 14242
rect 2957 14184 2962 14240
rect 3018 14184 3188 14240
rect 2957 14182 3188 14184
rect 2957 14179 3023 14182
rect 3182 14180 3188 14182
rect 3252 14180 3258 14244
rect 3550 14180 3556 14244
rect 3620 14242 3626 14244
rect 3693 14242 3759 14245
rect 3620 14240 3759 14242
rect 3620 14184 3698 14240
rect 3754 14184 3759 14240
rect 3620 14182 3759 14184
rect 3620 14180 3626 14182
rect 3693 14179 3759 14182
rect 4470 14180 4476 14244
rect 4540 14180 4546 14244
rect 6545 14242 6611 14245
rect 9952 14242 10012 14318
rect 15193 14315 15259 14318
rect 16438 14376 19307 14378
rect 16438 14320 19246 14376
rect 19302 14320 19307 14376
rect 16438 14318 19307 14320
rect 6545 14240 10012 14242
rect 6545 14184 6550 14240
rect 6606 14184 10012 14240
rect 6545 14182 10012 14184
rect 4478 14109 4538 14180
rect 6545 14179 6611 14182
rect 10542 14180 10548 14244
rect 10612 14242 10618 14244
rect 12249 14242 12315 14245
rect 10612 14240 12315 14242
rect 10612 14184 12254 14240
rect 12310 14184 12315 14240
rect 10612 14182 12315 14184
rect 10612 14180 10618 14182
rect 12249 14179 12315 14182
rect 15929 14242 15995 14245
rect 16246 14242 16252 14244
rect 15929 14240 16252 14242
rect 15929 14184 15934 14240
rect 15990 14184 16252 14240
rect 15929 14182 16252 14184
rect 15929 14179 15995 14182
rect 16246 14180 16252 14182
rect 16316 14180 16322 14244
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 2405 14106 2471 14109
rect 2630 14106 2636 14108
rect 2405 14104 2636 14106
rect 2405 14048 2410 14104
rect 2466 14048 2636 14104
rect 2405 14046 2636 14048
rect 2405 14043 2471 14046
rect 2630 14044 2636 14046
rect 2700 14044 2706 14108
rect 4429 14104 4538 14109
rect 6862 14106 6868 14108
rect 4429 14048 4434 14104
rect 4490 14048 4538 14104
rect 4429 14046 4538 14048
rect 5582 14046 6868 14106
rect 4429 14043 4495 14046
rect 4981 13970 5047 13973
rect 5582 13970 5642 14046
rect 6862 14044 6868 14046
rect 6932 14044 6938 14108
rect 9673 14106 9739 14109
rect 12198 14106 12204 14108
rect 9673 14104 12204 14106
rect 9673 14048 9678 14104
rect 9734 14048 12204 14104
rect 9673 14046 12204 14048
rect 9673 14043 9739 14046
rect 12198 14044 12204 14046
rect 12268 14044 12274 14108
rect 15929 14106 15995 14109
rect 16438 14106 16498 14318
rect 19241 14315 19307 14318
rect 16614 14180 16620 14244
rect 16684 14242 16690 14244
rect 19190 14242 19196 14244
rect 16684 14182 19196 14242
rect 16684 14180 16690 14182
rect 19190 14180 19196 14182
rect 19260 14180 19266 14244
rect 22737 14242 22803 14245
rect 23614 14242 23674 14696
rect 22737 14240 23674 14242
rect 22737 14184 22742 14240
rect 22798 14184 23674 14240
rect 22737 14182 23674 14184
rect 22737 14179 22803 14182
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 15929 14104 16498 14106
rect 15929 14048 15934 14104
rect 15990 14048 16498 14104
rect 15929 14046 16498 14048
rect 15929 14043 15995 14046
rect 16614 14044 16620 14108
rect 16684 14106 16690 14108
rect 16757 14106 16823 14109
rect 16684 14104 16823 14106
rect 16684 14048 16762 14104
rect 16818 14048 16823 14104
rect 16684 14046 16823 14048
rect 16684 14044 16690 14046
rect 16757 14043 16823 14046
rect 4981 13968 5642 13970
rect 4981 13912 4986 13968
rect 5042 13912 5642 13968
rect 4981 13910 5642 13912
rect 4981 13907 5047 13910
rect 6494 13908 6500 13972
rect 6564 13908 6570 13972
rect 7005 13970 7071 13973
rect 7230 13970 7236 13972
rect 7005 13968 7236 13970
rect 7005 13912 7010 13968
rect 7066 13912 7236 13968
rect 7005 13910 7236 13912
rect 0 13836 480 13864
rect 0 13772 60 13836
rect 124 13772 480 13836
rect 0 13744 480 13772
rect 3509 13834 3575 13837
rect 6502 13834 6562 13908
rect 7005 13907 7071 13910
rect 7230 13908 7236 13910
rect 7300 13908 7306 13972
rect 9305 13970 9371 13973
rect 9305 13968 9690 13970
rect 9305 13912 9310 13968
rect 9366 13912 9690 13968
rect 9305 13910 9690 13912
rect 9305 13907 9371 13910
rect 7414 13834 7420 13836
rect 3509 13832 7420 13834
rect 3509 13776 3514 13832
rect 3570 13776 7420 13832
rect 3509 13774 7420 13776
rect 3509 13771 3575 13774
rect 6456 13770 6562 13774
rect 7414 13772 7420 13774
rect 7484 13834 7490 13836
rect 9630 13834 9690 13910
rect 10174 13908 10180 13972
rect 10244 13970 10250 13972
rect 11329 13970 11395 13973
rect 10244 13968 11395 13970
rect 10244 13912 11334 13968
rect 11390 13912 11395 13968
rect 10244 13910 11395 13912
rect 10244 13908 10250 13910
rect 11329 13907 11395 13910
rect 12382 13908 12388 13972
rect 12452 13970 12458 13972
rect 13353 13970 13419 13973
rect 12452 13968 13419 13970
rect 12452 13912 13358 13968
rect 13414 13912 13419 13968
rect 12452 13910 13419 13912
rect 12452 13908 12458 13910
rect 13353 13907 13419 13910
rect 14038 13908 14044 13972
rect 14108 13970 14114 13972
rect 14181 13970 14247 13973
rect 14108 13968 14247 13970
rect 14108 13912 14186 13968
rect 14242 13912 14247 13968
rect 14108 13910 14247 13912
rect 14108 13908 14114 13910
rect 14181 13907 14247 13910
rect 14549 13970 14615 13973
rect 18873 13970 18939 13973
rect 14549 13968 18939 13970
rect 14549 13912 14554 13968
rect 14610 13912 18878 13968
rect 18934 13912 18939 13968
rect 14549 13910 18939 13912
rect 14549 13907 14615 13910
rect 18873 13907 18939 13910
rect 18045 13834 18111 13837
rect 7484 13774 9506 13834
rect 9630 13832 18111 13834
rect 9630 13776 18050 13832
rect 18106 13776 18111 13832
rect 9630 13774 18111 13776
rect 7484 13772 7490 13774
rect 54 13636 60 13700
rect 124 13698 130 13700
rect 2773 13698 2839 13701
rect 124 13696 2839 13698
rect 124 13640 2778 13696
rect 2834 13640 2839 13696
rect 124 13638 2839 13640
rect 124 13636 130 13638
rect 2773 13635 2839 13638
rect 3734 13636 3740 13700
rect 3804 13698 3810 13700
rect 4470 13698 4476 13700
rect 3804 13638 4476 13698
rect 3804 13636 3810 13638
rect 4470 13636 4476 13638
rect 4540 13636 4546 13700
rect 4654 13636 4660 13700
rect 4724 13698 4730 13700
rect 5942 13698 5948 13700
rect 4724 13638 5948 13698
rect 4724 13636 4730 13638
rect 5942 13636 5948 13638
rect 6012 13636 6018 13700
rect 6310 13636 6316 13700
rect 6380 13698 6386 13700
rect 6456 13698 6516 13770
rect 6380 13638 6516 13698
rect 9446 13698 9506 13774
rect 18045 13771 18111 13774
rect 10685 13698 10751 13701
rect 9446 13696 10751 13698
rect 9446 13640 10690 13696
rect 10746 13640 10751 13696
rect 9446 13638 10751 13640
rect 6380 13636 6386 13638
rect 10685 13635 10751 13638
rect 15878 13636 15884 13700
rect 15948 13698 15954 13700
rect 16021 13698 16087 13701
rect 23520 13698 24000 13728
rect 15948 13696 16087 13698
rect 15948 13640 16026 13696
rect 16082 13640 16087 13696
rect 15948 13638 16087 13640
rect 23484 13696 24000 13698
rect 23484 13640 23570 13696
rect 23626 13640 24000 13696
rect 23484 13638 24000 13640
rect 15948 13636 15954 13638
rect 16021 13635 16087 13638
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 23520 13608 24000 13638
rect 16944 13567 17264 13568
rect 3734 13500 3740 13564
rect 3804 13562 3810 13564
rect 3877 13562 3943 13565
rect 3804 13560 3943 13562
rect 3804 13504 3882 13560
rect 3938 13504 3943 13560
rect 3804 13502 3943 13504
rect 3804 13500 3810 13502
rect 3877 13499 3943 13502
rect 4654 13500 4660 13564
rect 4724 13562 4730 13564
rect 5349 13562 5415 13565
rect 4724 13560 5415 13562
rect 4724 13504 5354 13560
rect 5410 13504 5415 13560
rect 4724 13502 5415 13504
rect 4724 13500 4730 13502
rect 5349 13499 5415 13502
rect 7230 13500 7236 13564
rect 7300 13562 7306 13564
rect 7598 13562 7604 13564
rect 7300 13502 7604 13562
rect 7300 13500 7306 13502
rect 7598 13500 7604 13502
rect 7668 13500 7674 13564
rect 8109 13562 8175 13565
rect 8334 13562 8340 13564
rect 8109 13560 8340 13562
rect 8109 13504 8114 13560
rect 8170 13504 8340 13560
rect 8109 13502 8340 13504
rect 8109 13499 8175 13502
rect 8334 13500 8340 13502
rect 8404 13500 8410 13564
rect 14549 13562 14615 13565
rect 9400 13560 14615 13562
rect 9400 13504 14554 13560
rect 14610 13504 14615 13560
rect 9400 13502 14615 13504
rect 4613 13426 4679 13429
rect 4613 13424 6516 13426
rect 4613 13368 4618 13424
rect 4674 13368 6516 13424
rect 4613 13366 6516 13368
rect 4613 13363 4679 13366
rect 1117 13290 1183 13293
rect 1342 13290 1348 13292
rect 1117 13288 1348 13290
rect 1117 13232 1122 13288
rect 1178 13232 1348 13288
rect 1117 13230 1348 13232
rect 1117 13227 1183 13230
rect 1342 13228 1348 13230
rect 1412 13228 1418 13292
rect 3182 13228 3188 13292
rect 3252 13290 3258 13292
rect 4705 13290 4771 13293
rect 3252 13288 4771 13290
rect 3252 13232 4710 13288
rect 4766 13232 4771 13288
rect 3252 13230 4771 13232
rect 6456 13290 6516 13366
rect 7598 13364 7604 13428
rect 7668 13426 7674 13428
rect 8017 13426 8083 13429
rect 9400 13426 9460 13502
rect 14549 13499 14615 13502
rect 14774 13500 14780 13564
rect 14844 13562 14850 13564
rect 16665 13562 16731 13565
rect 14844 13560 16731 13562
rect 14844 13504 16670 13560
rect 16726 13504 16731 13560
rect 14844 13502 16731 13504
rect 14844 13500 14850 13502
rect 16665 13499 16731 13502
rect 18086 13500 18092 13564
rect 18156 13562 18162 13564
rect 18597 13562 18663 13565
rect 18156 13560 18663 13562
rect 18156 13504 18602 13560
rect 18658 13504 18663 13560
rect 18156 13502 18663 13504
rect 18156 13500 18162 13502
rect 18597 13499 18663 13502
rect 7668 13424 8083 13426
rect 7668 13368 8022 13424
rect 8078 13368 8083 13424
rect 7668 13366 8083 13368
rect 7668 13364 7674 13366
rect 8017 13363 8083 13366
rect 8388 13366 9460 13426
rect 9581 13426 9647 13429
rect 14641 13426 14707 13429
rect 9581 13424 14707 13426
rect 9581 13368 9586 13424
rect 9642 13368 14646 13424
rect 14702 13368 14707 13424
rect 9581 13366 14707 13368
rect 8388 13290 8448 13366
rect 9581 13363 9647 13366
rect 14641 13363 14707 13366
rect 17902 13364 17908 13428
rect 17972 13426 17978 13428
rect 17972 13366 20178 13426
rect 17972 13364 17978 13366
rect 6456 13230 8448 13290
rect 3252 13228 3258 13230
rect 4705 13227 4771 13230
rect 8518 13228 8524 13292
rect 8588 13290 8594 13292
rect 9990 13290 9996 13292
rect 8588 13230 9996 13290
rect 8588 13228 8594 13230
rect 9990 13228 9996 13230
rect 10060 13228 10066 13292
rect 15878 13228 15884 13292
rect 15948 13290 15954 13292
rect 18413 13290 18479 13293
rect 20118 13292 20178 13366
rect 15948 13288 18479 13290
rect 15948 13232 18418 13288
rect 18474 13232 18479 13288
rect 15948 13230 18479 13232
rect 15948 13228 15954 13230
rect 18413 13227 18479 13230
rect 20110 13228 20116 13292
rect 20180 13290 20186 13292
rect 20897 13290 20963 13293
rect 20180 13288 20963 13290
rect 20180 13232 20902 13288
rect 20958 13232 20963 13288
rect 20180 13230 20963 13232
rect 20180 13228 20186 13230
rect 20897 13227 20963 13230
rect 5809 13152 5875 13157
rect 5809 13096 5814 13152
rect 5870 13096 5875 13152
rect 5809 13091 5875 13096
rect 10542 13092 10548 13156
rect 10612 13154 10618 13156
rect 11421 13154 11487 13157
rect 10612 13152 11487 13154
rect 10612 13096 11426 13152
rect 11482 13096 11487 13152
rect 10612 13094 11487 13096
rect 10612 13092 10618 13094
rect 11421 13091 11487 13094
rect 15510 13092 15516 13156
rect 15580 13154 15586 13156
rect 19977 13154 20043 13157
rect 20805 13154 20871 13157
rect 15580 13152 20871 13154
rect 15580 13096 19982 13152
rect 20038 13096 20810 13152
rect 20866 13096 20871 13152
rect 15580 13094 20871 13096
rect 15580 13092 15586 13094
rect 19977 13091 20043 13094
rect 20805 13091 20871 13094
rect 4944 13088 5264 13089
rect 0 12928 480 13048
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 5441 13018 5507 13021
rect 5574 13018 5580 13020
rect 5441 13016 5580 13018
rect 5441 12960 5446 13016
rect 5502 12960 5580 13016
rect 5441 12958 5580 12960
rect 5441 12955 5507 12958
rect 5574 12956 5580 12958
rect 5644 12956 5650 13020
rect 62 12613 122 12928
rect 238 12820 244 12884
rect 308 12882 314 12884
rect 381 12882 447 12885
rect 308 12880 447 12882
rect 308 12824 386 12880
rect 442 12824 447 12880
rect 308 12822 447 12824
rect 308 12820 314 12822
rect 381 12819 447 12822
rect 4797 12882 4863 12885
rect 5812 12882 5872 13091
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 9765 13018 9831 13021
rect 10174 13018 10180 13020
rect 9765 13016 10180 13018
rect 9765 12960 9770 13016
rect 9826 12960 10180 13016
rect 9765 12958 10180 12960
rect 9765 12955 9831 12958
rect 10174 12956 10180 12958
rect 10244 12956 10250 13020
rect 14365 13018 14431 13021
rect 18597 13018 18663 13021
rect 14365 13016 18663 13018
rect 14365 12960 14370 13016
rect 14426 12960 18602 13016
rect 18658 12960 18663 13016
rect 14365 12958 18663 12960
rect 14365 12955 14431 12958
rect 18597 12955 18663 12958
rect 4797 12880 5872 12882
rect 4797 12824 4802 12880
rect 4858 12824 5872 12880
rect 4797 12822 5872 12824
rect 6177 12882 6243 12885
rect 8937 12882 9003 12885
rect 6177 12880 9003 12882
rect 6177 12824 6182 12880
rect 6238 12824 8942 12880
rect 8998 12824 9003 12880
rect 6177 12822 9003 12824
rect 4797 12819 4863 12822
rect 6177 12819 6243 12822
rect 8937 12819 9003 12822
rect 10777 12882 10843 12885
rect 13721 12882 13787 12885
rect 10777 12880 13787 12882
rect 10777 12824 10782 12880
rect 10838 12824 13726 12880
rect 13782 12824 13787 12880
rect 10777 12822 13787 12824
rect 10777 12819 10843 12822
rect 13721 12819 13787 12822
rect 2129 12746 2195 12749
rect 2814 12746 2820 12748
rect 2129 12744 2820 12746
rect 2129 12688 2134 12744
rect 2190 12688 2820 12744
rect 2129 12686 2820 12688
rect 2129 12683 2195 12686
rect 2814 12684 2820 12686
rect 2884 12746 2890 12748
rect 3417 12746 3483 12749
rect 2884 12744 3483 12746
rect 2884 12688 3422 12744
rect 3478 12688 3483 12744
rect 2884 12686 3483 12688
rect 2884 12684 2890 12686
rect 3417 12683 3483 12686
rect 4102 12684 4108 12748
rect 4172 12746 4178 12748
rect 4981 12746 5047 12749
rect 4172 12744 5047 12746
rect 4172 12688 4986 12744
rect 5042 12688 5047 12744
rect 4172 12686 5047 12688
rect 4172 12684 4178 12686
rect 4981 12683 5047 12686
rect 5625 12746 5691 12749
rect 8334 12746 8340 12748
rect 5625 12744 8340 12746
rect 5625 12688 5630 12744
rect 5686 12688 8340 12744
rect 5625 12686 8340 12688
rect 5625 12683 5691 12686
rect 8334 12684 8340 12686
rect 8404 12684 8410 12748
rect 8569 12746 8635 12749
rect 8702 12746 8708 12748
rect 8569 12744 8708 12746
rect 8569 12688 8574 12744
rect 8630 12688 8708 12744
rect 8569 12686 8708 12688
rect 8569 12683 8635 12686
rect 8702 12684 8708 12686
rect 8772 12684 8778 12748
rect 9121 12746 9187 12749
rect 9397 12746 9463 12749
rect 9121 12744 9463 12746
rect 9121 12688 9126 12744
rect 9182 12688 9402 12744
rect 9458 12688 9463 12744
rect 9121 12686 9463 12688
rect 9121 12683 9187 12686
rect 9397 12683 9463 12686
rect 9990 12684 9996 12748
rect 10060 12746 10066 12748
rect 12341 12746 12407 12749
rect 10060 12744 12407 12746
rect 10060 12688 12346 12744
rect 12402 12688 12407 12744
rect 10060 12686 12407 12688
rect 10060 12684 10066 12686
rect 12341 12683 12407 12686
rect 16798 12684 16804 12748
rect 16868 12746 16874 12748
rect 22277 12746 22343 12749
rect 16868 12744 22343 12746
rect 16868 12688 22282 12744
rect 22338 12688 22343 12744
rect 16868 12686 22343 12688
rect 16868 12684 16874 12686
rect 22277 12683 22343 12686
rect 13 12608 122 12613
rect 13 12552 18 12608
rect 74 12552 122 12608
rect 13 12550 122 12552
rect 1761 12610 1827 12613
rect 2814 12610 2820 12612
rect 1761 12608 2820 12610
rect 1761 12552 1766 12608
rect 1822 12552 2820 12608
rect 1761 12550 2820 12552
rect 13 12547 79 12550
rect 1761 12547 1827 12550
rect 2814 12548 2820 12550
rect 2884 12610 2890 12612
rect 8385 12610 8451 12613
rect 2884 12608 8451 12610
rect 2884 12552 8390 12608
rect 8446 12552 8451 12608
rect 2884 12550 8451 12552
rect 2884 12548 2890 12550
rect 8385 12547 8451 12550
rect 9622 12548 9628 12612
rect 9692 12610 9698 12612
rect 10961 12610 11027 12613
rect 11697 12610 11763 12613
rect 9692 12608 11763 12610
rect 9692 12552 10966 12608
rect 11022 12552 11702 12608
rect 11758 12552 11763 12608
rect 9692 12550 11763 12552
rect 9692 12548 9698 12550
rect 10961 12547 11027 12550
rect 11697 12547 11763 12550
rect 12433 12610 12499 12613
rect 13169 12610 13235 12613
rect 12433 12608 13235 12610
rect 12433 12552 12438 12608
rect 12494 12552 13174 12608
rect 13230 12552 13235 12608
rect 12433 12550 13235 12552
rect 12433 12547 12499 12550
rect 13169 12547 13235 12550
rect 14958 12548 14964 12612
rect 15028 12610 15034 12612
rect 16021 12610 16087 12613
rect 15028 12608 16087 12610
rect 15028 12552 16026 12608
rect 16082 12552 16087 12608
rect 15028 12550 16087 12552
rect 15028 12548 15034 12550
rect 16021 12547 16087 12550
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 23520 12520 24000 12640
rect 16944 12479 17264 12480
rect 3141 12472 3207 12477
rect 3141 12416 3146 12472
rect 3202 12416 3207 12472
rect 3141 12411 3207 12416
rect 4153 12474 4219 12477
rect 5625 12474 5691 12477
rect 8385 12474 8451 12477
rect 4153 12472 5691 12474
rect 4153 12416 4158 12472
rect 4214 12416 5630 12472
rect 5686 12416 5691 12472
rect 4153 12414 5691 12416
rect 4153 12411 4219 12414
rect 5625 12411 5691 12414
rect 5950 12472 8451 12474
rect 5950 12416 8390 12472
rect 8446 12416 8451 12472
rect 5950 12414 8451 12416
rect 0 12340 480 12368
rect 0 12276 60 12340
rect 124 12276 480 12340
rect 0 12248 480 12276
rect 1209 12338 1275 12341
rect 1342 12338 1348 12340
rect 1209 12336 1348 12338
rect 1209 12280 1214 12336
rect 1270 12280 1348 12336
rect 1209 12278 1348 12280
rect 1209 12275 1275 12278
rect 1342 12276 1348 12278
rect 1412 12276 1418 12340
rect 3144 12338 3204 12411
rect 3550 12338 3556 12340
rect 3144 12278 3556 12338
rect 3550 12276 3556 12278
rect 3620 12338 3626 12340
rect 5950 12338 6010 12414
rect 8385 12411 8451 12414
rect 12433 12474 12499 12477
rect 12566 12474 12572 12476
rect 12433 12472 12572 12474
rect 12433 12416 12438 12472
rect 12494 12416 12572 12472
rect 12433 12414 12572 12416
rect 12433 12411 12499 12414
rect 12566 12412 12572 12414
rect 12636 12474 12642 12476
rect 12985 12474 13051 12477
rect 12636 12472 13051 12474
rect 12636 12416 12990 12472
rect 13046 12416 13051 12472
rect 12636 12414 13051 12416
rect 12636 12412 12642 12414
rect 12985 12411 13051 12414
rect 14590 12412 14596 12476
rect 14660 12474 14666 12476
rect 14917 12474 14983 12477
rect 14660 12472 14983 12474
rect 14660 12416 14922 12472
rect 14978 12416 14983 12472
rect 14660 12414 14983 12416
rect 14660 12412 14666 12414
rect 14917 12411 14983 12414
rect 15561 12474 15627 12477
rect 16062 12474 16068 12476
rect 15561 12472 16068 12474
rect 15561 12416 15566 12472
rect 15622 12416 16068 12472
rect 15561 12414 16068 12416
rect 15561 12411 15627 12414
rect 16062 12412 16068 12414
rect 16132 12412 16138 12476
rect 3620 12278 6010 12338
rect 3620 12276 3626 12278
rect 6862 12276 6868 12340
rect 6932 12338 6938 12340
rect 7966 12338 7972 12340
rect 6932 12278 7972 12338
rect 6932 12276 6938 12278
rect 7966 12276 7972 12278
rect 8036 12276 8042 12340
rect 9121 12338 9187 12341
rect 10041 12338 10107 12341
rect 9121 12336 10107 12338
rect 9121 12280 9126 12336
rect 9182 12280 10046 12336
rect 10102 12280 10107 12336
rect 9121 12278 10107 12280
rect 9121 12275 9187 12278
rect 10041 12275 10107 12278
rect 10358 12276 10364 12340
rect 10428 12338 10434 12340
rect 11145 12338 11211 12341
rect 10428 12336 11211 12338
rect 10428 12280 11150 12336
rect 11206 12280 11211 12336
rect 10428 12278 11211 12280
rect 10428 12276 10434 12278
rect 11145 12275 11211 12278
rect 18454 12276 18460 12340
rect 18524 12338 18530 12340
rect 19885 12338 19951 12341
rect 18524 12336 19951 12338
rect 18524 12280 19890 12336
rect 19946 12280 19951 12336
rect 18524 12278 19951 12280
rect 18524 12276 18530 12278
rect 19885 12275 19951 12278
rect 20662 12276 20668 12340
rect 20732 12338 20738 12340
rect 21265 12338 21331 12341
rect 20732 12336 21331 12338
rect 20732 12280 21270 12336
rect 21326 12280 21331 12336
rect 20732 12278 21331 12280
rect 20732 12276 20738 12278
rect 21265 12275 21331 12278
rect 9857 12202 9923 12205
rect 568 12200 9923 12202
rect 568 12144 9862 12200
rect 9918 12144 9923 12200
rect 568 12142 9923 12144
rect 54 12004 60 12068
rect 124 12066 130 12068
rect 568 12066 628 12142
rect 9857 12139 9923 12142
rect 10501 12202 10567 12205
rect 21633 12202 21699 12205
rect 10501 12200 21699 12202
rect 10501 12144 10506 12200
rect 10562 12144 21638 12200
rect 21694 12144 21699 12200
rect 10501 12142 21699 12144
rect 10501 12139 10567 12142
rect 21633 12139 21699 12142
rect 124 12006 628 12066
rect 1945 12066 2011 12069
rect 3918 12066 3924 12068
rect 1945 12064 3924 12066
rect 1945 12008 1950 12064
rect 2006 12008 3924 12064
rect 1945 12006 3924 12008
rect 124 12004 130 12006
rect 1945 12003 2011 12006
rect 3918 12004 3924 12006
rect 3988 12004 3994 12068
rect 4102 12004 4108 12068
rect 4172 12066 4178 12068
rect 4337 12066 4403 12069
rect 4172 12064 4403 12066
rect 4172 12008 4342 12064
rect 4398 12008 4403 12064
rect 4172 12006 4403 12008
rect 4172 12004 4178 12006
rect 4337 12003 4403 12006
rect 6269 12066 6335 12069
rect 7966 12066 7972 12068
rect 6269 12064 7972 12066
rect 6269 12008 6274 12064
rect 6330 12008 7972 12064
rect 6269 12006 7972 12008
rect 6269 12003 6335 12006
rect 7966 12004 7972 12006
rect 8036 12004 8042 12068
rect 8385 12066 8451 12069
rect 8518 12066 8524 12068
rect 8385 12064 8524 12066
rect 8385 12008 8390 12064
rect 8446 12008 8524 12064
rect 8385 12006 8524 12008
rect 8385 12003 8451 12006
rect 8518 12004 8524 12006
rect 8588 12004 8594 12068
rect 8753 12066 8819 12069
rect 9438 12066 9444 12068
rect 8753 12064 9444 12066
rect 8753 12008 8758 12064
rect 8814 12008 9444 12064
rect 8753 12006 9444 12008
rect 8753 12003 8819 12006
rect 9438 12004 9444 12006
rect 9508 12004 9514 12068
rect 10174 12004 10180 12068
rect 10244 12066 10250 12068
rect 10910 12066 10916 12068
rect 10244 12006 10916 12066
rect 10244 12004 10250 12006
rect 10910 12004 10916 12006
rect 10980 12004 10986 12068
rect 12341 12066 12407 12069
rect 12566 12066 12572 12068
rect 12341 12064 12572 12066
rect 12341 12008 12346 12064
rect 12402 12008 12572 12064
rect 12341 12006 12572 12008
rect 12341 12003 12407 12006
rect 12566 12004 12572 12006
rect 12636 12004 12642 12068
rect 21357 12066 21423 12069
rect 23614 12066 23674 12520
rect 21357 12064 23674 12066
rect 21357 12008 21362 12064
rect 21418 12008 23674 12064
rect 21357 12006 23674 12008
rect 21357 12003 21423 12006
rect 4944 12000 5264 12001
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 13 11930 79 11933
rect 3550 11930 3556 11932
rect 13 11928 3556 11930
rect 13 11872 18 11928
rect 74 11872 3556 11928
rect 13 11870 3556 11872
rect 13 11867 79 11870
rect 3550 11868 3556 11870
rect 3620 11868 3626 11932
rect 4337 11930 4403 11933
rect 4521 11930 4587 11933
rect 4337 11928 4587 11930
rect 4337 11872 4342 11928
rect 4398 11872 4526 11928
rect 4582 11872 4587 11928
rect 4337 11870 4587 11872
rect 4337 11867 4403 11870
rect 4521 11867 4587 11870
rect 5809 11930 5875 11933
rect 9949 11930 10015 11933
rect 5809 11928 10015 11930
rect 5809 11872 5814 11928
rect 5870 11872 9954 11928
rect 10010 11872 10015 11928
rect 5809 11870 10015 11872
rect 5809 11867 5875 11870
rect 9949 11867 10015 11870
rect 10869 11930 10935 11933
rect 12750 11930 12756 11932
rect 10869 11928 12756 11930
rect 10869 11872 10874 11928
rect 10930 11872 12756 11928
rect 10869 11870 12756 11872
rect 10869 11867 10935 11870
rect 12750 11868 12756 11870
rect 12820 11868 12826 11932
rect 4245 11794 4311 11797
rect 7741 11794 7807 11797
rect 10726 11794 10732 11796
rect 4245 11792 10732 11794
rect 4245 11736 4250 11792
rect 4306 11736 7746 11792
rect 7802 11736 10732 11792
rect 4245 11734 10732 11736
rect 4245 11731 4311 11734
rect 7741 11731 7807 11734
rect 10726 11732 10732 11734
rect 10796 11732 10802 11796
rect 13905 11794 13971 11797
rect 17217 11794 17283 11797
rect 22737 11794 22803 11797
rect 13905 11792 22803 11794
rect 13905 11736 13910 11792
rect 13966 11736 17222 11792
rect 17278 11736 22742 11792
rect 22798 11736 22803 11792
rect 13905 11734 22803 11736
rect 13905 11731 13971 11734
rect 17217 11731 17283 11734
rect 22737 11731 22803 11734
rect 2589 11658 2655 11661
rect 11237 11658 11303 11661
rect 2589 11656 11303 11658
rect 2589 11600 2594 11656
rect 2650 11600 11242 11656
rect 11298 11600 11303 11656
rect 2589 11598 11303 11600
rect 2589 11595 2655 11598
rect 11237 11595 11303 11598
rect 12566 11596 12572 11660
rect 12636 11658 12642 11660
rect 12801 11658 12867 11661
rect 14181 11658 14247 11661
rect 15009 11658 15075 11661
rect 12636 11656 15075 11658
rect 12636 11600 12806 11656
rect 12862 11600 14186 11656
rect 14242 11600 15014 11656
rect 15070 11600 15075 11656
rect 12636 11598 15075 11600
rect 12636 11596 12642 11598
rect 12801 11595 12867 11598
rect 14181 11595 14247 11598
rect 15009 11595 15075 11598
rect 15694 11596 15700 11660
rect 15764 11658 15770 11660
rect 17493 11658 17559 11661
rect 15764 11656 17559 11658
rect 15764 11600 17498 11656
rect 17554 11600 17559 11656
rect 15764 11598 17559 11600
rect 15764 11596 15770 11598
rect 17493 11595 17559 11598
rect 0 11520 480 11552
rect 0 11464 18 11520
rect 74 11464 480 11520
rect 0 11432 480 11464
rect 2630 11460 2636 11524
rect 2700 11522 2706 11524
rect 4889 11522 4955 11525
rect 2700 11520 4955 11522
rect 2700 11464 4894 11520
rect 4950 11464 4955 11520
rect 2700 11462 4955 11464
rect 2700 11460 2706 11462
rect 4889 11459 4955 11462
rect 5257 11522 5323 11525
rect 5390 11522 5396 11524
rect 5257 11520 5396 11522
rect 5257 11464 5262 11520
rect 5318 11464 5396 11520
rect 5257 11462 5396 11464
rect 5257 11459 5323 11462
rect 5390 11460 5396 11462
rect 5460 11522 5466 11524
rect 9581 11522 9647 11525
rect 15142 11522 15148 11524
rect 5460 11462 8540 11522
rect 5460 11460 5466 11462
rect 8480 11389 8540 11462
rect 9581 11520 15148 11522
rect 9581 11464 9586 11520
rect 9642 11464 15148 11520
rect 9581 11462 15148 11464
rect 9581 11459 9647 11462
rect 15142 11460 15148 11462
rect 15212 11460 15218 11524
rect 18822 11460 18828 11524
rect 18892 11522 18898 11524
rect 19609 11522 19675 11525
rect 18892 11520 19675 11522
rect 18892 11464 19614 11520
rect 19670 11464 19675 11520
rect 18892 11462 19675 11464
rect 18892 11460 18898 11462
rect 19609 11459 19675 11462
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 23520 11432 24000 11552
rect 16944 11391 17264 11392
rect 1526 11324 1532 11388
rect 1596 11386 1602 11388
rect 5390 11386 5396 11388
rect 1596 11326 5396 11386
rect 1596 11324 1602 11326
rect 5390 11324 5396 11326
rect 5460 11324 5466 11388
rect 7230 11324 7236 11388
rect 7300 11386 7306 11388
rect 8334 11386 8340 11388
rect 7300 11326 8340 11386
rect 7300 11324 7306 11326
rect 8334 11324 8340 11326
rect 8404 11324 8410 11388
rect 8477 11384 8543 11389
rect 16757 11386 16823 11389
rect 22001 11386 22067 11389
rect 8477 11328 8482 11384
rect 8538 11328 8543 11384
rect 8477 11323 8543 11328
rect 9630 11384 16823 11386
rect 9630 11328 16762 11384
rect 16818 11328 16823 11384
rect 9630 11326 16823 11328
rect 1526 11188 1532 11252
rect 1596 11250 1602 11252
rect 2497 11250 2563 11253
rect 1596 11248 2563 11250
rect 1596 11192 2502 11248
rect 2558 11192 2563 11248
rect 1596 11190 2563 11192
rect 1596 11188 1602 11190
rect 2497 11187 2563 11190
rect 3550 11188 3556 11252
rect 3620 11250 3626 11252
rect 9630 11250 9690 11326
rect 16757 11323 16823 11326
rect 18094 11384 22067 11386
rect 18094 11328 22006 11384
rect 22062 11328 22067 11384
rect 18094 11326 22067 11328
rect 3620 11190 9690 11250
rect 3620 11188 3626 11190
rect 11462 11188 11468 11252
rect 11532 11250 11538 11252
rect 12065 11250 12131 11253
rect 11532 11248 12131 11250
rect 11532 11192 12070 11248
rect 12126 11192 12131 11248
rect 11532 11190 12131 11192
rect 11532 11188 11538 11190
rect 12065 11187 12131 11190
rect 12382 11188 12388 11252
rect 12452 11250 12458 11252
rect 18094 11250 18154 11326
rect 22001 11323 22067 11326
rect 12452 11190 18154 11250
rect 12452 11188 12458 11190
rect 18638 11188 18644 11252
rect 18708 11250 18714 11252
rect 22277 11250 22343 11253
rect 18708 11248 22343 11250
rect 18708 11192 22282 11248
rect 22338 11192 22343 11248
rect 18708 11190 22343 11192
rect 18708 11188 18714 11190
rect 22277 11187 22343 11190
rect 1393 11114 1459 11117
rect 5717 11114 5783 11117
rect 8109 11114 8175 11117
rect 1393 11112 5783 11114
rect 1393 11056 1398 11112
rect 1454 11056 5722 11112
rect 5778 11056 5783 11112
rect 1393 11054 5783 11056
rect 1393 11051 1459 11054
rect 5717 11051 5783 11054
rect 7468 11112 8175 11114
rect 7468 11056 8114 11112
rect 8170 11056 8175 11112
rect 7468 11054 8175 11056
rect 54 10916 60 10980
rect 124 10978 130 10980
rect 1209 10978 1275 10981
rect 124 10976 1275 10978
rect 124 10920 1214 10976
rect 1270 10920 1275 10976
rect 124 10918 1275 10920
rect 124 10916 130 10918
rect 1209 10915 1275 10918
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 3969 10842 4035 10845
rect 3052 10840 4035 10842
rect 3052 10784 3974 10840
rect 4030 10784 4035 10840
rect 3052 10782 4035 10784
rect 7468 10842 7528 11054
rect 8109 11051 8175 11054
rect 11278 11052 11284 11116
rect 11348 11114 11354 11116
rect 11421 11114 11487 11117
rect 13353 11114 13419 11117
rect 11348 11112 13419 11114
rect 11348 11056 11426 11112
rect 11482 11056 13358 11112
rect 13414 11056 13419 11112
rect 11348 11054 13419 11056
rect 11348 11052 11354 11054
rect 11421 11051 11487 11054
rect 13353 11051 13419 11054
rect 13905 11114 13971 11117
rect 23614 11114 23674 11432
rect 13905 11112 23674 11114
rect 13905 11056 13910 11112
rect 13966 11056 23674 11112
rect 13905 11054 23674 11056
rect 13905 11051 13971 11054
rect 7649 10978 7715 10981
rect 10174 10978 10180 10980
rect 7649 10976 10180 10978
rect 7649 10920 7654 10976
rect 7710 10920 10180 10976
rect 7649 10918 10180 10920
rect 7649 10915 7715 10918
rect 10174 10916 10180 10918
rect 10244 10916 10250 10980
rect 13445 10978 13511 10981
rect 15142 10978 15148 10980
rect 13445 10976 15148 10978
rect 13445 10920 13450 10976
rect 13506 10920 15148 10976
rect 13445 10918 15148 10920
rect 13445 10915 13511 10918
rect 15142 10916 15148 10918
rect 15212 10978 15218 10980
rect 15285 10978 15351 10981
rect 15212 10976 15351 10978
rect 15212 10920 15290 10976
rect 15346 10920 15351 10976
rect 15212 10918 15351 10920
rect 15212 10916 15218 10918
rect 15285 10915 15351 10918
rect 22001 10978 22067 10981
rect 23606 10978 23612 10980
rect 22001 10976 23612 10978
rect 22001 10920 22006 10976
rect 22062 10920 23612 10976
rect 22001 10918 23612 10920
rect 22001 10915 22067 10918
rect 23606 10916 23612 10918
rect 23676 10916 23682 10980
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 7649 10842 7715 10845
rect 7468 10840 7715 10842
rect 7468 10784 7654 10840
rect 7710 10784 7715 10840
rect 7468 10782 7715 10784
rect 0 10708 480 10736
rect 0 10644 60 10708
rect 124 10644 480 10708
rect 0 10616 480 10644
rect 1577 10706 1643 10709
rect 2681 10706 2747 10709
rect 3052 10706 3112 10782
rect 3969 10779 4035 10782
rect 7649 10779 7715 10782
rect 8334 10780 8340 10844
rect 8404 10842 8410 10844
rect 12433 10842 12499 10845
rect 8404 10840 12499 10842
rect 8404 10784 12438 10840
rect 12494 10784 12499 10840
rect 8404 10782 12499 10784
rect 8404 10780 8410 10782
rect 12433 10779 12499 10782
rect 13445 10842 13511 10845
rect 13670 10842 13676 10844
rect 13445 10840 13676 10842
rect 13445 10784 13450 10840
rect 13506 10784 13676 10840
rect 13445 10782 13676 10784
rect 13445 10779 13511 10782
rect 13670 10780 13676 10782
rect 13740 10780 13746 10844
rect 14641 10842 14707 10845
rect 19885 10842 19951 10845
rect 14641 10840 19951 10842
rect 14641 10784 14646 10840
rect 14702 10784 19890 10840
rect 19946 10784 19951 10840
rect 14641 10782 19951 10784
rect 14641 10779 14707 10782
rect 19885 10779 19951 10782
rect 1577 10704 3112 10706
rect 1577 10648 1582 10704
rect 1638 10648 2686 10704
rect 2742 10648 3112 10704
rect 1577 10646 3112 10648
rect 1577 10643 1643 10646
rect 2681 10643 2747 10646
rect 4286 10644 4292 10708
rect 4356 10706 4362 10708
rect 4521 10706 4587 10709
rect 4356 10704 4587 10706
rect 4356 10648 4526 10704
rect 4582 10648 4587 10704
rect 4356 10646 4587 10648
rect 4356 10644 4362 10646
rect 4521 10643 4587 10646
rect 6729 10706 6795 10709
rect 10685 10706 10751 10709
rect 11329 10706 11395 10709
rect 6729 10704 11395 10706
rect 6729 10648 6734 10704
rect 6790 10648 10690 10704
rect 10746 10648 11334 10704
rect 11390 10648 11395 10704
rect 6729 10646 11395 10648
rect 6729 10643 6795 10646
rect 10685 10643 10751 10646
rect 11329 10643 11395 10646
rect 12525 10706 12591 10709
rect 12750 10706 12756 10708
rect 12525 10704 12756 10706
rect 12525 10648 12530 10704
rect 12586 10648 12756 10704
rect 12525 10646 12756 10648
rect 12525 10643 12591 10646
rect 12750 10644 12756 10646
rect 12820 10644 12826 10708
rect 12985 10706 13051 10709
rect 13997 10706 14063 10709
rect 12985 10704 14063 10706
rect 12985 10648 12990 10704
rect 13046 10648 14002 10704
rect 14058 10648 14063 10704
rect 12985 10646 14063 10648
rect 12985 10643 13051 10646
rect 13997 10643 14063 10646
rect 15561 10706 15627 10709
rect 15561 10704 23674 10706
rect 15561 10648 15566 10704
rect 15622 10648 23674 10704
rect 15561 10646 23674 10648
rect 15561 10643 15627 10646
rect 3366 10508 3372 10572
rect 3436 10570 3442 10572
rect 3969 10570 4035 10573
rect 3436 10568 4035 10570
rect 3436 10512 3974 10568
rect 4030 10512 4035 10568
rect 3436 10510 4035 10512
rect 3436 10508 3442 10510
rect 3969 10507 4035 10510
rect 4286 10508 4292 10572
rect 4356 10570 4362 10572
rect 4705 10570 4771 10573
rect 4356 10568 4771 10570
rect 4356 10512 4710 10568
rect 4766 10512 4771 10568
rect 4356 10510 4771 10512
rect 4356 10508 4362 10510
rect 4705 10507 4771 10510
rect 4889 10570 4955 10573
rect 4889 10568 7528 10570
rect 4889 10512 4894 10568
rect 4950 10512 7528 10568
rect 4889 10510 7528 10512
rect 4889 10507 4955 10510
rect 1710 10372 1716 10436
rect 1780 10434 1786 10436
rect 5901 10434 5967 10437
rect 1780 10432 5967 10434
rect 1780 10376 5906 10432
rect 5962 10376 5967 10432
rect 1780 10374 5967 10376
rect 1780 10372 1786 10374
rect 5901 10371 5967 10374
rect 6729 10434 6795 10437
rect 7230 10434 7236 10436
rect 6729 10432 7236 10434
rect 6729 10376 6734 10432
rect 6790 10376 7236 10432
rect 6729 10374 7236 10376
rect 6729 10371 6795 10374
rect 7230 10372 7236 10374
rect 7300 10372 7306 10436
rect 7468 10434 7528 10510
rect 7598 10508 7604 10572
rect 7668 10570 7674 10572
rect 8109 10570 8175 10573
rect 7668 10568 8175 10570
rect 7668 10512 8114 10568
rect 8170 10512 8175 10568
rect 7668 10510 8175 10512
rect 7668 10508 7674 10510
rect 8109 10507 8175 10510
rect 9949 10570 10015 10573
rect 11329 10570 11395 10573
rect 16941 10570 17007 10573
rect 9949 10568 17007 10570
rect 9949 10512 9954 10568
rect 10010 10512 11334 10568
rect 11390 10512 16946 10568
rect 17002 10512 17007 10568
rect 9949 10510 17007 10512
rect 9949 10507 10015 10510
rect 11329 10507 11395 10510
rect 16941 10507 17007 10510
rect 18638 10508 18644 10572
rect 18708 10570 18714 10572
rect 21909 10570 21975 10573
rect 18708 10568 21975 10570
rect 18708 10512 21914 10568
rect 21970 10512 21975 10568
rect 18708 10510 21975 10512
rect 18708 10508 18714 10510
rect 21909 10507 21975 10510
rect 23614 10464 23674 10646
rect 8753 10434 8819 10437
rect 7468 10432 8819 10434
rect 7468 10376 8758 10432
rect 8814 10376 8819 10432
rect 7468 10374 8819 10376
rect 8753 10371 8819 10374
rect 10041 10434 10107 10437
rect 11278 10434 11284 10436
rect 10041 10432 11284 10434
rect 10041 10376 10046 10432
rect 10102 10376 11284 10432
rect 10041 10374 11284 10376
rect 10041 10371 10107 10374
rect 11278 10372 11284 10374
rect 11348 10434 11354 10436
rect 15285 10434 15351 10437
rect 11348 10432 15351 10434
rect 11348 10376 15290 10432
rect 15346 10376 15351 10432
rect 11348 10374 15351 10376
rect 11348 10372 11354 10374
rect 15285 10371 15351 10374
rect 19558 10372 19564 10436
rect 19628 10434 19634 10436
rect 20437 10434 20503 10437
rect 19628 10432 20503 10434
rect 19628 10376 20442 10432
rect 20498 10376 20503 10432
rect 19628 10374 20503 10376
rect 19628 10372 19634 10374
rect 20437 10371 20503 10374
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 23520 10344 24000 10464
rect 16944 10303 17264 10304
rect 1710 10236 1716 10300
rect 1780 10298 1786 10300
rect 2681 10298 2747 10301
rect 1780 10296 2747 10298
rect 1780 10240 2686 10296
rect 2742 10240 2747 10296
rect 1780 10238 2747 10240
rect 1780 10236 1786 10238
rect 2681 10235 2747 10238
rect 4102 10236 4108 10300
rect 4172 10298 4178 10300
rect 4337 10298 4403 10301
rect 7230 10298 7236 10300
rect 4172 10296 4403 10298
rect 4172 10240 4342 10296
rect 4398 10240 4403 10296
rect 4172 10238 4403 10240
rect 4172 10236 4178 10238
rect 4337 10235 4403 10238
rect 4478 10238 7236 10298
rect 2865 10162 2931 10165
rect 4478 10162 4538 10238
rect 7230 10236 7236 10238
rect 7300 10298 7306 10300
rect 8569 10298 8635 10301
rect 7300 10296 8635 10298
rect 7300 10240 8574 10296
rect 8630 10240 8635 10296
rect 7300 10238 8635 10240
rect 7300 10236 7306 10238
rect 8569 10235 8635 10238
rect 12566 10236 12572 10300
rect 12636 10298 12642 10300
rect 13353 10298 13419 10301
rect 12636 10296 13419 10298
rect 12636 10240 13358 10296
rect 13414 10240 13419 10296
rect 12636 10238 13419 10240
rect 12636 10236 12642 10238
rect 13353 10235 13419 10238
rect 13997 10298 14063 10301
rect 14222 10298 14228 10300
rect 13997 10296 14228 10298
rect 13997 10240 14002 10296
rect 14058 10240 14228 10296
rect 13997 10238 14228 10240
rect 13997 10235 14063 10238
rect 14222 10236 14228 10238
rect 14292 10236 14298 10300
rect 17401 10298 17467 10301
rect 17718 10298 17724 10300
rect 17401 10296 17724 10298
rect 17401 10240 17406 10296
rect 17462 10240 17724 10296
rect 17401 10238 17724 10240
rect 17401 10235 17467 10238
rect 17718 10236 17724 10238
rect 17788 10236 17794 10300
rect 21950 10236 21956 10300
rect 22020 10298 22026 10300
rect 22369 10298 22435 10301
rect 22020 10296 22435 10298
rect 22020 10240 22374 10296
rect 22430 10240 22435 10296
rect 22020 10238 22435 10240
rect 22020 10236 22026 10238
rect 22369 10235 22435 10238
rect 2865 10160 4538 10162
rect 2865 10104 2870 10160
rect 2926 10104 4538 10160
rect 2865 10102 4538 10104
rect 4705 10162 4771 10165
rect 6085 10162 6151 10165
rect 4705 10160 6151 10162
rect 4705 10104 4710 10160
rect 4766 10104 6090 10160
rect 6146 10104 6151 10160
rect 4705 10102 6151 10104
rect 2865 10099 2931 10102
rect 4705 10099 4771 10102
rect 6085 10099 6151 10102
rect 6637 10160 6703 10165
rect 6637 10104 6642 10160
rect 6698 10104 6703 10160
rect 6637 10099 6703 10104
rect 7833 10162 7899 10165
rect 11697 10162 11763 10165
rect 12893 10162 12959 10165
rect 7833 10160 12959 10162
rect 7833 10104 7838 10160
rect 7894 10104 11702 10160
rect 11758 10104 12898 10160
rect 12954 10104 12959 10160
rect 7833 10102 12959 10104
rect 7833 10099 7899 10102
rect 11697 10099 11763 10102
rect 12893 10099 12959 10102
rect 13353 10162 13419 10165
rect 15009 10162 15075 10165
rect 13353 10160 15075 10162
rect 13353 10104 13358 10160
rect 13414 10104 15014 10160
rect 15070 10104 15075 10160
rect 13353 10102 15075 10104
rect 13353 10099 13419 10102
rect 15009 10099 15075 10102
rect 15326 10100 15332 10164
rect 15396 10162 15402 10164
rect 17125 10162 17191 10165
rect 15396 10160 17191 10162
rect 15396 10104 17130 10160
rect 17186 10104 17191 10160
rect 15396 10102 17191 10104
rect 15396 10100 15402 10102
rect 17125 10099 17191 10102
rect 62 9966 3940 10026
rect 62 9920 122 9966
rect 0 9800 480 9920
rect 565 9890 631 9893
rect 2129 9890 2195 9893
rect 3734 9890 3740 9892
rect 565 9888 3740 9890
rect 565 9832 570 9888
rect 626 9832 2134 9888
rect 2190 9832 3740 9888
rect 565 9830 3740 9832
rect 565 9827 631 9830
rect 2129 9827 2195 9830
rect 3734 9828 3740 9830
rect 3804 9828 3810 9892
rect 3880 9890 3940 9966
rect 4286 9964 4292 10028
rect 4356 10026 4362 10028
rect 4889 10026 4955 10029
rect 4356 10024 4955 10026
rect 4356 9968 4894 10024
rect 4950 9968 4955 10024
rect 4356 9966 4955 9968
rect 6640 10028 6700 10099
rect 6640 9966 6684 10028
rect 4356 9964 4362 9966
rect 4889 9963 4955 9966
rect 6678 9964 6684 9966
rect 6748 9964 6754 10028
rect 8334 9964 8340 10028
rect 8404 10026 8410 10028
rect 11094 10026 11100 10028
rect 8404 9966 11100 10026
rect 8404 9964 8410 9966
rect 11094 9964 11100 9966
rect 11164 9964 11170 10028
rect 11646 9964 11652 10028
rect 11716 10026 11722 10028
rect 12617 10026 12683 10029
rect 14365 10026 14431 10029
rect 14733 10026 14799 10029
rect 16941 10026 17007 10029
rect 11716 10024 12683 10026
rect 11716 9968 12622 10024
rect 12678 9968 12683 10024
rect 11716 9966 12683 9968
rect 11716 9964 11722 9966
rect 12617 9963 12683 9966
rect 12804 10024 14431 10026
rect 12804 9968 14370 10024
rect 14426 9968 14431 10024
rect 12804 9966 14431 9968
rect 14606 10024 17007 10026
rect 14606 9968 14738 10024
rect 14794 9968 16946 10024
rect 17002 9968 17007 10024
rect 14606 9966 17007 9968
rect 4153 9890 4219 9893
rect 4429 9890 4495 9893
rect 3880 9888 4219 9890
rect 3880 9832 4158 9888
rect 4214 9832 4219 9888
rect 3880 9830 4219 9832
rect 4153 9827 4219 9830
rect 4294 9888 4495 9890
rect 4294 9832 4434 9888
rect 4490 9832 4495 9888
rect 4294 9830 4495 9832
rect 2129 9754 2195 9757
rect 2957 9754 3023 9757
rect 2129 9752 3023 9754
rect 2129 9696 2134 9752
rect 2190 9696 2962 9752
rect 3018 9696 3023 9752
rect 2129 9694 3023 9696
rect 2129 9691 2195 9694
rect 2957 9691 3023 9694
rect 3734 9692 3740 9756
rect 3804 9754 3810 9756
rect 4294 9754 4354 9830
rect 4429 9827 4495 9830
rect 4613 9888 4679 9893
rect 4613 9832 4618 9888
rect 4674 9832 4679 9888
rect 4613 9827 4679 9832
rect 5717 9890 5783 9893
rect 8569 9890 8635 9893
rect 5717 9888 8635 9890
rect 5717 9832 5722 9888
rect 5778 9832 8574 9888
rect 8630 9832 8635 9888
rect 5717 9830 8635 9832
rect 5717 9827 5783 9830
rect 8569 9827 8635 9830
rect 8702 9828 8708 9892
rect 8772 9890 8778 9892
rect 9438 9890 9444 9892
rect 8772 9830 9444 9890
rect 8772 9828 8778 9830
rect 9438 9828 9444 9830
rect 9508 9828 9514 9892
rect 10910 9828 10916 9892
rect 10980 9890 10986 9892
rect 11462 9890 11468 9892
rect 10980 9830 11468 9890
rect 10980 9828 10986 9830
rect 11462 9828 11468 9830
rect 11532 9828 11538 9892
rect 12249 9890 12315 9893
rect 12804 9890 12864 9966
rect 14365 9963 14431 9966
rect 14733 9963 14799 9966
rect 16941 9963 17007 9966
rect 18413 10026 18479 10029
rect 19977 10026 20043 10029
rect 18413 10024 20043 10026
rect 18413 9968 18418 10024
rect 18474 9968 19982 10024
rect 20038 9968 20043 10024
rect 18413 9966 20043 9968
rect 18413 9963 18479 9966
rect 19977 9963 20043 9966
rect 20294 9964 20300 10028
rect 20364 10026 20370 10028
rect 21449 10026 21515 10029
rect 20364 10024 21515 10026
rect 20364 9968 21454 10024
rect 21510 9968 21515 10024
rect 20364 9966 21515 9968
rect 20364 9964 20370 9966
rect 21449 9963 21515 9966
rect 20621 9890 20687 9893
rect 12249 9888 12864 9890
rect 12249 9832 12254 9888
rect 12310 9832 12864 9888
rect 12249 9830 12864 9832
rect 13356 9888 20687 9890
rect 13356 9832 20626 9888
rect 20682 9832 20687 9888
rect 13356 9830 20687 9832
rect 12249 9827 12315 9830
rect 4616 9754 4676 9827
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 3804 9694 4354 9754
rect 4432 9694 4676 9754
rect 3804 9692 3810 9694
rect 2589 9482 2655 9485
rect 62 9480 2655 9482
rect 62 9424 2594 9480
rect 2650 9424 2655 9480
rect 62 9422 2655 9424
rect 62 9104 122 9422
rect 2589 9419 2655 9422
rect 3233 9482 3299 9485
rect 3366 9482 3372 9484
rect 3233 9480 3372 9482
rect 3233 9424 3238 9480
rect 3294 9424 3372 9480
rect 3233 9422 3372 9424
rect 3233 9419 3299 9422
rect 3366 9420 3372 9422
rect 3436 9420 3442 9484
rect 4153 9482 4219 9485
rect 4432 9482 4492 9694
rect 5390 9692 5396 9756
rect 5460 9754 5466 9756
rect 5809 9754 5875 9757
rect 5460 9752 5875 9754
rect 5460 9696 5814 9752
rect 5870 9696 5875 9752
rect 5460 9694 5875 9696
rect 5460 9692 5466 9694
rect 5809 9691 5875 9694
rect 6085 9754 6151 9757
rect 7598 9754 7604 9756
rect 6085 9752 7604 9754
rect 6085 9696 6090 9752
rect 6146 9696 7604 9752
rect 6085 9694 7604 9696
rect 6085 9691 6151 9694
rect 7598 9692 7604 9694
rect 7668 9692 7674 9756
rect 8201 9754 8267 9757
rect 9622 9754 9628 9756
rect 8201 9752 9628 9754
rect 8201 9696 8206 9752
rect 8262 9696 9628 9752
rect 8201 9694 9628 9696
rect 8201 9691 8267 9694
rect 9622 9692 9628 9694
rect 9692 9692 9698 9756
rect 4654 9556 4660 9620
rect 4724 9618 4730 9620
rect 4981 9618 5047 9621
rect 4724 9616 5047 9618
rect 4724 9560 4986 9616
rect 5042 9560 5047 9616
rect 4724 9558 5047 9560
rect 4724 9556 4730 9558
rect 4981 9555 5047 9558
rect 5165 9618 5231 9621
rect 8702 9618 8708 9620
rect 5165 9616 8708 9618
rect 5165 9560 5170 9616
rect 5226 9560 8708 9616
rect 5165 9558 8708 9560
rect 5165 9555 5231 9558
rect 8702 9556 8708 9558
rect 8772 9556 8778 9620
rect 13356 9618 13416 9830
rect 20621 9827 20687 9830
rect 21582 9828 21588 9892
rect 21652 9890 21658 9892
rect 22277 9890 22343 9893
rect 21652 9888 22343 9890
rect 21652 9832 22282 9888
rect 22338 9832 22343 9888
rect 21652 9830 22343 9832
rect 21652 9828 21658 9830
rect 22277 9827 22343 9830
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 13537 9754 13603 9757
rect 14406 9754 14412 9756
rect 13537 9752 14412 9754
rect 13537 9696 13542 9752
rect 13598 9696 14412 9752
rect 13537 9694 14412 9696
rect 13537 9691 13603 9694
rect 14406 9692 14412 9694
rect 14476 9692 14482 9756
rect 18321 9754 18387 9757
rect 20294 9754 20300 9756
rect 18321 9752 20300 9754
rect 18321 9696 18326 9752
rect 18382 9696 20300 9752
rect 18321 9694 20300 9696
rect 18321 9691 18387 9694
rect 20294 9692 20300 9694
rect 20364 9692 20370 9756
rect 11056 9558 13416 9618
rect 11056 9485 11116 9558
rect 4153 9480 4492 9482
rect 4153 9424 4158 9480
rect 4214 9424 4492 9480
rect 4153 9422 4492 9424
rect 4889 9482 4955 9485
rect 7833 9482 7899 9485
rect 4889 9480 7899 9482
rect 4889 9424 4894 9480
rect 4950 9424 7838 9480
rect 7894 9424 7899 9480
rect 4889 9422 7899 9424
rect 4153 9419 4219 9422
rect 4889 9419 4955 9422
rect 7833 9419 7899 9422
rect 10910 9420 10916 9484
rect 10980 9482 10986 9484
rect 11053 9482 11119 9485
rect 10980 9480 11119 9482
rect 10980 9424 11058 9480
rect 11114 9424 11119 9480
rect 10980 9422 11119 9424
rect 10980 9420 10986 9422
rect 11053 9419 11119 9422
rect 11881 9482 11947 9485
rect 12249 9482 12315 9485
rect 11881 9480 12315 9482
rect 11881 9424 11886 9480
rect 11942 9424 12254 9480
rect 12310 9424 12315 9480
rect 11881 9422 12315 9424
rect 11881 9419 11947 9422
rect 12249 9419 12315 9422
rect 15009 9482 15075 9485
rect 21081 9482 21147 9485
rect 15009 9480 21147 9482
rect 15009 9424 15014 9480
rect 15070 9424 21086 9480
rect 21142 9424 21147 9480
rect 15009 9422 21147 9424
rect 15009 9419 15075 9422
rect 21081 9419 21147 9422
rect 1485 9346 1551 9349
rect 8753 9346 8819 9349
rect 1485 9344 8819 9346
rect 1485 9288 1490 9344
rect 1546 9288 8758 9344
rect 8814 9288 8819 9344
rect 1485 9286 8819 9288
rect 1485 9283 1551 9286
rect 8753 9283 8819 9286
rect 12198 9284 12204 9348
rect 12268 9346 12274 9348
rect 13813 9346 13879 9349
rect 12268 9344 13879 9346
rect 12268 9288 13818 9344
rect 13874 9288 13879 9344
rect 12268 9286 13879 9288
rect 12268 9284 12274 9286
rect 13813 9283 13879 9286
rect 22001 9346 22067 9349
rect 23520 9346 24000 9376
rect 22001 9344 24000 9346
rect 22001 9288 22006 9344
rect 22062 9288 24000 9344
rect 22001 9286 24000 9288
rect 22001 9283 22067 9286
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 23520 9256 24000 9286
rect 16944 9215 17264 9216
rect 974 9148 980 9212
rect 1044 9210 1050 9212
rect 1209 9210 1275 9213
rect 1044 9208 1275 9210
rect 1044 9152 1214 9208
rect 1270 9152 1275 9208
rect 1044 9150 1275 9152
rect 1044 9148 1050 9150
rect 1209 9147 1275 9150
rect 1894 9148 1900 9212
rect 1964 9210 1970 9212
rect 2037 9210 2103 9213
rect 1964 9208 2103 9210
rect 1964 9152 2042 9208
rect 2098 9152 2103 9208
rect 1964 9150 2103 9152
rect 1964 9148 1970 9150
rect 2037 9147 2103 9150
rect 3417 9210 3483 9213
rect 3734 9210 3740 9212
rect 3417 9208 3740 9210
rect 3417 9152 3422 9208
rect 3478 9152 3740 9208
rect 3417 9150 3740 9152
rect 3417 9147 3483 9150
rect 3734 9148 3740 9150
rect 3804 9148 3810 9212
rect 4429 9210 4495 9213
rect 4654 9210 4660 9212
rect 4429 9208 4660 9210
rect 4429 9152 4434 9208
rect 4490 9152 4660 9208
rect 4429 9150 4660 9152
rect 4429 9147 4495 9150
rect 4654 9148 4660 9150
rect 4724 9148 4730 9212
rect 4981 9210 5047 9213
rect 5390 9210 5396 9212
rect 4981 9208 5396 9210
rect 4981 9152 4986 9208
rect 5042 9152 5396 9208
rect 4981 9150 5396 9152
rect 4981 9147 5047 9150
rect 5390 9148 5396 9150
rect 5460 9148 5466 9212
rect 8753 9210 8819 9213
rect 5536 9208 8819 9210
rect 5536 9152 8758 9208
rect 8814 9152 8819 9208
rect 5536 9150 8819 9152
rect 0 8984 480 9104
rect 3049 9074 3115 9077
rect 5257 9074 5323 9077
rect 5536 9076 5596 9150
rect 8753 9147 8819 9150
rect 11646 9148 11652 9212
rect 11716 9210 11722 9212
rect 12157 9210 12223 9213
rect 11716 9208 12223 9210
rect 11716 9152 12162 9208
rect 12218 9152 12223 9208
rect 11716 9150 12223 9152
rect 11716 9148 11722 9150
rect 12157 9147 12223 9150
rect 18045 9210 18111 9213
rect 18270 9210 18276 9212
rect 18045 9208 18276 9210
rect 18045 9152 18050 9208
rect 18106 9152 18276 9208
rect 18045 9150 18276 9152
rect 18045 9147 18111 9150
rect 18270 9148 18276 9150
rect 18340 9148 18346 9212
rect 19374 9148 19380 9212
rect 19444 9210 19450 9212
rect 20161 9210 20227 9213
rect 19444 9208 20227 9210
rect 19444 9152 20166 9208
rect 20222 9152 20227 9208
rect 19444 9150 20227 9152
rect 19444 9148 19450 9150
rect 20161 9147 20227 9150
rect 5536 9074 5580 9076
rect 3049 9072 5323 9074
rect 3049 9016 3054 9072
rect 3110 9016 5262 9072
rect 5318 9016 5323 9072
rect 3049 9014 5323 9016
rect 3049 9011 3115 9014
rect 5257 9011 5323 9014
rect 5398 9014 5580 9074
rect 1209 8938 1275 8941
rect 1526 8938 1532 8940
rect 1209 8936 1532 8938
rect 1209 8880 1214 8936
rect 1270 8880 1532 8936
rect 1209 8878 1532 8880
rect 1209 8875 1275 8878
rect 1526 8876 1532 8878
rect 1596 8876 1602 8940
rect 3233 8938 3299 8941
rect 3734 8938 3740 8940
rect 3233 8936 3740 8938
rect 3233 8880 3238 8936
rect 3294 8880 3740 8936
rect 3233 8878 3740 8880
rect 3233 8875 3299 8878
rect 3734 8876 3740 8878
rect 3804 8938 3810 8940
rect 5398 8938 5458 9014
rect 5574 9012 5580 9014
rect 5644 9074 5650 9076
rect 7465 9074 7531 9077
rect 5644 9072 7531 9074
rect 5644 9016 7470 9072
rect 7526 9016 7531 9072
rect 5644 9014 7531 9016
rect 5644 9012 5650 9014
rect 7465 9011 7531 9014
rect 9765 9074 9831 9077
rect 10358 9074 10364 9076
rect 9765 9072 10364 9074
rect 9765 9016 9770 9072
rect 9826 9016 10364 9072
rect 9765 9014 10364 9016
rect 9765 9011 9831 9014
rect 10358 9012 10364 9014
rect 10428 9012 10434 9076
rect 14089 9074 14155 9077
rect 11470 9072 14155 9074
rect 11470 9016 14094 9072
rect 14150 9016 14155 9072
rect 11470 9014 14155 9016
rect 3804 8878 5458 8938
rect 5993 8938 6059 8941
rect 7046 8938 7052 8940
rect 5993 8936 7052 8938
rect 5993 8880 5998 8936
rect 6054 8880 7052 8936
rect 5993 8878 7052 8880
rect 3804 8876 3810 8878
rect 5993 8875 6059 8878
rect 7046 8876 7052 8878
rect 7116 8938 7122 8940
rect 7557 8938 7623 8941
rect 7116 8936 7623 8938
rect 7116 8880 7562 8936
rect 7618 8880 7623 8936
rect 7116 8878 7623 8880
rect 7116 8876 7122 8878
rect 7557 8875 7623 8878
rect 7782 8876 7788 8940
rect 7852 8938 7858 8940
rect 8702 8938 8708 8940
rect 7852 8878 8708 8938
rect 7852 8876 7858 8878
rect 8702 8876 8708 8878
rect 8772 8876 8778 8940
rect 8845 8938 8911 8941
rect 10358 8938 10364 8940
rect 8845 8936 10364 8938
rect 8845 8880 8850 8936
rect 8906 8880 10364 8936
rect 8845 8878 10364 8880
rect 8845 8875 8911 8878
rect 10358 8876 10364 8878
rect 10428 8938 10434 8940
rect 11470 8938 11530 9014
rect 14089 9011 14155 9014
rect 16665 9074 16731 9077
rect 17217 9074 17283 9077
rect 16665 9072 17283 9074
rect 16665 9016 16670 9072
rect 16726 9016 17222 9072
rect 17278 9016 17283 9072
rect 16665 9014 17283 9016
rect 16665 9011 16731 9014
rect 17217 9011 17283 9014
rect 19926 9012 19932 9076
rect 19996 9074 20002 9076
rect 21725 9074 21791 9077
rect 19996 9072 21791 9074
rect 19996 9016 21730 9072
rect 21786 9016 21791 9072
rect 19996 9014 21791 9016
rect 19996 9012 20002 9014
rect 21725 9011 21791 9014
rect 10428 8878 11530 8938
rect 11605 8938 11671 8941
rect 12198 8938 12204 8940
rect 11605 8936 12204 8938
rect 11605 8880 11610 8936
rect 11666 8880 12204 8936
rect 11605 8878 12204 8880
rect 10428 8876 10434 8878
rect 11605 8875 11671 8878
rect 12198 8876 12204 8878
rect 12268 8876 12274 8940
rect 13670 8938 13676 8940
rect 12758 8878 13676 8938
rect 1761 8802 1827 8805
rect 2078 8802 2084 8804
rect 1761 8800 2084 8802
rect 1761 8744 1766 8800
rect 1822 8744 2084 8800
rect 1761 8742 2084 8744
rect 1761 8739 1827 8742
rect 2078 8740 2084 8742
rect 2148 8740 2154 8804
rect 2998 8740 3004 8804
rect 3068 8802 3074 8804
rect 3877 8802 3943 8805
rect 3068 8800 3943 8802
rect 3068 8744 3882 8800
rect 3938 8744 3943 8800
rect 3068 8742 3943 8744
rect 3068 8740 3074 8742
rect 3877 8739 3943 8742
rect 4102 8740 4108 8804
rect 4172 8802 4178 8804
rect 4245 8802 4311 8805
rect 4172 8800 4311 8802
rect 4172 8744 4250 8800
rect 4306 8744 4311 8800
rect 4172 8742 4311 8744
rect 4172 8740 4178 8742
rect 4245 8739 4311 8742
rect 6269 8802 6335 8805
rect 8293 8802 8359 8805
rect 6269 8800 8359 8802
rect 6269 8744 6274 8800
rect 6330 8744 8298 8800
rect 8354 8744 8359 8800
rect 6269 8742 8359 8744
rect 6269 8739 6335 8742
rect 8293 8739 8359 8742
rect 8569 8802 8635 8805
rect 10685 8802 10751 8805
rect 11278 8802 11284 8804
rect 8569 8800 11284 8802
rect 8569 8744 8574 8800
rect 8630 8744 10690 8800
rect 10746 8744 11284 8800
rect 8569 8742 11284 8744
rect 8569 8739 8635 8742
rect 10685 8739 10751 8742
rect 11278 8740 11284 8742
rect 11348 8740 11354 8804
rect 11605 8802 11671 8805
rect 11881 8802 11947 8805
rect 11605 8800 11947 8802
rect 11605 8744 11610 8800
rect 11666 8744 11886 8800
rect 11942 8744 11947 8800
rect 11605 8742 11947 8744
rect 11605 8739 11671 8742
rect 11881 8739 11947 8742
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 2129 8666 2195 8669
rect 3550 8666 3556 8668
rect 2129 8664 3556 8666
rect 2129 8608 2134 8664
rect 2190 8608 3556 8664
rect 2129 8606 3556 8608
rect 2129 8603 2195 8606
rect 3550 8604 3556 8606
rect 3620 8604 3626 8668
rect 3693 8666 3759 8669
rect 4429 8666 4495 8669
rect 12758 8666 12818 8878
rect 13670 8876 13676 8878
rect 13740 8876 13746 8940
rect 13997 8938 14063 8941
rect 14406 8938 14412 8940
rect 13997 8936 14412 8938
rect 13997 8880 14002 8936
rect 14058 8880 14412 8936
rect 13997 8878 14412 8880
rect 13997 8875 14063 8878
rect 14406 8876 14412 8878
rect 14476 8876 14482 8940
rect 16246 8876 16252 8940
rect 16316 8938 16322 8940
rect 16665 8938 16731 8941
rect 16316 8936 16731 8938
rect 16316 8880 16670 8936
rect 16726 8880 16731 8936
rect 16316 8878 16731 8880
rect 16316 8876 16322 8878
rect 16665 8875 16731 8878
rect 19558 8876 19564 8940
rect 19628 8938 19634 8940
rect 21265 8938 21331 8941
rect 19628 8936 21331 8938
rect 19628 8880 21270 8936
rect 21326 8880 21331 8936
rect 19628 8878 21331 8880
rect 19628 8876 19634 8878
rect 21265 8875 21331 8878
rect 14089 8802 14155 8805
rect 19425 8802 19491 8805
rect 14089 8800 19491 8802
rect 14089 8744 14094 8800
rect 14150 8744 19430 8800
rect 19486 8744 19491 8800
rect 14089 8742 19491 8744
rect 14089 8739 14155 8742
rect 19425 8739 19491 8742
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 3693 8664 4495 8666
rect 3693 8608 3698 8664
rect 3754 8608 4434 8664
rect 4490 8608 4495 8664
rect 3693 8606 4495 8608
rect 3693 8603 3759 8606
rect 4429 8603 4495 8606
rect 8296 8606 12818 8666
rect 1945 8530 2011 8533
rect 7833 8530 7899 8533
rect 1945 8528 7899 8530
rect 1945 8472 1950 8528
rect 2006 8472 7838 8528
rect 7894 8472 7899 8528
rect 1945 8470 7899 8472
rect 1945 8467 2011 8470
rect 7833 8467 7899 8470
rect 1117 8394 1183 8397
rect 2262 8394 2268 8396
rect 1117 8392 2268 8394
rect 1117 8336 1122 8392
rect 1178 8336 2268 8392
rect 1117 8334 2268 8336
rect 1117 8331 1183 8334
rect 2262 8332 2268 8334
rect 2332 8332 2338 8396
rect 2589 8394 2655 8397
rect 8017 8394 8083 8397
rect 2589 8392 8083 8394
rect 2589 8336 2594 8392
rect 2650 8336 8022 8392
rect 8078 8336 8083 8392
rect 2589 8334 8083 8336
rect 2589 8331 2655 8334
rect 8017 8331 8083 8334
rect 0 8168 480 8288
rect 2681 8258 2747 8261
rect 2998 8258 3004 8260
rect 2681 8256 3004 8258
rect 2681 8200 2686 8256
rect 2742 8200 3004 8256
rect 2681 8198 3004 8200
rect 2681 8195 2747 8198
rect 2998 8196 3004 8198
rect 3068 8196 3074 8260
rect 3233 8258 3299 8261
rect 4245 8258 4311 8261
rect 3233 8256 4311 8258
rect 3233 8200 3238 8256
rect 3294 8200 4250 8256
rect 4306 8200 4311 8256
rect 3233 8198 4311 8200
rect 3233 8195 3299 8198
rect 4245 8195 4311 8198
rect 4654 8196 4660 8260
rect 4724 8258 4730 8260
rect 7833 8258 7899 8261
rect 4724 8256 7899 8258
rect 4724 8200 7838 8256
rect 7894 8200 7899 8256
rect 4724 8198 7899 8200
rect 4724 8196 4730 8198
rect 7833 8195 7899 8198
rect 62 7714 122 8168
rect 1393 8122 1459 8125
rect 2497 8122 2563 8125
rect 1393 8120 2563 8122
rect 1393 8064 1398 8120
rect 1454 8064 2502 8120
rect 2558 8064 2563 8120
rect 1393 8062 2563 8064
rect 1393 8059 1459 8062
rect 2132 7853 2192 8062
rect 2497 8059 2563 8062
rect 3693 8122 3759 8125
rect 8296 8122 8356 8606
rect 8477 8530 8543 8533
rect 13721 8530 13787 8533
rect 8477 8528 13787 8530
rect 8477 8472 8482 8528
rect 8538 8472 13726 8528
rect 13782 8472 13787 8528
rect 8477 8470 13787 8472
rect 8477 8467 8543 8470
rect 13721 8467 13787 8470
rect 13854 8468 13860 8532
rect 13924 8530 13930 8532
rect 22001 8530 22067 8533
rect 13924 8528 22067 8530
rect 13924 8472 22006 8528
rect 22062 8472 22067 8528
rect 13924 8470 22067 8472
rect 13924 8468 13930 8470
rect 22001 8467 22067 8470
rect 8753 8392 8819 8397
rect 8753 8336 8758 8392
rect 8814 8336 8819 8392
rect 8753 8331 8819 8336
rect 9765 8394 9831 8397
rect 10542 8394 10548 8396
rect 9765 8392 10548 8394
rect 9765 8336 9770 8392
rect 9826 8336 10548 8392
rect 9765 8334 10548 8336
rect 9765 8331 9831 8334
rect 10542 8332 10548 8334
rect 10612 8332 10618 8396
rect 11329 8394 11395 8397
rect 13077 8394 13143 8397
rect 11329 8392 13143 8394
rect 11329 8336 11334 8392
rect 11390 8336 13082 8392
rect 13138 8336 13143 8392
rect 11329 8334 13143 8336
rect 11329 8331 11395 8334
rect 13077 8331 13143 8334
rect 8477 8258 8543 8261
rect 8756 8258 8816 8331
rect 8477 8256 8816 8258
rect 8477 8200 8482 8256
rect 8538 8200 8816 8256
rect 8477 8198 8816 8200
rect 8477 8195 8543 8198
rect 11830 8196 11836 8260
rect 11900 8258 11906 8260
rect 13353 8258 13419 8261
rect 14457 8258 14523 8261
rect 11900 8256 14523 8258
rect 11900 8200 13358 8256
rect 13414 8200 14462 8256
rect 14518 8200 14523 8256
rect 11900 8198 14523 8200
rect 11900 8196 11906 8198
rect 13353 8195 13419 8198
rect 14457 8195 14523 8198
rect 20437 8258 20503 8261
rect 23520 8258 24000 8288
rect 20437 8256 24000 8258
rect 20437 8200 20442 8256
rect 20498 8200 24000 8256
rect 20437 8198 24000 8200
rect 20437 8195 20503 8198
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 23520 8168 24000 8198
rect 16944 8127 17264 8128
rect 3693 8120 8356 8122
rect 3693 8064 3698 8120
rect 3754 8064 8356 8120
rect 3693 8062 8356 8064
rect 3693 8059 3759 8062
rect 10358 8060 10364 8124
rect 10428 8122 10434 8124
rect 10777 8122 10843 8125
rect 10428 8120 10843 8122
rect 10428 8064 10782 8120
rect 10838 8064 10843 8120
rect 10428 8062 10843 8064
rect 10428 8060 10434 8062
rect 10777 8059 10843 8062
rect 11462 8060 11468 8124
rect 11532 8122 11538 8124
rect 11830 8122 11836 8124
rect 11532 8062 11836 8122
rect 11532 8060 11538 8062
rect 11830 8060 11836 8062
rect 11900 8122 11906 8124
rect 14089 8122 14155 8125
rect 11900 8120 14155 8122
rect 11900 8064 14094 8120
rect 14150 8064 14155 8120
rect 11900 8062 14155 8064
rect 11900 8060 11906 8062
rect 14089 8059 14155 8062
rect 2957 7986 3023 7989
rect 6177 7986 6243 7989
rect 2957 7984 6243 7986
rect 2957 7928 2962 7984
rect 3018 7928 6182 7984
rect 6238 7928 6243 7984
rect 2957 7926 6243 7928
rect 2957 7923 3023 7926
rect 6177 7923 6243 7926
rect 7097 7986 7163 7989
rect 20713 7986 20779 7989
rect 7097 7984 20779 7986
rect 7097 7928 7102 7984
rect 7158 7928 20718 7984
rect 20774 7928 20779 7984
rect 7097 7926 20779 7928
rect 7097 7923 7163 7926
rect 20713 7923 20779 7926
rect 2129 7848 2195 7853
rect 2129 7792 2134 7848
rect 2190 7792 2195 7848
rect 2129 7787 2195 7792
rect 3550 7788 3556 7852
rect 3620 7850 3626 7852
rect 5349 7850 5415 7853
rect 3620 7848 5415 7850
rect 3620 7792 5354 7848
rect 5410 7792 5415 7848
rect 3620 7790 5415 7792
rect 3620 7788 3626 7790
rect 5349 7787 5415 7790
rect 5625 7850 5691 7853
rect 5758 7850 5764 7852
rect 5625 7848 5764 7850
rect 5625 7792 5630 7848
rect 5686 7792 5764 7848
rect 5625 7790 5764 7792
rect 5625 7787 5691 7790
rect 5758 7788 5764 7790
rect 5828 7788 5834 7852
rect 6545 7850 6611 7853
rect 6678 7850 6684 7852
rect 6545 7848 6684 7850
rect 6545 7792 6550 7848
rect 6606 7792 6684 7848
rect 6545 7790 6684 7792
rect 6545 7787 6611 7790
rect 6678 7788 6684 7790
rect 6748 7788 6754 7852
rect 6862 7788 6868 7852
rect 6932 7850 6938 7852
rect 12157 7850 12223 7853
rect 15561 7850 15627 7853
rect 21633 7850 21699 7853
rect 6932 7848 12223 7850
rect 6932 7792 12162 7848
rect 12218 7792 12223 7848
rect 6932 7790 12223 7792
rect 6932 7788 6938 7790
rect 12157 7787 12223 7790
rect 12758 7848 15627 7850
rect 12758 7792 15566 7848
rect 15622 7792 15627 7848
rect 12758 7790 15627 7792
rect 2405 7714 2471 7717
rect 62 7712 2471 7714
rect 62 7656 2410 7712
rect 2466 7656 2471 7712
rect 62 7654 2471 7656
rect 2405 7651 2471 7654
rect 5758 7652 5764 7716
rect 5828 7714 5834 7716
rect 8569 7714 8635 7717
rect 5828 7712 8635 7714
rect 5828 7656 8574 7712
rect 8630 7656 8635 7712
rect 5828 7654 8635 7656
rect 5828 7652 5834 7654
rect 8569 7651 8635 7654
rect 10777 7714 10843 7717
rect 12758 7714 12818 7790
rect 15561 7787 15627 7790
rect 19290 7848 21699 7850
rect 19290 7792 21638 7848
rect 21694 7792 21699 7848
rect 19290 7790 21699 7792
rect 14181 7714 14247 7717
rect 19290 7714 19350 7790
rect 21633 7787 21699 7790
rect 10777 7712 12818 7714
rect 10777 7656 10782 7712
rect 10838 7656 12818 7712
rect 10777 7654 12818 7656
rect 13356 7712 19350 7714
rect 13356 7656 14186 7712
rect 14242 7656 19350 7712
rect 13356 7654 19350 7656
rect 10777 7651 10843 7654
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 2998 7516 3004 7580
rect 3068 7578 3074 7580
rect 3141 7578 3207 7581
rect 3068 7576 3207 7578
rect 3068 7520 3146 7576
rect 3202 7520 3207 7576
rect 3068 7518 3207 7520
rect 3068 7516 3074 7518
rect 3141 7515 3207 7518
rect 6177 7578 6243 7581
rect 8385 7578 8451 7581
rect 9121 7578 9187 7581
rect 6177 7576 7850 7578
rect 6177 7520 6182 7576
rect 6238 7520 7850 7576
rect 6177 7518 7850 7520
rect 6177 7515 6243 7518
rect 0 7440 480 7472
rect 0 7384 110 7440
rect 166 7384 480 7440
rect 0 7352 480 7384
rect 1853 7442 1919 7445
rect 3417 7442 3483 7445
rect 7281 7442 7347 7445
rect 1853 7440 3112 7442
rect 1853 7384 1858 7440
rect 1914 7384 3112 7440
rect 1853 7382 3112 7384
rect 1853 7379 1919 7382
rect 3052 7306 3112 7382
rect 3417 7440 7347 7442
rect 3417 7384 3422 7440
rect 3478 7384 7286 7440
rect 7342 7384 7347 7440
rect 3417 7382 7347 7384
rect 7790 7442 7850 7518
rect 8385 7576 9187 7578
rect 8385 7520 8390 7576
rect 8446 7520 9126 7576
rect 9182 7520 9187 7576
rect 8385 7518 9187 7520
rect 8385 7515 8451 7518
rect 9121 7515 9187 7518
rect 9397 7578 9463 7581
rect 12014 7578 12020 7580
rect 9397 7576 12020 7578
rect 9397 7520 9402 7576
rect 9458 7520 12020 7576
rect 9397 7518 12020 7520
rect 9397 7515 9463 7518
rect 12014 7516 12020 7518
rect 12084 7516 12090 7580
rect 9806 7442 9812 7444
rect 7790 7382 9812 7442
rect 3417 7379 3483 7382
rect 7281 7379 7347 7382
rect 9806 7380 9812 7382
rect 9876 7380 9882 7444
rect 12893 7442 12959 7445
rect 13356 7442 13416 7654
rect 14181 7651 14247 7654
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 13486 7516 13492 7580
rect 13556 7578 13562 7580
rect 14733 7578 14799 7581
rect 13556 7576 14799 7578
rect 13556 7520 14738 7576
rect 14794 7520 14799 7576
rect 13556 7518 14799 7520
rect 13556 7516 13562 7518
rect 14733 7515 14799 7518
rect 18321 7578 18387 7581
rect 18454 7578 18460 7580
rect 18321 7576 18460 7578
rect 18321 7520 18326 7576
rect 18382 7520 18460 7576
rect 18321 7518 18460 7520
rect 18321 7515 18387 7518
rect 18454 7516 18460 7518
rect 18524 7516 18530 7580
rect 12893 7440 13416 7442
rect 12893 7384 12898 7440
rect 12954 7384 13416 7440
rect 12893 7382 13416 7384
rect 15009 7442 15075 7445
rect 19793 7442 19859 7445
rect 15009 7440 19859 7442
rect 15009 7384 15014 7440
rect 15070 7384 19798 7440
rect 19854 7384 19859 7440
rect 15009 7382 19859 7384
rect 12893 7379 12959 7382
rect 15009 7379 15075 7382
rect 19793 7379 19859 7382
rect 10501 7306 10567 7309
rect 3052 7304 10567 7306
rect 3052 7248 10506 7304
rect 10562 7248 10567 7304
rect 3052 7246 10567 7248
rect 10501 7243 10567 7246
rect 10961 7306 11027 7309
rect 15009 7306 15075 7309
rect 10961 7304 15075 7306
rect 10961 7248 10966 7304
rect 11022 7248 15014 7304
rect 15070 7248 15075 7304
rect 10961 7246 15075 7248
rect 10961 7243 11027 7246
rect 15009 7243 15075 7246
rect 15561 7306 15627 7309
rect 19241 7306 19307 7309
rect 15561 7304 19307 7306
rect 15561 7248 15566 7304
rect 15622 7248 19246 7304
rect 19302 7248 19307 7304
rect 15561 7246 19307 7248
rect 15561 7243 15627 7246
rect 19241 7243 19307 7246
rect 2630 7108 2636 7172
rect 2700 7170 2706 7172
rect 2957 7170 3023 7173
rect 2700 7168 3023 7170
rect 2700 7112 2962 7168
rect 3018 7112 3023 7168
rect 2700 7110 3023 7112
rect 2700 7108 2706 7110
rect 2957 7107 3023 7110
rect 3417 7170 3483 7173
rect 3969 7170 4035 7173
rect 3417 7168 4035 7170
rect 3417 7112 3422 7168
rect 3478 7112 3974 7168
rect 4030 7112 4035 7168
rect 3417 7110 4035 7112
rect 3417 7107 3483 7110
rect 3969 7107 4035 7110
rect 4153 7170 4219 7173
rect 4286 7170 4292 7172
rect 4153 7168 4292 7170
rect 4153 7112 4158 7168
rect 4214 7112 4292 7168
rect 4153 7110 4292 7112
rect 4153 7107 4219 7110
rect 4286 7108 4292 7110
rect 4356 7108 4362 7172
rect 5993 7170 6059 7173
rect 6126 7170 6132 7172
rect 5993 7168 6132 7170
rect 5993 7112 5998 7168
rect 6054 7112 6132 7168
rect 5993 7110 6132 7112
rect 5993 7107 6059 7110
rect 6126 7108 6132 7110
rect 6196 7108 6202 7172
rect 6545 7170 6611 7173
rect 6678 7170 6684 7172
rect 6545 7168 6684 7170
rect 6545 7112 6550 7168
rect 6606 7112 6684 7168
rect 6545 7110 6684 7112
rect 6545 7107 6611 7110
rect 6678 7108 6684 7110
rect 6748 7108 6754 7172
rect 9397 7170 9463 7173
rect 15745 7170 15811 7173
rect 23520 7170 24000 7200
rect 9397 7168 15811 7170
rect 9397 7112 9402 7168
rect 9458 7112 15750 7168
rect 15806 7112 15811 7168
rect 9397 7110 15811 7112
rect 23484 7168 24000 7170
rect 23484 7112 23570 7168
rect 23626 7112 24000 7168
rect 23484 7110 24000 7112
rect 9397 7107 9463 7110
rect 15745 7107 15811 7110
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 23520 7080 24000 7110
rect 16944 7039 17264 7040
rect 7005 7034 7071 7037
rect 62 7032 7071 7034
rect 62 6976 7010 7032
rect 7066 6976 7071 7032
rect 62 6974 7071 6976
rect 62 6656 122 6974
rect 7005 6971 7071 6974
rect 3049 6898 3115 6901
rect 11881 6898 11947 6901
rect 3049 6896 11947 6898
rect 3049 6840 3054 6896
rect 3110 6840 11886 6896
rect 11942 6840 11947 6896
rect 3049 6838 11947 6840
rect 3049 6835 3115 6838
rect 11881 6835 11947 6838
rect 13905 6898 13971 6901
rect 18137 6898 18203 6901
rect 13905 6896 18203 6898
rect 13905 6840 13910 6896
rect 13966 6840 18142 6896
rect 18198 6840 18203 6896
rect 13905 6838 18203 6840
rect 13905 6835 13971 6838
rect 18137 6835 18203 6838
rect 2037 6762 2103 6765
rect 3969 6762 4035 6765
rect 4889 6762 4955 6765
rect 2037 6760 4035 6762
rect 2037 6704 2042 6760
rect 2098 6704 3974 6760
rect 4030 6704 4035 6760
rect 2037 6702 4035 6704
rect 2037 6699 2103 6702
rect 3969 6699 4035 6702
rect 4110 6760 4955 6762
rect 4110 6704 4894 6760
rect 4950 6704 4955 6760
rect 4110 6702 4955 6704
rect 0 6536 480 6656
rect 1669 6626 1735 6629
rect 4110 6626 4170 6702
rect 4889 6699 4955 6702
rect 5165 6762 5231 6765
rect 7782 6762 7788 6764
rect 5165 6760 7788 6762
rect 5165 6704 5170 6760
rect 5226 6704 7788 6760
rect 5165 6702 7788 6704
rect 5165 6699 5231 6702
rect 7782 6700 7788 6702
rect 7852 6762 7858 6764
rect 8385 6762 8451 6765
rect 7852 6760 8451 6762
rect 7852 6704 8390 6760
rect 8446 6704 8451 6760
rect 7852 6702 8451 6704
rect 7852 6700 7858 6702
rect 8385 6699 8451 6702
rect 12801 6762 12867 6765
rect 20621 6762 20687 6765
rect 12801 6760 20687 6762
rect 12801 6704 12806 6760
rect 12862 6704 20626 6760
rect 20682 6704 20687 6760
rect 12801 6702 20687 6704
rect 12801 6699 12867 6702
rect 20621 6699 20687 6702
rect 1669 6624 4170 6626
rect 1669 6568 1674 6624
rect 1730 6568 4170 6624
rect 1669 6566 4170 6568
rect 1669 6563 1735 6566
rect 6126 6564 6132 6628
rect 6196 6626 6202 6628
rect 8109 6626 8175 6629
rect 6196 6624 8175 6626
rect 6196 6568 8114 6624
rect 8170 6568 8175 6624
rect 6196 6566 8175 6568
rect 6196 6564 6202 6566
rect 8109 6563 8175 6566
rect 22185 6626 22251 6629
rect 22185 6624 23674 6626
rect 22185 6568 22190 6624
rect 22246 6568 23674 6624
rect 22185 6566 23674 6568
rect 22185 6563 22251 6566
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 2078 6428 2084 6492
rect 2148 6490 2154 6492
rect 2681 6490 2747 6493
rect 2148 6488 2747 6490
rect 2148 6432 2686 6488
rect 2742 6432 2747 6488
rect 2148 6430 2747 6432
rect 2148 6428 2154 6430
rect 2681 6427 2747 6430
rect 2814 6428 2820 6492
rect 2884 6490 2890 6492
rect 3969 6490 4035 6493
rect 9673 6490 9739 6493
rect 11145 6490 11211 6493
rect 2884 6488 4035 6490
rect 2884 6432 3974 6488
rect 4030 6432 4035 6488
rect 2884 6430 4035 6432
rect 2884 6428 2890 6430
rect 3969 6427 4035 6430
rect 5996 6488 11211 6490
rect 5996 6432 9678 6488
rect 9734 6432 11150 6488
rect 11206 6432 11211 6488
rect 5996 6430 11211 6432
rect 1577 6354 1643 6357
rect 62 6352 1643 6354
rect 62 6296 1582 6352
rect 1638 6296 1643 6352
rect 62 6294 1643 6296
rect 62 5976 122 6294
rect 1577 6291 1643 6294
rect 4153 6354 4219 6357
rect 5996 6354 6056 6430
rect 9673 6427 9739 6430
rect 11145 6427 11211 6430
rect 14365 6490 14431 6493
rect 20713 6492 20779 6493
rect 20662 6490 20668 6492
rect 14365 6488 20668 6490
rect 20732 6488 20779 6492
rect 14365 6432 14370 6488
rect 14426 6432 20668 6488
rect 20774 6432 20779 6488
rect 14365 6430 20668 6432
rect 14365 6427 14431 6430
rect 20662 6428 20668 6430
rect 20732 6428 20779 6432
rect 20713 6427 20779 6428
rect 4153 6352 6056 6354
rect 4153 6296 4158 6352
rect 4214 6296 6056 6352
rect 4153 6294 6056 6296
rect 6269 6354 6335 6357
rect 16849 6354 16915 6357
rect 6269 6352 16915 6354
rect 6269 6296 6274 6352
rect 6330 6296 16854 6352
rect 16910 6296 16915 6352
rect 6269 6294 16915 6296
rect 4153 6291 4219 6294
rect 6269 6291 6335 6294
rect 16849 6291 16915 6294
rect 17585 6354 17651 6357
rect 19926 6354 19932 6356
rect 17585 6352 19932 6354
rect 17585 6296 17590 6352
rect 17646 6296 19932 6352
rect 17585 6294 19932 6296
rect 17585 6291 17651 6294
rect 19926 6292 19932 6294
rect 19996 6292 20002 6356
rect 2865 6218 2931 6221
rect 3182 6218 3188 6220
rect 2865 6216 3188 6218
rect 2865 6160 2870 6216
rect 2926 6160 3188 6216
rect 2865 6158 3188 6160
rect 2865 6155 2931 6158
rect 3182 6156 3188 6158
rect 3252 6156 3258 6220
rect 3877 6218 3943 6221
rect 4102 6218 4108 6220
rect 3877 6216 4108 6218
rect 3877 6160 3882 6216
rect 3938 6160 4108 6216
rect 3877 6158 4108 6160
rect 3877 6155 3943 6158
rect 4102 6156 4108 6158
rect 4172 6156 4178 6220
rect 4286 6156 4292 6220
rect 4356 6218 4362 6220
rect 4429 6218 4495 6221
rect 4356 6216 4495 6218
rect 4356 6160 4434 6216
rect 4490 6160 4495 6216
rect 4356 6158 4495 6160
rect 4356 6156 4362 6158
rect 4429 6155 4495 6158
rect 5809 6218 5875 6221
rect 5942 6218 5948 6220
rect 5809 6216 5948 6218
rect 5809 6160 5814 6216
rect 5870 6160 5948 6216
rect 5809 6158 5948 6160
rect 5809 6155 5875 6158
rect 5942 6156 5948 6158
rect 6012 6156 6018 6220
rect 7598 6156 7604 6220
rect 7668 6218 7674 6220
rect 15837 6218 15903 6221
rect 7668 6216 15903 6218
rect 7668 6160 15842 6216
rect 15898 6160 15903 6216
rect 7668 6158 15903 6160
rect 7668 6156 7674 6158
rect 15837 6155 15903 6158
rect 16573 6218 16639 6221
rect 17534 6218 17540 6220
rect 16573 6216 17540 6218
rect 16573 6160 16578 6216
rect 16634 6160 17540 6216
rect 16573 6158 17540 6160
rect 16573 6155 16639 6158
rect 17534 6156 17540 6158
rect 17604 6156 17610 6220
rect 23614 6112 23674 6566
rect 1485 6082 1551 6085
rect 1710 6082 1716 6084
rect 1485 6080 1716 6082
rect 1485 6024 1490 6080
rect 1546 6024 1716 6080
rect 1485 6022 1716 6024
rect 1485 6019 1551 6022
rect 1710 6020 1716 6022
rect 1780 6020 1786 6084
rect 2681 6082 2747 6085
rect 7281 6082 7347 6085
rect 2681 6080 7347 6082
rect 2681 6024 2686 6080
rect 2742 6024 7286 6080
rect 7342 6024 7347 6080
rect 2681 6022 7347 6024
rect 2681 6019 2747 6022
rect 7281 6019 7347 6022
rect 9673 6082 9739 6085
rect 16798 6082 16804 6084
rect 9673 6080 16804 6082
rect 9673 6024 9678 6080
rect 9734 6024 16804 6080
rect 9673 6022 16804 6024
rect 9673 6019 9739 6022
rect 16798 6020 16804 6022
rect 16868 6020 16874 6084
rect 18822 6020 18828 6084
rect 18892 6082 18898 6084
rect 18965 6082 19031 6085
rect 18892 6080 19031 6082
rect 18892 6024 18970 6080
rect 19026 6024 19031 6080
rect 18892 6022 19031 6024
rect 18892 6020 18898 6022
rect 18965 6019 19031 6022
rect 8944 6016 9264 6017
rect 0 5856 480 5976
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 23520 5992 24000 6112
rect 16944 5951 17264 5952
rect 1342 5884 1348 5948
rect 1412 5946 1418 5948
rect 2221 5946 2287 5949
rect 8293 5946 8359 5949
rect 8569 5946 8635 5949
rect 1412 5944 8635 5946
rect 1412 5888 2226 5944
rect 2282 5888 8298 5944
rect 8354 5888 8574 5944
rect 8630 5888 8635 5944
rect 1412 5886 8635 5888
rect 1412 5884 1418 5886
rect 2221 5883 2287 5886
rect 8293 5883 8359 5886
rect 8569 5883 8635 5886
rect 9397 5946 9463 5949
rect 16481 5946 16547 5949
rect 9397 5944 16547 5946
rect 9397 5888 9402 5944
rect 9458 5888 16486 5944
rect 16542 5888 16547 5944
rect 9397 5886 16547 5888
rect 9397 5883 9463 5886
rect 16481 5883 16547 5886
rect 17677 5946 17743 5949
rect 18086 5946 18092 5948
rect 17677 5944 18092 5946
rect 17677 5888 17682 5944
rect 17738 5888 18092 5944
rect 17677 5886 18092 5888
rect 17677 5883 17743 5886
rect 18086 5884 18092 5886
rect 18156 5884 18162 5948
rect 3877 5810 3943 5813
rect 4470 5810 4476 5812
rect 3877 5808 4476 5810
rect 3877 5752 3882 5808
rect 3938 5752 4476 5808
rect 3877 5750 4476 5752
rect 3877 5747 3943 5750
rect 4470 5748 4476 5750
rect 4540 5810 4546 5812
rect 5165 5810 5231 5813
rect 4540 5808 5231 5810
rect 4540 5752 5170 5808
rect 5226 5752 5231 5808
rect 4540 5750 5231 5752
rect 4540 5748 4546 5750
rect 5165 5747 5231 5750
rect 6637 5810 6703 5813
rect 9990 5810 9996 5812
rect 6637 5808 9996 5810
rect 6637 5752 6642 5808
rect 6698 5752 9996 5808
rect 6637 5750 9996 5752
rect 6637 5747 6703 5750
rect 9990 5748 9996 5750
rect 10060 5748 10066 5812
rect 10133 5810 10199 5813
rect 18321 5810 18387 5813
rect 10133 5808 18387 5810
rect 10133 5752 10138 5808
rect 10194 5752 18326 5808
rect 18382 5752 18387 5808
rect 10133 5750 18387 5752
rect 10133 5747 10199 5750
rect 18321 5747 18387 5750
rect 4061 5674 4127 5677
rect 6177 5674 6243 5677
rect 4061 5672 6243 5674
rect 4061 5616 4066 5672
rect 4122 5616 6182 5672
rect 6238 5616 6243 5672
rect 4061 5614 6243 5616
rect 4061 5611 4127 5614
rect 6177 5611 6243 5614
rect 7833 5674 7899 5677
rect 17861 5674 17927 5677
rect 7833 5672 17927 5674
rect 7833 5616 7838 5672
rect 7894 5616 17866 5672
rect 17922 5616 17927 5672
rect 7833 5614 17927 5616
rect 7833 5611 7899 5614
rect 17861 5611 17927 5614
rect 4470 5476 4476 5540
rect 4540 5538 4546 5540
rect 4705 5538 4771 5541
rect 4540 5536 4771 5538
rect 4540 5480 4710 5536
rect 4766 5480 4771 5536
rect 4540 5478 4771 5480
rect 4540 5476 4546 5478
rect 4705 5475 4771 5478
rect 5574 5476 5580 5540
rect 5644 5538 5650 5540
rect 9949 5538 10015 5541
rect 5644 5536 10015 5538
rect 5644 5480 9954 5536
rect 10010 5480 10015 5536
rect 5644 5478 10015 5480
rect 5644 5476 5650 5478
rect 9949 5475 10015 5478
rect 10726 5476 10732 5540
rect 10796 5538 10802 5540
rect 11094 5538 11100 5540
rect 10796 5478 11100 5538
rect 10796 5476 10802 5478
rect 11094 5476 11100 5478
rect 11164 5476 11170 5540
rect 11646 5476 11652 5540
rect 11716 5538 11722 5540
rect 11789 5538 11855 5541
rect 11716 5536 11855 5538
rect 11716 5480 11794 5536
rect 11850 5480 11855 5536
rect 11716 5478 11855 5480
rect 11716 5476 11722 5478
rect 11789 5475 11855 5478
rect 16297 5538 16363 5541
rect 18689 5538 18755 5541
rect 16297 5536 18755 5538
rect 16297 5480 16302 5536
rect 16358 5480 18694 5536
rect 18750 5480 18755 5536
rect 16297 5478 18755 5480
rect 16297 5475 16363 5478
rect 18689 5475 18755 5478
rect 22645 5538 22711 5541
rect 22645 5536 23674 5538
rect 22645 5480 22650 5536
rect 22706 5480 23674 5536
rect 22645 5478 23674 5480
rect 22645 5475 22711 5478
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 9029 5402 9095 5405
rect 10041 5402 10107 5405
rect 9029 5400 10107 5402
rect 9029 5344 9034 5400
rect 9090 5344 10046 5400
rect 10102 5344 10107 5400
rect 9029 5342 10107 5344
rect 9029 5339 9095 5342
rect 10041 5339 10107 5342
rect 10317 5402 10383 5405
rect 12382 5402 12388 5404
rect 10317 5400 12388 5402
rect 10317 5344 10322 5400
rect 10378 5344 12388 5400
rect 10317 5342 12388 5344
rect 10317 5339 10383 5342
rect 12382 5340 12388 5342
rect 12452 5340 12458 5404
rect 13537 5402 13603 5405
rect 14365 5402 14431 5405
rect 13537 5400 14431 5402
rect 13537 5344 13542 5400
rect 13598 5344 14370 5400
rect 14426 5344 14431 5400
rect 13537 5342 14431 5344
rect 13537 5339 13603 5342
rect 14365 5339 14431 5342
rect 14549 5402 14615 5405
rect 17861 5402 17927 5405
rect 14549 5400 17927 5402
rect 14549 5344 14554 5400
rect 14610 5344 17866 5400
rect 17922 5344 17927 5400
rect 14549 5342 17927 5344
rect 14549 5339 14615 5342
rect 17861 5339 17927 5342
rect 19241 5400 19307 5405
rect 19241 5344 19246 5400
rect 19302 5344 19307 5400
rect 19241 5339 19307 5344
rect 5257 5266 5323 5269
rect 15653 5266 15719 5269
rect 5257 5264 15719 5266
rect 5257 5208 5262 5264
rect 5318 5208 15658 5264
rect 15714 5208 15719 5264
rect 5257 5206 15719 5208
rect 5257 5203 5323 5206
rect 15653 5203 15719 5206
rect 16389 5266 16455 5269
rect 18413 5266 18479 5269
rect 16389 5264 18479 5266
rect 16389 5208 16394 5264
rect 16450 5208 18418 5264
rect 18474 5208 18479 5264
rect 16389 5206 18479 5208
rect 16389 5203 16455 5206
rect 18413 5203 18479 5206
rect 0 5128 480 5160
rect 0 5072 18 5128
rect 74 5072 480 5128
rect 0 5040 480 5072
rect 4153 5130 4219 5133
rect 8937 5130 9003 5133
rect 4153 5128 9003 5130
rect 4153 5072 4158 5128
rect 4214 5072 8942 5128
rect 8998 5072 9003 5128
rect 4153 5070 9003 5072
rect 4153 5067 4219 5070
rect 8937 5067 9003 5070
rect 12801 5130 12867 5133
rect 14038 5130 14044 5132
rect 12801 5128 14044 5130
rect 12801 5072 12806 5128
rect 12862 5072 14044 5128
rect 12801 5070 14044 5072
rect 12801 5067 12867 5070
rect 14038 5068 14044 5070
rect 14108 5068 14114 5132
rect 15142 5068 15148 5132
rect 15212 5130 15218 5132
rect 15469 5130 15535 5133
rect 15212 5128 15535 5130
rect 15212 5072 15474 5128
rect 15530 5072 15535 5128
rect 15212 5070 15535 5072
rect 15212 5068 15218 5070
rect 15469 5067 15535 5070
rect 16113 5130 16179 5133
rect 19244 5130 19304 5339
rect 16113 5128 19304 5130
rect 16113 5072 16118 5128
rect 16174 5072 19304 5128
rect 16113 5070 19304 5072
rect 16113 5067 16179 5070
rect 19742 5068 19748 5132
rect 19812 5130 19818 5132
rect 20529 5130 20595 5133
rect 19812 5128 20595 5130
rect 19812 5072 20534 5128
rect 20590 5072 20595 5128
rect 19812 5070 20595 5072
rect 19812 5068 19818 5070
rect 20529 5067 20595 5070
rect 20662 5068 20668 5132
rect 20732 5130 20738 5132
rect 22277 5130 22343 5133
rect 20732 5128 22343 5130
rect 20732 5072 22282 5128
rect 22338 5072 22343 5128
rect 20732 5070 22343 5072
rect 20732 5068 20738 5070
rect 22277 5067 22343 5070
rect 23614 5024 23674 5478
rect 1894 4932 1900 4996
rect 1964 4994 1970 4996
rect 5993 4994 6059 4997
rect 1964 4992 6059 4994
rect 1964 4936 5998 4992
rect 6054 4936 6059 4992
rect 1964 4934 6059 4936
rect 1964 4932 1970 4934
rect 5993 4931 6059 4934
rect 7833 4994 7899 4997
rect 8150 4994 8156 4996
rect 7833 4992 8156 4994
rect 7833 4936 7838 4992
rect 7894 4936 8156 4992
rect 7833 4934 8156 4936
rect 7833 4931 7899 4934
rect 8150 4932 8156 4934
rect 8220 4932 8226 4996
rect 9857 4994 9923 4997
rect 9990 4994 9996 4996
rect 9857 4992 9996 4994
rect 9857 4936 9862 4992
rect 9918 4936 9996 4992
rect 9857 4934 9996 4936
rect 9857 4931 9923 4934
rect 9990 4932 9996 4934
rect 10060 4932 10066 4996
rect 10133 4994 10199 4997
rect 11830 4994 11836 4996
rect 10133 4992 11836 4994
rect 10133 4936 10138 4992
rect 10194 4936 11836 4992
rect 10133 4934 11836 4936
rect 10133 4931 10199 4934
rect 11830 4932 11836 4934
rect 11900 4932 11906 4996
rect 12566 4932 12572 4996
rect 12636 4994 12642 4996
rect 12801 4994 12867 4997
rect 12636 4992 12867 4994
rect 12636 4936 12806 4992
rect 12862 4936 12867 4992
rect 12636 4934 12867 4936
rect 12636 4932 12642 4934
rect 12801 4931 12867 4934
rect 17493 4994 17559 4997
rect 20989 4994 21055 4997
rect 17493 4992 21055 4994
rect 17493 4936 17498 4992
rect 17554 4936 20994 4992
rect 21050 4936 21055 4992
rect 17493 4934 21055 4936
rect 17493 4931 17559 4934
rect 20989 4931 21055 4934
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 23520 4904 24000 5024
rect 16944 4863 17264 4864
rect 238 4858 244 4860
rect 62 4798 244 4858
rect 62 4344 122 4798
rect 238 4796 244 4798
rect 308 4796 314 4860
rect 4705 4858 4771 4861
rect 5758 4858 5764 4860
rect 4705 4856 5764 4858
rect 4705 4800 4710 4856
rect 4766 4800 5764 4856
rect 4705 4798 5764 4800
rect 4705 4795 4771 4798
rect 5758 4796 5764 4798
rect 5828 4796 5834 4860
rect 6494 4796 6500 4860
rect 6564 4858 6570 4860
rect 6637 4858 6703 4861
rect 6564 4856 6703 4858
rect 6564 4800 6642 4856
rect 6698 4800 6703 4856
rect 6564 4798 6703 4800
rect 6564 4796 6570 4798
rect 6637 4795 6703 4798
rect 7966 4796 7972 4860
rect 8036 4858 8042 4860
rect 8109 4858 8175 4861
rect 8036 4856 8175 4858
rect 8036 4800 8114 4856
rect 8170 4800 8175 4856
rect 8036 4798 8175 4800
rect 8036 4796 8042 4798
rect 8109 4795 8175 4798
rect 9673 4858 9739 4861
rect 9806 4858 9812 4860
rect 9673 4856 9812 4858
rect 9673 4800 9678 4856
rect 9734 4800 9812 4856
rect 9673 4798 9812 4800
rect 9673 4795 9739 4798
rect 9806 4796 9812 4798
rect 9876 4796 9882 4860
rect 10174 4796 10180 4860
rect 10244 4858 10250 4860
rect 10593 4858 10659 4861
rect 16757 4858 16823 4861
rect 10244 4856 16823 4858
rect 10244 4800 10598 4856
rect 10654 4800 16762 4856
rect 16818 4800 16823 4856
rect 10244 4798 16823 4800
rect 10244 4796 10250 4798
rect 10593 4795 10659 4798
rect 16757 4795 16823 4798
rect 19149 4858 19215 4861
rect 20110 4858 20116 4860
rect 19149 4856 20116 4858
rect 19149 4800 19154 4856
rect 19210 4800 20116 4856
rect 19149 4798 20116 4800
rect 19149 4795 19215 4798
rect 20110 4796 20116 4798
rect 20180 4796 20186 4860
rect 3734 4660 3740 4724
rect 3804 4722 3810 4724
rect 3969 4722 4035 4725
rect 3804 4720 4035 4722
rect 3804 4664 3974 4720
rect 4030 4664 4035 4720
rect 3804 4662 4035 4664
rect 3804 4660 3810 4662
rect 3969 4659 4035 4662
rect 4429 4722 4495 4725
rect 13721 4722 13787 4725
rect 4429 4720 13787 4722
rect 4429 4664 4434 4720
rect 4490 4664 13726 4720
rect 13782 4664 13787 4720
rect 4429 4662 13787 4664
rect 4429 4659 4495 4662
rect 13721 4659 13787 4662
rect 16113 4722 16179 4725
rect 19609 4722 19675 4725
rect 16113 4720 19675 4722
rect 16113 4664 16118 4720
rect 16174 4664 19614 4720
rect 19670 4664 19675 4720
rect 16113 4662 19675 4664
rect 16113 4659 16179 4662
rect 19609 4659 19675 4662
rect 19926 4660 19932 4724
rect 19996 4722 20002 4724
rect 20069 4722 20135 4725
rect 22461 4722 22527 4725
rect 19996 4720 22527 4722
rect 19996 4664 20074 4720
rect 20130 4664 22466 4720
rect 22522 4664 22527 4720
rect 19996 4662 22527 4664
rect 19996 4660 20002 4662
rect 20069 4659 20135 4662
rect 22461 4659 22527 4662
rect 3509 4586 3575 4589
rect 8385 4586 8451 4589
rect 9489 4586 9555 4589
rect 3509 4584 9555 4586
rect 3509 4528 3514 4584
rect 3570 4528 8390 4584
rect 8446 4528 9494 4584
rect 9550 4528 9555 4584
rect 3509 4526 9555 4528
rect 3509 4523 3575 4526
rect 8385 4523 8451 4526
rect 9489 4523 9555 4526
rect 10225 4586 10291 4589
rect 12566 4586 12572 4588
rect 10225 4584 12572 4586
rect 10225 4528 10230 4584
rect 10286 4528 12572 4584
rect 10225 4526 12572 4528
rect 10225 4523 10291 4526
rect 12566 4524 12572 4526
rect 12636 4524 12642 4588
rect 12893 4586 12959 4589
rect 14365 4586 14431 4589
rect 17861 4586 17927 4589
rect 20345 4586 20411 4589
rect 12893 4584 17927 4586
rect 12893 4528 12898 4584
rect 12954 4528 14370 4584
rect 14426 4528 17866 4584
rect 17922 4528 17927 4584
rect 12893 4526 17927 4528
rect 12893 4523 12959 4526
rect 14365 4523 14431 4526
rect 17861 4523 17927 4526
rect 18048 4584 20411 4586
rect 18048 4528 20350 4584
rect 20406 4528 20411 4584
rect 18048 4526 20411 4528
rect 5901 4450 5967 4453
rect 8017 4450 8083 4453
rect 5901 4448 8083 4450
rect 5901 4392 5906 4448
rect 5962 4392 8022 4448
rect 8078 4392 8083 4448
rect 5901 4390 8083 4392
rect 5901 4387 5967 4390
rect 8017 4387 8083 4390
rect 8845 4450 8911 4453
rect 9990 4450 9996 4452
rect 8845 4448 9996 4450
rect 8845 4392 8850 4448
rect 8906 4392 9996 4448
rect 8845 4390 9996 4392
rect 8845 4387 8911 4390
rect 9990 4388 9996 4390
rect 10060 4388 10066 4452
rect 11329 4450 11395 4453
rect 15929 4450 15995 4453
rect 18048 4450 18108 4526
rect 20345 4523 20411 4526
rect 10136 4448 11395 4450
rect 10136 4392 11334 4448
rect 11390 4392 11395 4448
rect 10136 4390 11395 4392
rect 4944 4384 5264 4385
rect 0 4224 480 4344
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 790 4252 796 4316
rect 860 4314 866 4316
rect 2681 4314 2747 4317
rect 860 4312 2747 4314
rect 860 4256 2686 4312
rect 2742 4256 2747 4312
rect 860 4254 2747 4256
rect 860 4252 866 4254
rect 2681 4251 2747 4254
rect 6085 4314 6151 4317
rect 6310 4314 6316 4316
rect 6085 4312 6316 4314
rect 6085 4256 6090 4312
rect 6146 4256 6316 4312
rect 6085 4254 6316 4256
rect 6085 4251 6151 4254
rect 6310 4252 6316 4254
rect 6380 4252 6386 4316
rect 6729 4314 6795 4317
rect 7230 4314 7236 4316
rect 6729 4312 7236 4314
rect 6729 4256 6734 4312
rect 6790 4256 7236 4312
rect 6729 4254 7236 4256
rect 6729 4251 6795 4254
rect 7230 4252 7236 4254
rect 7300 4252 7306 4316
rect 7557 4314 7623 4317
rect 7741 4314 7807 4317
rect 7557 4312 7807 4314
rect 7557 4256 7562 4312
rect 7618 4256 7746 4312
rect 7802 4256 7807 4312
rect 7557 4254 7807 4256
rect 7557 4251 7623 4254
rect 7741 4251 7807 4254
rect 8017 4314 8083 4317
rect 8334 4314 8340 4316
rect 8017 4312 8340 4314
rect 8017 4256 8022 4312
rect 8078 4256 8340 4312
rect 8017 4254 8340 4256
rect 8017 4251 8083 4254
rect 8334 4252 8340 4254
rect 8404 4252 8410 4316
rect 8518 4252 8524 4316
rect 8588 4252 8594 4316
rect 9765 4314 9831 4317
rect 10136 4314 10196 4390
rect 11329 4387 11395 4390
rect 13770 4448 18108 4450
rect 13770 4392 15934 4448
rect 15990 4392 18108 4448
rect 13770 4390 18108 4392
rect 18873 4450 18939 4453
rect 19885 4450 19951 4453
rect 18873 4448 19951 4450
rect 18873 4392 18878 4448
rect 18934 4392 19890 4448
rect 19946 4392 19951 4448
rect 18873 4390 19951 4392
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 9078 4254 9690 4314
rect 3417 4178 3483 4181
rect 4153 4178 4219 4181
rect 3417 4176 4219 4178
rect 3417 4120 3422 4176
rect 3478 4120 4158 4176
rect 4214 4120 4219 4176
rect 3417 4118 4219 4120
rect 3417 4115 3483 4118
rect 4153 4115 4219 4118
rect 4429 4178 4495 4181
rect 6678 4178 6684 4180
rect 4429 4176 6684 4178
rect 4429 4120 4434 4176
rect 4490 4120 6684 4176
rect 4429 4118 6684 4120
rect 4429 4115 4495 4118
rect 6678 4116 6684 4118
rect 6748 4116 6754 4180
rect 7925 4178 7991 4181
rect 8526 4178 8586 4252
rect 7925 4176 8586 4178
rect 7925 4120 7930 4176
rect 7986 4120 8586 4176
rect 7925 4118 8586 4120
rect 7925 4115 7991 4118
rect 2313 4042 2379 4045
rect 62 4040 2379 4042
rect 62 3984 2318 4040
rect 2374 3984 2379 4040
rect 62 3982 2379 3984
rect 62 3528 122 3982
rect 2313 3979 2379 3982
rect 3233 4042 3299 4045
rect 5533 4042 5599 4045
rect 3233 4040 5599 4042
rect 3233 3984 3238 4040
rect 3294 3984 5538 4040
rect 5594 3984 5599 4040
rect 3233 3982 5599 3984
rect 3233 3979 3299 3982
rect 5533 3979 5599 3982
rect 7005 4042 7071 4045
rect 8661 4042 8727 4045
rect 7005 4040 8727 4042
rect 7005 3984 7010 4040
rect 7066 3984 8666 4040
rect 8722 3984 8727 4040
rect 7005 3982 8727 3984
rect 9078 4042 9138 4254
rect 9213 4178 9279 4181
rect 9438 4178 9444 4180
rect 9213 4176 9444 4178
rect 9213 4120 9218 4176
rect 9274 4120 9444 4176
rect 9213 4118 9444 4120
rect 9213 4115 9279 4118
rect 9438 4116 9444 4118
rect 9508 4116 9514 4180
rect 9630 4178 9690 4254
rect 9765 4312 10196 4314
rect 9765 4256 9770 4312
rect 9826 4256 10196 4312
rect 9765 4254 10196 4256
rect 10593 4314 10659 4317
rect 10726 4314 10732 4316
rect 10593 4312 10732 4314
rect 10593 4256 10598 4312
rect 10654 4256 10732 4312
rect 10593 4254 10732 4256
rect 9765 4251 9831 4254
rect 10593 4251 10659 4254
rect 10726 4252 10732 4254
rect 10796 4252 10802 4316
rect 9857 4178 9923 4181
rect 9630 4176 9923 4178
rect 9630 4120 9862 4176
rect 9918 4120 9923 4176
rect 9630 4118 9923 4120
rect 9857 4115 9923 4118
rect 10133 4176 10199 4181
rect 10133 4120 10138 4176
rect 10194 4120 10199 4176
rect 10133 4115 10199 4120
rect 10317 4178 10383 4181
rect 13770 4178 13830 4390
rect 15929 4387 15995 4390
rect 18873 4387 18939 4390
rect 19885 4387 19951 4390
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 14089 4314 14155 4317
rect 18505 4314 18571 4317
rect 14089 4312 18571 4314
rect 14089 4256 14094 4312
rect 14150 4256 18510 4312
rect 18566 4256 18571 4312
rect 14089 4254 18571 4256
rect 14089 4251 14155 4254
rect 18505 4251 18571 4254
rect 18781 4314 18847 4317
rect 18965 4314 19031 4317
rect 18781 4312 19031 4314
rect 18781 4256 18786 4312
rect 18842 4256 18970 4312
rect 19026 4256 19031 4312
rect 18781 4254 19031 4256
rect 18781 4251 18847 4254
rect 18965 4251 19031 4254
rect 10317 4176 13830 4178
rect 10317 4120 10322 4176
rect 10378 4120 13830 4176
rect 10317 4118 13830 4120
rect 15285 4178 15351 4181
rect 18965 4178 19031 4181
rect 15285 4176 19031 4178
rect 15285 4120 15290 4176
rect 15346 4120 18970 4176
rect 19026 4120 19031 4176
rect 15285 4118 19031 4120
rect 10317 4115 10383 4118
rect 15285 4115 15351 4118
rect 18965 4115 19031 4118
rect 19977 4178 20043 4181
rect 21725 4178 21791 4181
rect 19977 4176 21791 4178
rect 19977 4120 19982 4176
rect 20038 4120 21730 4176
rect 21786 4120 21791 4176
rect 19977 4118 21791 4120
rect 19977 4115 20043 4118
rect 21725 4115 21791 4118
rect 9581 4042 9647 4045
rect 10136 4042 10196 4115
rect 9078 4008 9322 4042
rect 9581 4040 9690 4042
rect 9078 3982 9460 4008
rect 7005 3979 7071 3982
rect 8661 3979 8727 3982
rect 9262 3948 9460 3982
rect 9581 3984 9586 4040
rect 9642 4008 9690 4040
rect 9768 4008 10196 4042
rect 9642 3984 10196 4008
rect 9581 3982 10196 3984
rect 9581 3979 9828 3982
rect 9630 3948 9828 3979
rect 4102 3844 4108 3908
rect 4172 3906 4178 3908
rect 7046 3906 7052 3908
rect 4172 3846 7052 3906
rect 4172 3844 4178 3846
rect 7046 3844 7052 3846
rect 7116 3906 7122 3908
rect 8109 3906 8175 3909
rect 7116 3904 8175 3906
rect 7116 3848 8114 3904
rect 8170 3848 8175 3904
rect 7116 3846 8175 3848
rect 7116 3844 7122 3846
rect 8109 3843 8175 3846
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 1393 3770 1459 3773
rect 6126 3770 6132 3772
rect 1393 3768 6132 3770
rect 1393 3712 1398 3768
rect 1454 3712 6132 3768
rect 1393 3710 6132 3712
rect 1393 3707 1459 3710
rect 6126 3708 6132 3710
rect 6196 3708 6202 3772
rect 6494 3708 6500 3772
rect 6564 3770 6570 3772
rect 7465 3770 7531 3773
rect 6564 3768 7531 3770
rect 6564 3712 7470 3768
rect 7526 3712 7531 3768
rect 6564 3710 7531 3712
rect 6564 3708 6570 3710
rect 7465 3707 7531 3710
rect 7966 3708 7972 3772
rect 8036 3770 8042 3772
rect 8201 3770 8267 3773
rect 8036 3768 8267 3770
rect 8036 3712 8206 3768
rect 8262 3712 8267 3768
rect 8036 3710 8267 3712
rect 8036 3708 8042 3710
rect 8201 3707 8267 3710
rect 2446 3572 2452 3636
rect 2516 3634 2522 3636
rect 2681 3634 2747 3637
rect 2516 3632 2747 3634
rect 2516 3576 2686 3632
rect 2742 3576 2747 3632
rect 2516 3574 2747 3576
rect 2516 3572 2522 3574
rect 2681 3571 2747 3574
rect 3918 3572 3924 3636
rect 3988 3634 3994 3636
rect 4153 3634 4219 3637
rect 3988 3632 4219 3634
rect 3988 3576 4158 3632
rect 4214 3576 4219 3632
rect 3988 3574 4219 3576
rect 3988 3572 3994 3574
rect 4153 3571 4219 3574
rect 5574 3572 5580 3636
rect 5644 3634 5650 3636
rect 5717 3634 5783 3637
rect 5644 3632 5783 3634
rect 5644 3576 5722 3632
rect 5778 3576 5783 3632
rect 5644 3574 5783 3576
rect 5644 3572 5650 3574
rect 5717 3571 5783 3574
rect 5901 3634 5967 3637
rect 8109 3634 8175 3637
rect 5901 3632 8175 3634
rect 5901 3576 5906 3632
rect 5962 3576 8114 3632
rect 8170 3576 8175 3632
rect 5901 3574 8175 3576
rect 5901 3571 5967 3574
rect 8109 3571 8175 3574
rect 8293 3634 8359 3637
rect 9400 3634 9460 3948
rect 9952 3637 10012 3982
rect 10358 3980 10364 4044
rect 10428 4042 10434 4044
rect 10961 4042 11027 4045
rect 12065 4042 12131 4045
rect 18873 4042 18939 4045
rect 10428 4040 11944 4042
rect 10428 3984 10966 4040
rect 11022 3984 11944 4040
rect 10428 3982 11944 3984
rect 10428 3980 10434 3982
rect 10961 3979 11027 3982
rect 10133 3906 10199 3909
rect 10869 3906 10935 3909
rect 10133 3904 10935 3906
rect 10133 3848 10138 3904
rect 10194 3848 10874 3904
rect 10930 3848 10935 3904
rect 10133 3846 10935 3848
rect 11884 3906 11944 3982
rect 12065 4040 18939 4042
rect 12065 3984 12070 4040
rect 12126 3984 18878 4040
rect 18934 3984 18939 4040
rect 12065 3982 18939 3984
rect 12065 3979 12131 3982
rect 18873 3979 18939 3982
rect 19057 4042 19123 4045
rect 19517 4042 19583 4045
rect 19057 4040 19583 4042
rect 19057 3984 19062 4040
rect 19118 3984 19522 4040
rect 19578 3984 19583 4040
rect 19057 3982 19583 3984
rect 19057 3979 19123 3982
rect 19517 3979 19583 3982
rect 15745 3906 15811 3909
rect 11884 3904 15811 3906
rect 11884 3848 15750 3904
rect 15806 3848 15811 3904
rect 11884 3846 15811 3848
rect 10133 3843 10199 3846
rect 10869 3843 10935 3846
rect 15745 3843 15811 3846
rect 17401 3906 17467 3909
rect 18137 3906 18203 3909
rect 18454 3906 18460 3908
rect 17401 3904 18460 3906
rect 17401 3848 17406 3904
rect 17462 3848 18142 3904
rect 18198 3848 18460 3904
rect 17401 3846 18460 3848
rect 17401 3843 17467 3846
rect 18137 3843 18203 3846
rect 18454 3844 18460 3846
rect 18524 3844 18530 3908
rect 23520 3906 24000 3936
rect 23484 3904 24000 3906
rect 23484 3848 23570 3904
rect 23626 3848 24000 3904
rect 23484 3846 24000 3848
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 23520 3816 24000 3846
rect 16944 3775 17264 3776
rect 10317 3770 10383 3773
rect 15653 3770 15719 3773
rect 10317 3768 15719 3770
rect 10317 3712 10322 3768
rect 10378 3712 15658 3768
rect 15714 3712 15719 3768
rect 10317 3710 15719 3712
rect 10317 3707 10383 3710
rect 15653 3707 15719 3710
rect 15837 3770 15903 3773
rect 16205 3770 16271 3773
rect 15837 3768 16271 3770
rect 15837 3712 15842 3768
rect 15898 3712 16210 3768
rect 16266 3712 16271 3768
rect 15837 3710 16271 3712
rect 15837 3707 15903 3710
rect 16205 3707 16271 3710
rect 8293 3632 9460 3634
rect 8293 3576 8298 3632
rect 8354 3576 9460 3632
rect 8293 3574 9460 3576
rect 9949 3632 10015 3637
rect 9949 3576 9954 3632
rect 10010 3576 10015 3632
rect 8293 3571 8359 3574
rect 9949 3571 10015 3576
rect 10542 3572 10548 3636
rect 10612 3634 10618 3636
rect 10869 3634 10935 3637
rect 10612 3632 10935 3634
rect 10612 3576 10874 3632
rect 10930 3576 10935 3632
rect 10612 3574 10935 3576
rect 10612 3572 10618 3574
rect 10869 3571 10935 3574
rect 12750 3572 12756 3636
rect 12820 3634 12826 3636
rect 13169 3634 13235 3637
rect 13721 3634 13787 3637
rect 12820 3632 13235 3634
rect 12820 3576 13174 3632
rect 13230 3576 13235 3632
rect 12820 3574 13235 3576
rect 12820 3572 12826 3574
rect 13169 3571 13235 3574
rect 13310 3632 13787 3634
rect 13310 3576 13726 3632
rect 13782 3576 13787 3632
rect 13310 3574 13787 3576
rect 0 3408 480 3528
rect 2589 3498 2655 3501
rect 6361 3498 6427 3501
rect 2589 3496 6427 3498
rect 2589 3440 2594 3496
rect 2650 3440 6366 3496
rect 6422 3440 6427 3496
rect 2589 3438 6427 3440
rect 2589 3435 2655 3438
rect 6361 3435 6427 3438
rect 7097 3498 7163 3501
rect 10910 3498 10916 3500
rect 7097 3496 10916 3498
rect 7097 3440 7102 3496
rect 7158 3440 10916 3496
rect 7097 3438 10916 3440
rect 7097 3435 7163 3438
rect 10910 3436 10916 3438
rect 10980 3436 10986 3500
rect 12065 3498 12131 3501
rect 13310 3498 13370 3574
rect 13721 3571 13787 3574
rect 14038 3572 14044 3636
rect 14108 3634 14114 3636
rect 22001 3634 22067 3637
rect 14108 3632 22067 3634
rect 14108 3576 22006 3632
rect 22062 3576 22067 3632
rect 14108 3574 22067 3576
rect 14108 3572 14114 3574
rect 22001 3571 22067 3574
rect 12065 3496 13370 3498
rect 12065 3440 12070 3496
rect 12126 3440 13370 3496
rect 12065 3438 13370 3440
rect 12065 3435 12131 3438
rect 13670 3436 13676 3500
rect 13740 3498 13746 3500
rect 15745 3498 15811 3501
rect 13740 3496 15811 3498
rect 13740 3440 15750 3496
rect 15806 3440 15811 3496
rect 13740 3438 15811 3440
rect 13740 3436 13746 3438
rect 15745 3435 15811 3438
rect 16021 3498 16087 3501
rect 16614 3498 16620 3500
rect 16021 3496 16620 3498
rect 16021 3440 16026 3496
rect 16082 3440 16620 3496
rect 16021 3438 16620 3440
rect 16021 3435 16087 3438
rect 16614 3436 16620 3438
rect 16684 3498 16690 3500
rect 19885 3498 19951 3501
rect 16684 3496 19951 3498
rect 16684 3440 19890 3496
rect 19946 3440 19951 3496
rect 16684 3438 19951 3440
rect 16684 3436 16690 3438
rect 19885 3435 19951 3438
rect 6453 3362 6519 3365
rect 8293 3362 8359 3365
rect 6453 3360 8359 3362
rect 6453 3304 6458 3360
rect 6514 3304 8298 3360
rect 8354 3304 8359 3360
rect 6453 3302 8359 3304
rect 6453 3299 6519 3302
rect 8293 3299 8359 3302
rect 8569 3362 8635 3365
rect 12617 3362 12683 3365
rect 8569 3360 12683 3362
rect 8569 3304 8574 3360
rect 8630 3304 12622 3360
rect 12678 3304 12683 3360
rect 8569 3302 12683 3304
rect 8569 3299 8635 3302
rect 12617 3299 12683 3302
rect 15653 3362 15719 3365
rect 18689 3362 18755 3365
rect 15653 3360 18755 3362
rect 15653 3304 15658 3360
rect 15714 3304 18694 3360
rect 18750 3304 18755 3360
rect 15653 3302 18755 3304
rect 15653 3299 15719 3302
rect 18689 3299 18755 3302
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 1669 3226 1735 3229
rect 62 3224 1735 3226
rect 62 3168 1674 3224
rect 1730 3168 1735 3224
rect 62 3166 1735 3168
rect 62 2712 122 3166
rect 1669 3163 1735 3166
rect 7005 3226 7071 3229
rect 11605 3226 11671 3229
rect 7005 3224 11671 3226
rect 7005 3168 7010 3224
rect 7066 3168 11610 3224
rect 11666 3168 11671 3224
rect 7005 3166 11671 3168
rect 7005 3163 7071 3166
rect 11605 3163 11671 3166
rect 15653 3226 15719 3229
rect 15878 3226 15884 3228
rect 15653 3224 15884 3226
rect 15653 3168 15658 3224
rect 15714 3168 15884 3224
rect 15653 3166 15884 3168
rect 15653 3163 15719 3166
rect 15878 3164 15884 3166
rect 15948 3164 15954 3228
rect 606 3028 612 3092
rect 676 3090 682 3092
rect 2405 3090 2471 3093
rect 676 3088 2471 3090
rect 676 3032 2410 3088
rect 2466 3032 2471 3088
rect 676 3030 2471 3032
rect 676 3028 682 3030
rect 2405 3027 2471 3030
rect 3693 3090 3759 3093
rect 6494 3090 6500 3092
rect 3693 3088 6500 3090
rect 3693 3032 3698 3088
rect 3754 3032 6500 3088
rect 3693 3030 6500 3032
rect 3693 3027 3759 3030
rect 6494 3028 6500 3030
rect 6564 3028 6570 3092
rect 6729 3090 6795 3093
rect 6862 3090 6868 3092
rect 6729 3088 6868 3090
rect 6729 3032 6734 3088
rect 6790 3032 6868 3088
rect 6729 3030 6868 3032
rect 6729 3027 6795 3030
rect 6862 3028 6868 3030
rect 6932 3028 6938 3092
rect 7414 3028 7420 3092
rect 7484 3090 7490 3092
rect 9213 3090 9279 3093
rect 7484 3088 9279 3090
rect 7484 3032 9218 3088
rect 9274 3032 9279 3088
rect 7484 3030 9279 3032
rect 7484 3028 7490 3030
rect 9213 3027 9279 3030
rect 9622 3028 9628 3092
rect 9692 3090 9698 3092
rect 10685 3090 10751 3093
rect 9692 3088 10751 3090
rect 9692 3032 10690 3088
rect 10746 3032 10751 3088
rect 9692 3030 10751 3032
rect 9692 3028 9698 3030
rect 10685 3027 10751 3030
rect 12709 3090 12775 3093
rect 13670 3090 13676 3092
rect 12709 3088 13676 3090
rect 12709 3032 12714 3088
rect 12770 3032 13676 3088
rect 12709 3030 13676 3032
rect 12709 3027 12775 3030
rect 13670 3028 13676 3030
rect 13740 3028 13746 3092
rect 15009 3090 15075 3093
rect 13816 3088 15075 3090
rect 13816 3032 15014 3088
rect 15070 3032 15075 3088
rect 13816 3030 15075 3032
rect 2313 2954 2379 2957
rect 3366 2954 3372 2956
rect 2313 2952 3372 2954
rect 2313 2896 2318 2952
rect 2374 2896 3372 2952
rect 2313 2894 3372 2896
rect 2313 2891 2379 2894
rect 3366 2892 3372 2894
rect 3436 2954 3442 2956
rect 7005 2954 7071 2957
rect 3436 2952 7071 2954
rect 3436 2896 7010 2952
rect 7066 2896 7071 2952
rect 3436 2894 7071 2896
rect 3436 2892 3442 2894
rect 7005 2891 7071 2894
rect 8702 2892 8708 2956
rect 8772 2954 8778 2956
rect 8845 2954 8911 2957
rect 8772 2952 8911 2954
rect 8772 2896 8850 2952
rect 8906 2896 8911 2952
rect 8772 2894 8911 2896
rect 8772 2892 8778 2894
rect 8845 2891 8911 2894
rect 9029 2954 9095 2957
rect 9397 2954 9463 2957
rect 9029 2952 9463 2954
rect 9029 2896 9034 2952
rect 9090 2896 9402 2952
rect 9458 2896 9463 2952
rect 9029 2894 9463 2896
rect 9029 2891 9095 2894
rect 9397 2891 9463 2894
rect 10225 2954 10291 2957
rect 13816 2954 13876 3030
rect 15009 3027 15075 3030
rect 16113 3090 16179 3093
rect 19609 3090 19675 3093
rect 20069 3090 20135 3093
rect 23606 3090 23612 3092
rect 16113 3088 20135 3090
rect 16113 3032 16118 3088
rect 16174 3032 19614 3088
rect 19670 3032 20074 3088
rect 20130 3032 20135 3088
rect 16113 3030 20135 3032
rect 16113 3027 16179 3030
rect 19609 3027 19675 3030
rect 20069 3027 20135 3030
rect 23246 3030 23612 3090
rect 10225 2952 13876 2954
rect 10225 2896 10230 2952
rect 10286 2896 13876 2952
rect 10225 2894 13876 2896
rect 10225 2891 10291 2894
rect 14406 2892 14412 2956
rect 14476 2954 14482 2956
rect 17493 2954 17559 2957
rect 23246 2954 23306 3030
rect 23606 3028 23612 3030
rect 23676 3028 23682 3092
rect 14476 2952 23306 2954
rect 14476 2896 17498 2952
rect 17554 2896 23306 2952
rect 14476 2894 23306 2896
rect 14476 2892 14482 2894
rect 17493 2891 17559 2894
rect 5533 2818 5599 2821
rect 7557 2818 7623 2821
rect 8661 2818 8727 2821
rect 5533 2816 8727 2818
rect 5533 2760 5538 2816
rect 5594 2760 7562 2816
rect 7618 2760 8666 2816
rect 8722 2760 8727 2816
rect 5533 2758 8727 2760
rect 5533 2755 5599 2758
rect 7557 2755 7623 2758
rect 8661 2755 8727 2758
rect 11145 2818 11211 2821
rect 12198 2818 12204 2820
rect 11145 2816 12204 2818
rect 11145 2760 11150 2816
rect 11206 2760 12204 2816
rect 11145 2758 12204 2760
rect 11145 2755 11211 2758
rect 12198 2756 12204 2758
rect 12268 2756 12274 2820
rect 12566 2756 12572 2820
rect 12636 2818 12642 2820
rect 16021 2818 16087 2821
rect 12636 2816 16087 2818
rect 12636 2760 16026 2816
rect 16082 2760 16087 2816
rect 12636 2758 16087 2760
rect 12636 2756 12642 2758
rect 16021 2755 16087 2758
rect 18822 2756 18828 2820
rect 18892 2818 18898 2820
rect 22093 2818 22159 2821
rect 23520 2820 24000 2848
rect 23520 2818 23612 2820
rect 18892 2816 22159 2818
rect 18892 2760 22098 2816
rect 22154 2760 22159 2816
rect 18892 2758 22159 2760
rect 23484 2758 23612 2818
rect 18892 2756 18898 2758
rect 22093 2755 22159 2758
rect 23520 2756 23612 2758
rect 23676 2756 24000 2820
rect 8944 2752 9264 2753
rect 0 2592 480 2712
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 23520 2728 24000 2756
rect 16944 2687 17264 2688
rect 1342 2620 1348 2684
rect 1412 2682 1418 2684
rect 4061 2682 4127 2685
rect 1412 2680 4127 2682
rect 1412 2624 4066 2680
rect 4122 2624 4127 2680
rect 1412 2622 4127 2624
rect 1412 2620 1418 2622
rect 4061 2619 4127 2622
rect 7005 2682 7071 2685
rect 7598 2682 7604 2684
rect 7005 2680 7604 2682
rect 7005 2624 7010 2680
rect 7066 2624 7604 2680
rect 7005 2622 7604 2624
rect 7005 2619 7071 2622
rect 7598 2620 7604 2622
rect 7668 2620 7674 2684
rect 10041 2682 10107 2685
rect 11881 2682 11947 2685
rect 10041 2680 11947 2682
rect 10041 2624 10046 2680
rect 10102 2624 11886 2680
rect 11942 2624 11947 2680
rect 10041 2622 11947 2624
rect 10041 2619 10107 2622
rect 11881 2619 11947 2622
rect 17401 2682 17467 2685
rect 18873 2682 18939 2685
rect 17401 2680 18939 2682
rect 17401 2624 17406 2680
rect 17462 2624 18878 2680
rect 18934 2624 18939 2680
rect 17401 2622 18939 2624
rect 17401 2619 17467 2622
rect 18873 2619 18939 2622
rect 4797 2546 4863 2549
rect 12617 2546 12683 2549
rect 4797 2544 12683 2546
rect 4797 2488 4802 2544
rect 4858 2488 12622 2544
rect 12678 2488 12683 2544
rect 4797 2486 12683 2488
rect 4797 2483 4863 2486
rect 12617 2483 12683 2486
rect 12893 2546 12959 2549
rect 14457 2546 14523 2549
rect 12893 2544 14523 2546
rect 12893 2488 12898 2544
rect 12954 2488 14462 2544
rect 14518 2488 14523 2544
rect 12893 2486 14523 2488
rect 12893 2483 12959 2486
rect 14457 2483 14523 2486
rect 17217 2546 17283 2549
rect 17350 2546 17356 2548
rect 17217 2544 17356 2546
rect 17217 2488 17222 2544
rect 17278 2488 17356 2544
rect 17217 2486 17356 2488
rect 17217 2483 17283 2486
rect 17350 2484 17356 2486
rect 17420 2484 17426 2548
rect 3601 2410 3667 2413
rect 62 2408 3667 2410
rect 62 2352 3606 2408
rect 3662 2352 3667 2408
rect 62 2350 3667 2352
rect 62 1896 122 2350
rect 3601 2347 3667 2350
rect 6637 2410 6703 2413
rect 6637 2408 13830 2410
rect 6637 2352 6642 2408
rect 6698 2352 13830 2408
rect 6637 2350 13830 2352
rect 6637 2347 6703 2350
rect 6494 2212 6500 2276
rect 6564 2274 6570 2276
rect 12709 2274 12775 2277
rect 6564 2272 12775 2274
rect 6564 2216 12714 2272
rect 12770 2216 12775 2272
rect 6564 2214 12775 2216
rect 13770 2274 13830 2350
rect 14774 2348 14780 2412
rect 14844 2410 14850 2412
rect 21725 2410 21791 2413
rect 14844 2408 21791 2410
rect 14844 2352 21730 2408
rect 21786 2352 21791 2408
rect 14844 2350 21791 2352
rect 14844 2348 14850 2350
rect 21725 2347 21791 2350
rect 19885 2274 19951 2277
rect 13770 2272 19951 2274
rect 13770 2216 19890 2272
rect 19946 2216 19951 2272
rect 13770 2214 19951 2216
rect 6564 2212 6570 2214
rect 12709 2211 12775 2214
rect 19885 2211 19951 2214
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 4286 1940 4292 2004
rect 4356 2002 4362 2004
rect 9397 2002 9463 2005
rect 21725 2002 21791 2005
rect 23606 2002 23612 2004
rect 4356 2000 21791 2002
rect 4356 1944 9402 2000
rect 9458 1944 21730 2000
rect 21786 1944 21791 2000
rect 4356 1942 21791 1944
rect 4356 1940 4362 1942
rect 9397 1939 9463 1942
rect 21725 1939 21791 1942
rect 23246 1942 23612 2002
rect 0 1776 480 1896
rect 3141 1866 3207 1869
rect 12525 1866 12591 1869
rect 3141 1864 12591 1866
rect 3141 1808 3146 1864
rect 3202 1808 12530 1864
rect 12586 1808 12591 1864
rect 3141 1806 12591 1808
rect 3141 1803 3207 1806
rect 12525 1803 12591 1806
rect 14733 1866 14799 1869
rect 23246 1866 23306 1942
rect 23606 1940 23612 1942
rect 23676 1940 23682 2004
rect 14733 1864 23306 1866
rect 14733 1808 14738 1864
rect 14794 1808 23306 1864
rect 14733 1806 23306 1808
rect 14733 1803 14799 1806
rect 2313 1730 2379 1733
rect 12801 1730 12867 1733
rect 23520 1732 24000 1760
rect 23520 1730 23612 1732
rect 2313 1728 12867 1730
rect 2313 1672 2318 1728
rect 2374 1672 12806 1728
rect 12862 1672 12867 1728
rect 2313 1670 12867 1672
rect 23484 1670 23612 1730
rect 2313 1667 2379 1670
rect 12801 1667 12867 1670
rect 23520 1668 23612 1670
rect 23676 1668 24000 1732
rect 23520 1640 24000 1668
rect 565 1594 631 1597
rect 62 1592 631 1594
rect 62 1536 570 1592
rect 626 1536 631 1592
rect 62 1534 631 1536
rect 62 1080 122 1534
rect 565 1531 631 1534
rect 8477 1458 8543 1461
rect 18045 1458 18111 1461
rect 8477 1456 18111 1458
rect 8477 1400 8482 1456
rect 8538 1400 18050 1456
rect 18106 1400 18111 1456
rect 8477 1398 18111 1400
rect 8477 1395 8543 1398
rect 18045 1395 18111 1398
rect 11421 1322 11487 1325
rect 20713 1322 20779 1325
rect 11421 1320 20779 1322
rect 11421 1264 11426 1320
rect 11482 1264 20718 1320
rect 20774 1264 20779 1320
rect 11421 1262 20779 1264
rect 11421 1259 11487 1262
rect 20713 1259 20779 1262
rect 3325 1186 3391 1189
rect 19333 1186 19399 1189
rect 3325 1184 19399 1186
rect 3325 1128 3330 1184
rect 3386 1128 19338 1184
rect 19394 1128 19399 1184
rect 3325 1126 19399 1128
rect 3325 1123 3391 1126
rect 19333 1123 19399 1126
rect 19558 1124 19564 1188
rect 19628 1186 19634 1188
rect 19628 1126 23674 1186
rect 19628 1124 19634 1126
rect 0 960 480 1080
rect 6361 1050 6427 1053
rect 12382 1050 12388 1052
rect 6361 1048 12388 1050
rect 6361 992 6366 1048
rect 6422 992 12388 1048
rect 6361 990 12388 992
rect 6361 987 6427 990
rect 12382 988 12388 990
rect 12452 988 12458 1052
rect 6913 914 6979 917
rect 16389 914 16455 917
rect 6913 912 16455 914
rect 6913 856 6918 912
rect 6974 856 16394 912
rect 16450 856 16455 912
rect 6913 854 16455 856
rect 6913 851 6979 854
rect 16389 851 16455 854
rect 5625 778 5691 781
rect 62 776 5691 778
rect 62 720 5630 776
rect 5686 720 5691 776
rect 62 718 5691 720
rect 62 400 122 718
rect 5625 715 5691 718
rect 8753 778 8819 781
rect 20253 778 20319 781
rect 8753 776 20319 778
rect 8753 720 8758 776
rect 8814 720 20258 776
rect 20314 720 20319 776
rect 8753 718 20319 720
rect 8753 715 8819 718
rect 20253 715 20319 718
rect 23614 672 23674 1126
rect 11697 642 11763 645
rect 20345 642 20411 645
rect 11697 640 20411 642
rect 11697 584 11702 640
rect 11758 584 20350 640
rect 20406 584 20411 640
rect 11697 582 20411 584
rect 11697 579 11763 582
rect 20345 579 20411 582
rect 23520 552 24000 672
rect 8109 506 8175 509
rect 19701 506 19767 509
rect 8109 504 19767 506
rect 8109 448 8114 504
rect 8170 448 19706 504
rect 19762 448 19767 504
rect 8109 446 19767 448
rect 8109 443 8175 446
rect 19701 443 19767 446
rect 0 280 480 400
rect 7741 370 7807 373
rect 22277 370 22343 373
rect 7741 368 22343 370
rect 7741 312 7746 368
rect 7802 312 22282 368
rect 22338 312 22343 368
rect 7741 310 22343 312
rect 7741 307 7807 310
rect 22277 307 22343 310
rect 4613 232 4679 237
rect 4613 176 4618 232
rect 4674 176 4679 232
rect 4613 171 4679 176
rect 6821 234 6887 237
rect 14089 234 14155 237
rect 6821 232 14155 234
rect 6821 176 6826 232
rect 6882 176 14094 232
rect 14150 176 14155 232
rect 6821 174 14155 176
rect 6821 171 6887 174
rect 14089 171 14155 174
rect 289 98 355 101
rect 422 98 428 100
rect 289 96 428 98
rect 289 40 294 96
rect 350 40 428 96
rect 289 38 428 40
rect 289 35 355 38
rect 422 36 428 38
rect 492 36 498 100
rect 4616 98 4676 171
rect 14917 98 14983 101
rect 4616 96 14983 98
rect 4616 40 14922 96
rect 14978 40 14983 96
rect 4616 38 14983 40
rect 14917 35 14983 38
rect 20662 36 20668 100
rect 20732 98 20738 100
rect 21449 98 21515 101
rect 20732 96 21515 98
rect 20732 40 21454 96
rect 21510 40 21515 96
rect 20732 38 21515 40
rect 20732 36 20738 38
rect 21449 35 21515 38
<< via3 >>
rect 3556 23020 3620 23084
rect 2820 22884 2884 22948
rect 7972 22748 8036 22812
rect 17908 22612 17972 22676
rect 3924 22476 3988 22540
rect 15700 22340 15764 22404
rect 1900 22204 1964 22268
rect 12388 22204 12452 22268
rect 4660 22068 4724 22132
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 10548 21524 10612 21588
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 3188 20980 3252 21044
rect 4108 20980 4172 21044
rect 9812 20980 9876 21044
rect 9628 20878 9692 20942
rect 244 20708 308 20772
rect 10180 20708 10244 20772
rect 12756 20708 12820 20772
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 3372 20436 3436 20500
rect 8708 20300 8772 20364
rect 7052 20164 7116 20228
rect 19564 20164 19628 20228
rect 23612 20164 23676 20228
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 9444 20028 9508 20092
rect 244 19756 308 19820
rect 7420 19756 7484 19820
rect 2084 19484 2148 19548
rect 3556 19212 3620 19276
rect 5764 19620 5828 19684
rect 8156 19620 8220 19684
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 5396 19484 5460 19548
rect 6868 19348 6932 19412
rect 17356 19484 17420 19548
rect 13676 19348 13740 19412
rect 1164 19076 1228 19140
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 7604 18940 7668 19004
rect 14044 18940 14108 19004
rect 4108 18804 4172 18868
rect 1532 18532 1596 18596
rect 6500 18668 6564 18732
rect 14596 18668 14660 18732
rect 10180 18532 10244 18596
rect 12756 18532 12820 18596
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 6316 18396 6380 18460
rect 8340 18396 8404 18460
rect 19932 18396 19996 18460
rect 612 18260 676 18324
rect 8708 18260 8772 18324
rect 3740 18124 3804 18188
rect 980 17988 1044 18052
rect 8524 17988 8588 18052
rect 15332 17988 15396 18052
rect 15884 17988 15948 18052
rect 17540 17988 17604 18052
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 60 17852 124 17916
rect 1348 17852 1412 17916
rect 14228 17852 14292 17916
rect 2820 17716 2884 17780
rect 8708 17716 8772 17780
rect 3004 17580 3068 17644
rect 4660 17580 4724 17644
rect 9628 17580 9692 17644
rect 796 17444 860 17508
rect 796 17308 860 17372
rect 5764 17444 5828 17508
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 7604 17308 7668 17372
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 9444 17308 9508 17372
rect 11652 17172 11716 17236
rect 1716 16900 1780 16964
rect 3556 16900 3620 16964
rect 4476 16900 4540 16964
rect 5396 16900 5460 16964
rect 7236 16900 7300 16964
rect 14964 16900 15028 16964
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 60 16628 124 16692
rect 4292 16764 4356 16828
rect 11836 16628 11900 16692
rect 6684 16492 6748 16556
rect 7788 16492 7852 16556
rect 13676 16492 13740 16556
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 3924 16220 3988 16284
rect 7604 16220 7668 16284
rect 11468 16220 11532 16284
rect 4108 15812 4172 15876
rect 5948 15812 6012 15876
rect 2268 15540 2332 15604
rect 14412 15948 14476 16012
rect 12756 15812 12820 15876
rect 17356 15812 17420 15876
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 11100 15540 11164 15604
rect 3924 15404 3988 15468
rect 7788 15404 7852 15468
rect 11284 15404 11348 15468
rect 18460 15404 18524 15468
rect 19932 15404 19996 15468
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 2084 15132 2148 15196
rect 3372 15132 3436 15196
rect 12572 15132 12636 15196
rect 16068 15132 16132 15196
rect 17724 15132 17788 15196
rect 10732 14996 10796 15060
rect 2084 14860 2148 14924
rect 12020 14860 12084 14924
rect 3372 14784 3436 14788
rect 3372 14728 3386 14784
rect 3386 14728 3436 14784
rect 3372 14724 3436 14728
rect 6132 14588 6196 14652
rect 13492 14724 13556 14788
rect 15516 14724 15580 14788
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 8340 14588 8404 14652
rect 7420 14452 7484 14516
rect 15148 14452 15212 14516
rect 2452 14180 2516 14244
rect 3188 14180 3252 14244
rect 3556 14180 3620 14244
rect 4476 14180 4540 14244
rect 10548 14180 10612 14244
rect 16252 14180 16316 14244
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 2636 14044 2700 14108
rect 6868 14044 6932 14108
rect 12204 14044 12268 14108
rect 16620 14180 16684 14244
rect 19196 14180 19260 14244
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 16620 14044 16684 14108
rect 6500 13908 6564 13972
rect 60 13772 124 13836
rect 7236 13908 7300 13972
rect 7420 13772 7484 13836
rect 10180 13908 10244 13972
rect 12388 13908 12452 13972
rect 14044 13908 14108 13972
rect 60 13636 124 13700
rect 3740 13636 3804 13700
rect 4476 13636 4540 13700
rect 4660 13636 4724 13700
rect 5948 13636 6012 13700
rect 6316 13636 6380 13700
rect 15884 13636 15948 13700
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 3740 13500 3804 13564
rect 4660 13500 4724 13564
rect 7236 13500 7300 13564
rect 7604 13500 7668 13564
rect 8340 13500 8404 13564
rect 1348 13228 1412 13292
rect 3188 13228 3252 13292
rect 7604 13364 7668 13428
rect 14780 13500 14844 13564
rect 18092 13500 18156 13564
rect 17908 13364 17972 13428
rect 8524 13228 8588 13292
rect 9996 13228 10060 13292
rect 15884 13228 15948 13292
rect 20116 13228 20180 13292
rect 10548 13092 10612 13156
rect 15516 13092 15580 13156
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 5580 12956 5644 13020
rect 244 12820 308 12884
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 10180 12956 10244 13020
rect 2820 12684 2884 12748
rect 4108 12684 4172 12748
rect 8340 12684 8404 12748
rect 8708 12684 8772 12748
rect 9996 12684 10060 12748
rect 16804 12684 16868 12748
rect 2820 12548 2884 12612
rect 9628 12548 9692 12612
rect 14964 12548 15028 12612
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 60 12276 124 12340
rect 1348 12276 1412 12340
rect 3556 12276 3620 12340
rect 12572 12412 12636 12476
rect 14596 12412 14660 12476
rect 16068 12412 16132 12476
rect 6868 12276 6932 12340
rect 7972 12276 8036 12340
rect 10364 12276 10428 12340
rect 18460 12276 18524 12340
rect 20668 12276 20732 12340
rect 60 12004 124 12068
rect 3924 12004 3988 12068
rect 4108 12004 4172 12068
rect 7972 12004 8036 12068
rect 8524 12004 8588 12068
rect 9444 12004 9508 12068
rect 10180 12004 10244 12068
rect 10916 12004 10980 12068
rect 12572 12004 12636 12068
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 3556 11868 3620 11932
rect 12756 11868 12820 11932
rect 10732 11732 10796 11796
rect 12572 11596 12636 11660
rect 15700 11596 15764 11660
rect 2636 11460 2700 11524
rect 5396 11460 5460 11524
rect 15148 11460 15212 11524
rect 18828 11460 18892 11524
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 1532 11324 1596 11388
rect 5396 11324 5460 11388
rect 7236 11324 7300 11388
rect 8340 11324 8404 11388
rect 1532 11188 1596 11252
rect 3556 11188 3620 11252
rect 11468 11188 11532 11252
rect 12388 11188 12452 11252
rect 18644 11188 18708 11252
rect 60 10916 124 10980
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 11284 11052 11348 11116
rect 10180 10916 10244 10980
rect 15148 10916 15212 10980
rect 23612 10916 23676 10980
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 60 10644 124 10708
rect 8340 10780 8404 10844
rect 13676 10780 13740 10844
rect 4292 10644 4356 10708
rect 12756 10644 12820 10708
rect 3372 10508 3436 10572
rect 4292 10508 4356 10572
rect 1716 10372 1780 10436
rect 7236 10372 7300 10436
rect 7604 10508 7668 10572
rect 18644 10508 18708 10572
rect 11284 10372 11348 10436
rect 19564 10372 19628 10436
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 1716 10236 1780 10300
rect 4108 10236 4172 10300
rect 7236 10236 7300 10300
rect 12572 10236 12636 10300
rect 14228 10236 14292 10300
rect 17724 10236 17788 10300
rect 21956 10236 22020 10300
rect 15332 10100 15396 10164
rect 3740 9828 3804 9892
rect 4292 9964 4356 10028
rect 6684 9964 6748 10028
rect 8340 9964 8404 10028
rect 11100 9964 11164 10028
rect 11652 9964 11716 10028
rect 3740 9692 3804 9756
rect 8708 9828 8772 9892
rect 9444 9828 9508 9892
rect 10916 9828 10980 9892
rect 11468 9828 11532 9892
rect 20300 9964 20364 10028
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 3372 9420 3436 9484
rect 5396 9692 5460 9756
rect 7604 9692 7668 9756
rect 9628 9692 9692 9756
rect 4660 9556 4724 9620
rect 8708 9556 8772 9620
rect 21588 9828 21652 9892
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 14412 9692 14476 9756
rect 20300 9692 20364 9756
rect 10916 9420 10980 9484
rect 12204 9284 12268 9348
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 980 9148 1044 9212
rect 1900 9148 1964 9212
rect 3740 9148 3804 9212
rect 4660 9148 4724 9212
rect 5396 9148 5460 9212
rect 11652 9148 11716 9212
rect 18276 9148 18340 9212
rect 19380 9148 19444 9212
rect 1532 8876 1596 8940
rect 3740 8876 3804 8940
rect 5580 9012 5644 9076
rect 10364 9012 10428 9076
rect 7052 8876 7116 8940
rect 7788 8876 7852 8940
rect 8708 8876 8772 8940
rect 10364 8876 10428 8940
rect 19932 9012 19996 9076
rect 12204 8876 12268 8940
rect 2084 8740 2148 8804
rect 3004 8740 3068 8804
rect 4108 8740 4172 8804
rect 11284 8740 11348 8804
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 3556 8604 3620 8668
rect 13676 8876 13740 8940
rect 14412 8876 14476 8940
rect 16252 8876 16316 8940
rect 19564 8876 19628 8940
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 2268 8332 2332 8396
rect 3004 8196 3068 8260
rect 4660 8196 4724 8260
rect 13860 8468 13924 8532
rect 10548 8332 10612 8396
rect 11836 8196 11900 8260
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 10364 8060 10428 8124
rect 11468 8060 11532 8124
rect 11836 8060 11900 8124
rect 3556 7788 3620 7852
rect 5764 7788 5828 7852
rect 6684 7788 6748 7852
rect 6868 7788 6932 7852
rect 5764 7652 5828 7716
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 3004 7516 3068 7580
rect 12020 7516 12084 7580
rect 9812 7380 9876 7444
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 13492 7516 13556 7580
rect 18460 7516 18524 7580
rect 2636 7108 2700 7172
rect 4292 7108 4356 7172
rect 6132 7108 6196 7172
rect 6684 7108 6748 7172
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 7788 6700 7852 6764
rect 6132 6564 6196 6628
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 2084 6428 2148 6492
rect 2820 6428 2884 6492
rect 20668 6488 20732 6492
rect 20668 6432 20718 6488
rect 20718 6432 20732 6488
rect 20668 6428 20732 6432
rect 19932 6292 19996 6356
rect 3188 6156 3252 6220
rect 4108 6156 4172 6220
rect 4292 6156 4356 6220
rect 5948 6156 6012 6220
rect 7604 6156 7668 6220
rect 17540 6156 17604 6220
rect 1716 6020 1780 6084
rect 16804 6020 16868 6084
rect 18828 6020 18892 6084
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 1348 5884 1412 5948
rect 18092 5884 18156 5948
rect 4476 5748 4540 5812
rect 9996 5748 10060 5812
rect 4476 5476 4540 5540
rect 5580 5476 5644 5540
rect 10732 5476 10796 5540
rect 11100 5476 11164 5540
rect 11652 5476 11716 5540
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 12388 5340 12452 5404
rect 14044 5068 14108 5132
rect 15148 5068 15212 5132
rect 19748 5068 19812 5132
rect 20668 5068 20732 5132
rect 1900 4932 1964 4996
rect 8156 4932 8220 4996
rect 9996 4932 10060 4996
rect 11836 4932 11900 4996
rect 12572 4932 12636 4996
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 244 4796 308 4860
rect 5764 4796 5828 4860
rect 6500 4796 6564 4860
rect 7972 4796 8036 4860
rect 9812 4796 9876 4860
rect 10180 4796 10244 4860
rect 20116 4796 20180 4860
rect 3740 4660 3804 4724
rect 19932 4660 19996 4724
rect 12572 4524 12636 4588
rect 9996 4388 10060 4452
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 796 4252 860 4316
rect 6316 4252 6380 4316
rect 7236 4252 7300 4316
rect 8340 4252 8404 4316
rect 8524 4252 8588 4316
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 6684 4116 6748 4180
rect 9444 4116 9508 4180
rect 10732 4252 10796 4316
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 4108 3844 4172 3908
rect 7052 3844 7116 3908
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 6132 3708 6196 3772
rect 6500 3708 6564 3772
rect 7972 3708 8036 3772
rect 2452 3572 2516 3636
rect 3924 3572 3988 3636
rect 5580 3572 5644 3636
rect 10364 3980 10428 4044
rect 18460 3844 18524 3908
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 10548 3572 10612 3636
rect 12756 3572 12820 3636
rect 10916 3436 10980 3500
rect 14044 3572 14108 3636
rect 13676 3436 13740 3500
rect 16620 3436 16684 3500
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 15884 3164 15948 3228
rect 612 3028 676 3092
rect 6500 3028 6564 3092
rect 6868 3028 6932 3092
rect 7420 3028 7484 3092
rect 9628 3028 9692 3092
rect 13676 3028 13740 3092
rect 3372 2892 3436 2956
rect 8708 2892 8772 2956
rect 14412 2892 14476 2956
rect 23612 3028 23676 3092
rect 12204 2756 12268 2820
rect 12572 2756 12636 2820
rect 18828 2756 18892 2820
rect 23612 2756 23676 2820
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 1348 2620 1412 2684
rect 7604 2620 7668 2684
rect 17356 2484 17420 2548
rect 6500 2212 6564 2276
rect 14780 2348 14844 2412
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 4292 1940 4356 2004
rect 23612 1940 23676 2004
rect 23612 1668 23676 1732
rect 19564 1124 19628 1188
rect 12388 988 12452 1052
rect 428 36 492 100
rect 20668 36 20732 100
<< metal4 >>
rect 3555 23084 3621 23085
rect 3555 23020 3556 23084
rect 3620 23020 3621 23084
rect 3555 23019 3621 23020
rect 2819 22948 2885 22949
rect 2819 22884 2820 22948
rect 2884 22884 2885 22948
rect 2819 22883 2885 22884
rect 1899 22268 1965 22269
rect 1899 22204 1900 22268
rect 1964 22204 1965 22268
rect 1899 22203 1965 22204
rect 243 20772 309 20773
rect 243 20770 244 20772
rect 62 20710 244 20770
rect 62 17917 122 20710
rect 243 20708 244 20710
rect 308 20708 309 20772
rect 243 20707 309 20708
rect 243 19820 309 19821
rect 243 19756 244 19820
rect 308 19756 309 19820
rect 243 19755 309 19756
rect 59 17916 125 17917
rect 59 17852 60 17916
rect 124 17852 125 17916
rect 59 17851 125 17852
rect 59 16692 125 16693
rect 59 16628 60 16692
rect 124 16628 125 16692
rect 59 16627 125 16628
rect 62 13837 122 16627
rect 59 13836 125 13837
rect 59 13772 60 13836
rect 124 13772 125 13836
rect 59 13771 125 13772
rect 62 13701 122 13771
rect 59 13700 125 13701
rect 59 13636 60 13700
rect 124 13636 125 13700
rect 59 13635 125 13636
rect 62 12746 122 13635
rect 246 12885 306 19755
rect 243 12884 309 12885
rect 243 12820 244 12884
rect 308 12820 309 12884
rect 243 12819 309 12820
rect 62 12686 306 12746
rect 59 12340 125 12341
rect 59 12276 60 12340
rect 124 12276 125 12340
rect 59 12275 125 12276
rect 62 12069 122 12275
rect 59 12068 125 12069
rect 59 12004 60 12068
rect 124 12004 125 12068
rect 59 12003 125 12004
rect 59 10980 125 10981
rect 59 10916 60 10980
rect 124 10916 125 10980
rect 59 10915 125 10916
rect 62 10709 122 10915
rect 59 10708 125 10709
rect 59 10644 60 10708
rect 124 10644 125 10708
rect 59 10643 125 10644
rect 246 4861 306 12686
rect 243 4860 309 4861
rect 243 4796 244 4860
rect 308 4796 309 4860
rect 243 4795 309 4796
rect 430 101 490 19942
rect 1163 19140 1229 19141
rect 1163 19076 1164 19140
rect 1228 19076 1229 19140
rect 1163 19075 1229 19076
rect 611 18324 677 18325
rect 611 18260 612 18324
rect 676 18260 677 18324
rect 611 18259 677 18260
rect 614 3093 674 18259
rect 798 17509 858 18582
rect 979 18052 1045 18053
rect 979 17988 980 18052
rect 1044 17988 1045 18052
rect 979 17987 1045 17988
rect 795 17508 861 17509
rect 795 17444 796 17508
rect 860 17444 861 17508
rect 795 17443 861 17444
rect 795 17372 861 17373
rect 795 17308 796 17372
rect 860 17308 861 17372
rect 795 17307 861 17308
rect 798 4317 858 17307
rect 982 9213 1042 17987
rect 979 9212 1045 9213
rect 979 9148 980 9212
rect 1044 9148 1045 9212
rect 979 9147 1045 9148
rect 795 4316 861 4317
rect 795 4252 796 4316
rect 860 4252 861 4316
rect 795 4251 861 4252
rect 1166 4170 1226 19075
rect 1531 18596 1597 18597
rect 1531 18532 1532 18596
rect 1596 18532 1597 18596
rect 1531 18531 1597 18532
rect 1347 17916 1413 17917
rect 1347 17852 1348 17916
rect 1412 17852 1413 17916
rect 1347 17851 1413 17852
rect 1350 13293 1410 17851
rect 1347 13292 1413 13293
rect 1347 13228 1348 13292
rect 1412 13228 1413 13292
rect 1347 13227 1413 13228
rect 1347 12340 1413 12341
rect 1347 12276 1348 12340
rect 1412 12276 1413 12340
rect 1347 12275 1413 12276
rect 1350 5949 1410 12275
rect 1534 11389 1594 18531
rect 1715 16964 1781 16965
rect 1715 16900 1716 16964
rect 1780 16900 1781 16964
rect 1715 16899 1781 16900
rect 1531 11388 1597 11389
rect 1531 11324 1532 11388
rect 1596 11324 1597 11388
rect 1531 11323 1597 11324
rect 1531 11252 1597 11253
rect 1531 11188 1532 11252
rect 1596 11188 1597 11252
rect 1531 11187 1597 11188
rect 1534 8941 1594 11187
rect 1718 10437 1778 16899
rect 1715 10436 1781 10437
rect 1715 10372 1716 10436
rect 1780 10372 1781 10436
rect 1715 10371 1781 10372
rect 1715 10300 1781 10301
rect 1715 10236 1716 10300
rect 1780 10236 1781 10300
rect 1715 10235 1781 10236
rect 1531 8940 1597 8941
rect 1531 8876 1532 8940
rect 1596 8876 1597 8940
rect 1531 8875 1597 8876
rect 1718 6085 1778 10235
rect 1902 9213 1962 22203
rect 2083 19548 2149 19549
rect 2083 19484 2084 19548
rect 2148 19484 2149 19548
rect 2083 19483 2149 19484
rect 2086 15197 2146 19483
rect 2267 15604 2333 15605
rect 2267 15540 2268 15604
rect 2332 15540 2333 15604
rect 2267 15539 2333 15540
rect 2083 15196 2149 15197
rect 2083 15132 2084 15196
rect 2148 15132 2149 15196
rect 2083 15131 2149 15132
rect 2083 14924 2149 14925
rect 2083 14860 2084 14924
rect 2148 14860 2149 14924
rect 2083 14859 2149 14860
rect 1899 9212 1965 9213
rect 1899 9148 1900 9212
rect 1964 9148 1965 9212
rect 1899 9147 1965 9148
rect 2086 9074 2146 14859
rect 1902 9014 2146 9074
rect 1715 6084 1781 6085
rect 1715 6020 1716 6084
rect 1780 6020 1781 6084
rect 1715 6019 1781 6020
rect 1347 5948 1413 5949
rect 1347 5884 1348 5948
rect 1412 5884 1413 5948
rect 1347 5883 1413 5884
rect 1902 4997 1962 9014
rect 2083 8804 2149 8805
rect 2083 8740 2084 8804
rect 2148 8740 2149 8804
rect 2083 8739 2149 8740
rect 2086 6493 2146 8739
rect 2270 8397 2330 15539
rect 2454 14245 2514 19262
rect 2822 18730 2882 22883
rect 3187 21044 3253 21045
rect 3187 20980 3188 21044
rect 3252 20980 3253 21044
rect 3187 20979 3253 20980
rect 2638 18670 2882 18730
rect 2451 14244 2517 14245
rect 2451 14180 2452 14244
rect 2516 14180 2517 14244
rect 2451 14179 2517 14180
rect 2267 8396 2333 8397
rect 2267 8332 2268 8396
rect 2332 8332 2333 8396
rect 2267 8331 2333 8332
rect 2083 6492 2149 6493
rect 2083 6428 2084 6492
rect 2148 6428 2149 6492
rect 2083 6427 2149 6428
rect 1899 4996 1965 4997
rect 1899 4932 1900 4996
rect 1964 4932 1965 4996
rect 1899 4931 1965 4932
rect 1166 4110 1410 4170
rect 611 3092 677 3093
rect 611 3028 612 3092
rect 676 3028 677 3092
rect 611 3027 677 3028
rect 1350 2685 1410 4110
rect 2454 3637 2514 14179
rect 2638 14109 2698 18670
rect 2819 17780 2885 17781
rect 2819 17716 2820 17780
rect 2884 17716 2885 17780
rect 2819 17715 2885 17716
rect 2635 14108 2701 14109
rect 2635 14044 2636 14108
rect 2700 14044 2701 14108
rect 2635 14043 2701 14044
rect 2822 12749 2882 17715
rect 3003 17644 3069 17645
rect 3003 17580 3004 17644
rect 3068 17580 3069 17644
rect 3003 17579 3069 17580
rect 2819 12748 2885 12749
rect 2819 12684 2820 12748
rect 2884 12684 2885 12748
rect 2819 12683 2885 12684
rect 2819 12612 2885 12613
rect 2819 12548 2820 12612
rect 2884 12548 2885 12612
rect 2819 12547 2885 12548
rect 2635 11524 2701 11525
rect 2635 11460 2636 11524
rect 2700 11460 2701 11524
rect 2635 11459 2701 11460
rect 2638 7173 2698 11459
rect 2635 7172 2701 7173
rect 2635 7108 2636 7172
rect 2700 7108 2701 7172
rect 2635 7107 2701 7108
rect 2822 6493 2882 12547
rect 3006 8805 3066 17579
rect 3190 14245 3250 20979
rect 3371 20500 3437 20501
rect 3371 20436 3372 20500
rect 3436 20436 3437 20500
rect 3371 20435 3437 20436
rect 3374 15197 3434 20435
rect 3558 19277 3618 23019
rect 7971 22812 8037 22813
rect 7971 22748 7972 22812
rect 8036 22748 8037 22812
rect 7971 22747 8037 22748
rect 3923 22540 3989 22541
rect 3923 22476 3924 22540
rect 3988 22476 3989 22540
rect 3923 22475 3989 22476
rect 3555 19276 3621 19277
rect 3555 19212 3556 19276
rect 3620 19212 3621 19276
rect 3555 19211 3621 19212
rect 3558 16965 3618 19211
rect 3739 18188 3805 18189
rect 3739 18124 3740 18188
rect 3804 18124 3805 18188
rect 3739 18123 3805 18124
rect 3555 16964 3621 16965
rect 3555 16900 3556 16964
rect 3620 16900 3621 16964
rect 3555 16899 3621 16900
rect 3371 15196 3437 15197
rect 3371 15132 3372 15196
rect 3436 15132 3437 15196
rect 3371 15131 3437 15132
rect 3371 14788 3437 14789
rect 3371 14724 3372 14788
rect 3436 14724 3437 14788
rect 3371 14723 3437 14724
rect 3187 14244 3253 14245
rect 3187 14180 3188 14244
rect 3252 14180 3253 14244
rect 3187 14179 3253 14180
rect 3187 13292 3253 13293
rect 3187 13228 3188 13292
rect 3252 13228 3253 13292
rect 3187 13227 3253 13228
rect 3003 8804 3069 8805
rect 3003 8740 3004 8804
rect 3068 8740 3069 8804
rect 3003 8739 3069 8740
rect 3003 8260 3069 8261
rect 3003 8196 3004 8260
rect 3068 8196 3069 8260
rect 3003 8195 3069 8196
rect 3006 7581 3066 8195
rect 3003 7580 3069 7581
rect 3003 7516 3004 7580
rect 3068 7516 3069 7580
rect 3003 7515 3069 7516
rect 2819 6492 2885 6493
rect 2819 6428 2820 6492
rect 2884 6428 2885 6492
rect 2819 6427 2885 6428
rect 3190 6221 3250 13227
rect 3374 10573 3434 14723
rect 3555 14244 3621 14245
rect 3555 14180 3556 14244
rect 3620 14180 3621 14244
rect 3555 14179 3621 14180
rect 3558 12341 3618 14179
rect 3742 13701 3802 18123
rect 3926 16285 3986 22475
rect 4659 22132 4725 22133
rect 4659 22068 4660 22132
rect 4724 22068 4725 22132
rect 4659 22067 4725 22068
rect 4107 21044 4173 21045
rect 4107 20980 4108 21044
rect 4172 20980 4173 21044
rect 4107 20979 4173 20980
rect 4110 18869 4170 20979
rect 4107 18868 4173 18869
rect 4107 18804 4108 18868
rect 4172 18804 4173 18868
rect 4107 18803 4173 18804
rect 4662 17645 4722 22067
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 7051 20228 7117 20229
rect 7051 20164 7052 20228
rect 7116 20164 7117 20228
rect 7051 20163 7117 20164
rect 5763 19684 5829 19685
rect 5763 19620 5764 19684
rect 5828 19620 5829 19684
rect 5763 19619 5829 19620
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 5395 19548 5461 19549
rect 5395 19484 5396 19548
rect 5460 19484 5461 19548
rect 5395 19483 5461 19484
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4659 17644 4725 17645
rect 4659 17580 4660 17644
rect 4724 17580 4725 17644
rect 4659 17579 4725 17580
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4475 16964 4541 16965
rect 4475 16900 4476 16964
rect 4540 16900 4541 16964
rect 4475 16899 4541 16900
rect 4291 16828 4357 16829
rect 4291 16764 4292 16828
rect 4356 16764 4357 16828
rect 4291 16763 4357 16764
rect 3923 16284 3989 16285
rect 3923 16220 3924 16284
rect 3988 16220 3989 16284
rect 3923 16219 3989 16220
rect 4107 15876 4173 15877
rect 4107 15812 4108 15876
rect 4172 15812 4173 15876
rect 4107 15811 4173 15812
rect 3923 15468 3989 15469
rect 3923 15404 3924 15468
rect 3988 15404 3989 15468
rect 3923 15403 3989 15404
rect 3739 13700 3805 13701
rect 3739 13636 3740 13700
rect 3804 13636 3805 13700
rect 3739 13635 3805 13636
rect 3739 13564 3805 13565
rect 3739 13500 3740 13564
rect 3804 13500 3805 13564
rect 3739 13499 3805 13500
rect 3555 12340 3621 12341
rect 3555 12276 3556 12340
rect 3620 12276 3621 12340
rect 3555 12275 3621 12276
rect 3555 11932 3621 11933
rect 3555 11868 3556 11932
rect 3620 11868 3621 11932
rect 3555 11867 3621 11868
rect 3558 11253 3618 11867
rect 3555 11252 3621 11253
rect 3555 11188 3556 11252
rect 3620 11188 3621 11252
rect 3555 11187 3621 11188
rect 3371 10572 3437 10573
rect 3371 10508 3372 10572
rect 3436 10508 3437 10572
rect 3371 10507 3437 10508
rect 3371 9484 3437 9485
rect 3371 9420 3372 9484
rect 3436 9420 3437 9484
rect 3371 9419 3437 9420
rect 3187 6220 3253 6221
rect 3187 6156 3188 6220
rect 3252 6156 3253 6220
rect 3187 6155 3253 6156
rect 2451 3636 2517 3637
rect 2451 3572 2452 3636
rect 2516 3572 2517 3636
rect 2451 3571 2517 3572
rect 3374 2957 3434 9419
rect 3558 8669 3618 11187
rect 3742 10026 3802 13499
rect 3926 12069 3986 15403
rect 4110 12749 4170 15811
rect 4107 12748 4173 12749
rect 4107 12684 4108 12748
rect 4172 12684 4173 12748
rect 4107 12683 4173 12684
rect 3923 12068 3989 12069
rect 3923 12004 3924 12068
rect 3988 12004 3989 12068
rect 3923 12003 3989 12004
rect 4107 12068 4173 12069
rect 4107 12004 4108 12068
rect 4172 12004 4173 12068
rect 4107 12003 4173 12004
rect 4110 10301 4170 12003
rect 4294 10709 4354 16763
rect 4478 14922 4538 16899
rect 4432 14862 4538 14922
rect 4944 16352 5264 17376
rect 5398 17234 5458 19483
rect 5766 17509 5826 19619
rect 6867 19412 6933 19413
rect 6867 19348 6868 19412
rect 6932 19348 6933 19412
rect 6867 19347 6933 19348
rect 6499 18732 6565 18733
rect 6499 18668 6500 18732
rect 6564 18668 6565 18732
rect 6499 18667 6565 18668
rect 6315 18460 6381 18461
rect 6315 18396 6316 18460
rect 6380 18396 6381 18460
rect 6315 18395 6381 18396
rect 5763 17508 5829 17509
rect 5763 17444 5764 17508
rect 5828 17444 5829 17508
rect 5763 17443 5829 17444
rect 5398 17174 5826 17234
rect 5395 16964 5461 16965
rect 5395 16900 5396 16964
rect 5460 16900 5461 16964
rect 5395 16899 5461 16900
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4432 14245 4492 14862
rect 4432 14244 4541 14245
rect 4432 14182 4476 14244
rect 4475 14180 4476 14182
rect 4540 14180 4541 14244
rect 4475 14179 4541 14180
rect 4662 13701 4722 14502
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4475 13700 4541 13701
rect 4475 13636 4476 13700
rect 4540 13636 4541 13700
rect 4475 13635 4541 13636
rect 4659 13700 4725 13701
rect 4659 13636 4660 13700
rect 4724 13636 4725 13700
rect 4659 13635 4725 13636
rect 4291 10708 4357 10709
rect 4291 10644 4292 10708
rect 4356 10644 4357 10708
rect 4291 10643 4357 10644
rect 4291 10572 4357 10573
rect 4291 10508 4292 10572
rect 4356 10508 4357 10572
rect 4291 10507 4357 10508
rect 4107 10300 4173 10301
rect 4107 10236 4108 10300
rect 4172 10236 4173 10300
rect 4107 10235 4173 10236
rect 4294 10162 4354 10507
rect 4110 10102 4354 10162
rect 3742 9966 3940 10026
rect 3739 9892 3805 9893
rect 3739 9828 3740 9892
rect 3804 9890 3805 9892
rect 3880 9890 3940 9966
rect 4110 9890 4170 10102
rect 4291 10028 4357 10029
rect 4291 10026 4292 10028
rect 3804 9830 4170 9890
rect 4248 9964 4292 10026
rect 4356 9964 4357 10028
rect 4248 9963 4357 9964
rect 3804 9828 3805 9830
rect 3739 9827 3805 9828
rect 3739 9756 3805 9757
rect 3739 9692 3740 9756
rect 3804 9692 3805 9756
rect 3739 9691 3805 9692
rect 3742 9213 3802 9691
rect 3880 9690 3940 9830
rect 3880 9630 3986 9690
rect 3739 9212 3805 9213
rect 3739 9148 3740 9212
rect 3804 9148 3805 9212
rect 3739 9147 3805 9148
rect 3739 8940 3805 8941
rect 3739 8876 3740 8940
rect 3804 8876 3805 8940
rect 3739 8875 3805 8876
rect 3555 8668 3621 8669
rect 3555 8604 3556 8668
rect 3620 8604 3621 8668
rect 3555 8603 3621 8604
rect 3558 7853 3618 8603
rect 3555 7852 3621 7853
rect 3555 7788 3556 7852
rect 3620 7788 3621 7852
rect 3555 7787 3621 7788
rect 3742 4725 3802 8875
rect 3739 4724 3805 4725
rect 3739 4660 3740 4724
rect 3804 4660 3805 4724
rect 3739 4659 3805 4660
rect 3926 3637 3986 9630
rect 4248 9618 4308 9963
rect 4248 9558 4354 9618
rect 4107 8804 4173 8805
rect 4107 8740 4108 8804
rect 4172 8740 4173 8804
rect 4107 8739 4173 8740
rect 4110 7034 4170 8739
rect 4294 7173 4354 9558
rect 4291 7172 4357 7173
rect 4291 7108 4292 7172
rect 4356 7108 4357 7172
rect 4291 7107 4357 7108
rect 4110 6974 4354 7034
rect 4294 6221 4354 6974
rect 4107 6220 4173 6221
rect 4107 6156 4108 6220
rect 4172 6156 4173 6220
rect 4107 6155 4173 6156
rect 4291 6220 4357 6221
rect 4291 6156 4292 6220
rect 4356 6156 4357 6220
rect 4291 6155 4357 6156
rect 4110 3909 4170 6155
rect 4107 3908 4173 3909
rect 4107 3844 4108 3908
rect 4172 3844 4173 3908
rect 4107 3843 4173 3844
rect 3923 3636 3989 3637
rect 3923 3572 3924 3636
rect 3988 3572 3989 3636
rect 3923 3571 3989 3572
rect 3371 2956 3437 2957
rect 3371 2892 3372 2956
rect 3436 2892 3437 2956
rect 3371 2891 3437 2892
rect 1347 2684 1413 2685
rect 1347 2620 1348 2684
rect 1412 2620 1413 2684
rect 1347 2619 1413 2620
rect 4294 2005 4354 6155
rect 4478 5813 4538 13635
rect 4659 13564 4725 13565
rect 4659 13500 4660 13564
rect 4724 13500 4725 13564
rect 4659 13499 4725 13500
rect 4662 9621 4722 13499
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 5398 11525 5458 16899
rect 5579 13020 5645 13021
rect 5579 12956 5580 13020
rect 5644 12956 5645 13020
rect 5579 12955 5645 12956
rect 5395 11524 5461 11525
rect 5395 11460 5396 11524
rect 5460 11460 5461 11524
rect 5395 11459 5461 11460
rect 5395 11388 5461 11389
rect 5395 11324 5396 11388
rect 5460 11324 5461 11388
rect 5395 11323 5461 11324
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 4659 9212 4725 9213
rect 4659 9148 4660 9212
rect 4724 9148 4725 9212
rect 4659 9147 4725 9148
rect 4662 8261 4722 9147
rect 4944 8736 5264 9760
rect 5398 9757 5458 11323
rect 5395 9756 5461 9757
rect 5395 9692 5396 9756
rect 5460 9692 5461 9756
rect 5395 9691 5461 9692
rect 5395 9212 5461 9213
rect 5395 9148 5396 9212
rect 5460 9148 5461 9212
rect 5395 9147 5461 9148
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4659 8260 4725 8261
rect 4659 8196 4660 8260
rect 4724 8196 4725 8260
rect 4659 8195 4725 8196
rect 4475 5812 4541 5813
rect 4475 5748 4476 5812
rect 4540 5748 4541 5812
rect 4475 5747 4541 5748
rect 4475 5540 4541 5541
rect 4475 5476 4476 5540
rect 4540 5538 4541 5540
rect 4662 5538 4722 8195
rect 4540 5478 4722 5538
rect 4944 7648 5264 8672
rect 5398 8394 5458 9147
rect 5582 9077 5642 12955
rect 5579 9076 5645 9077
rect 5579 9012 5580 9076
rect 5644 9012 5645 9076
rect 5579 9011 5645 9012
rect 5398 8334 5642 8394
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4540 5476 4541 5478
rect 4475 5475 4541 5476
rect 4944 5472 5264 6496
rect 5582 5541 5642 8334
rect 5766 7853 5826 17174
rect 5947 15876 6013 15877
rect 5947 15812 5948 15876
rect 6012 15812 6013 15876
rect 5947 15811 6013 15812
rect 5950 13701 6010 15811
rect 6318 15602 6378 18395
rect 6088 15542 6378 15602
rect 6502 15602 6562 18667
rect 6683 16556 6749 16557
rect 6683 16492 6684 16556
rect 6748 16492 6749 16556
rect 6683 16491 6749 16492
rect 6502 15542 6608 15602
rect 6088 15058 6148 15542
rect 6088 14998 6194 15058
rect 6134 14653 6194 14998
rect 6131 14652 6197 14653
rect 6131 14588 6132 14652
rect 6196 14588 6197 14652
rect 6131 14587 6197 14588
rect 6318 14106 6378 15182
rect 6548 15058 6608 15542
rect 6088 14046 6378 14106
rect 6502 14998 6608 15058
rect 5947 13700 6013 13701
rect 5947 13636 5948 13700
rect 6012 13636 6013 13700
rect 6088 13698 6148 14046
rect 6502 13973 6562 14998
rect 6499 13972 6565 13973
rect 6499 13908 6500 13972
rect 6564 13908 6565 13972
rect 6499 13907 6565 13908
rect 6315 13700 6381 13701
rect 6088 13638 6194 13698
rect 5947 13635 6013 13636
rect 5763 7852 5829 7853
rect 5763 7788 5764 7852
rect 5828 7788 5829 7852
rect 5763 7787 5829 7788
rect 5763 7716 5829 7717
rect 5763 7652 5764 7716
rect 5828 7652 5829 7716
rect 5763 7651 5829 7652
rect 5579 5540 5645 5541
rect 5579 5476 5580 5540
rect 5644 5476 5645 5540
rect 5579 5475 5645 5476
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 5582 3637 5642 5475
rect 5766 4861 5826 7651
rect 5950 6221 6010 13635
rect 6134 7173 6194 13638
rect 6315 13636 6316 13700
rect 6380 13636 6381 13700
rect 6686 13698 6746 16491
rect 6870 14109 6930 19347
rect 6867 14108 6933 14109
rect 6867 14044 6868 14108
rect 6932 14044 6933 14108
rect 6867 14043 6933 14044
rect 7054 13970 7114 20163
rect 7419 19820 7485 19821
rect 7419 19756 7420 19820
rect 7484 19756 7485 19820
rect 7419 19755 7485 19756
rect 7235 16964 7301 16965
rect 7235 16900 7236 16964
rect 7300 16900 7301 16964
rect 7235 16899 7301 16900
rect 7238 13973 7298 16899
rect 7422 14517 7482 19755
rect 7603 19004 7669 19005
rect 7603 18940 7604 19004
rect 7668 18940 7669 19004
rect 7603 18939 7669 18940
rect 7606 17373 7666 18939
rect 7603 17372 7669 17373
rect 7603 17308 7604 17372
rect 7668 17308 7669 17372
rect 7603 17307 7669 17308
rect 7787 16556 7853 16557
rect 7787 16492 7788 16556
rect 7852 16492 7853 16556
rect 7787 16491 7853 16492
rect 7603 16284 7669 16285
rect 7603 16220 7604 16284
rect 7668 16220 7669 16284
rect 7603 16219 7669 16220
rect 7419 14516 7485 14517
rect 7419 14452 7420 14516
rect 7484 14452 7485 14516
rect 7419 14451 7485 14452
rect 6870 13910 7114 13970
rect 7235 13972 7301 13973
rect 6870 13830 6930 13910
rect 7235 13908 7236 13972
rect 7300 13908 7301 13972
rect 7235 13907 7301 13908
rect 7419 13836 7485 13837
rect 6870 13770 7114 13830
rect 7419 13772 7420 13836
rect 7484 13772 7485 13836
rect 7419 13771 7485 13772
rect 6315 13635 6381 13636
rect 6502 13638 6746 13698
rect 6131 7172 6197 7173
rect 6131 7108 6132 7172
rect 6196 7108 6197 7172
rect 6131 7107 6197 7108
rect 6131 6628 6197 6629
rect 6131 6564 6132 6628
rect 6196 6564 6197 6628
rect 6131 6563 6197 6564
rect 5947 6220 6013 6221
rect 5947 6156 5948 6220
rect 6012 6156 6013 6220
rect 5947 6155 6013 6156
rect 5763 4860 5829 4861
rect 5763 4796 5764 4860
rect 5828 4796 5829 4860
rect 5763 4795 5829 4796
rect 6134 3773 6194 6563
rect 6318 4317 6378 13635
rect 6502 4861 6562 13638
rect 6867 12340 6933 12341
rect 6867 12276 6868 12340
rect 6932 12276 6933 12340
rect 6867 12275 6933 12276
rect 6683 10028 6749 10029
rect 6683 9964 6684 10028
rect 6748 9964 6749 10028
rect 6683 9963 6749 9964
rect 6686 7853 6746 9963
rect 6870 7986 6930 12275
rect 7054 8941 7114 13770
rect 7235 13564 7301 13565
rect 7235 13500 7236 13564
rect 7300 13500 7301 13564
rect 7235 13499 7301 13500
rect 7238 11389 7298 13499
rect 7235 11388 7301 11389
rect 7235 11324 7236 11388
rect 7300 11324 7301 11388
rect 7235 11323 7301 11324
rect 7238 10437 7298 11323
rect 7235 10436 7301 10437
rect 7235 10372 7236 10436
rect 7300 10372 7301 10436
rect 7235 10371 7301 10372
rect 7235 10300 7301 10301
rect 7235 10236 7236 10300
rect 7300 10236 7301 10300
rect 7235 10235 7301 10236
rect 7051 8940 7117 8941
rect 7051 8876 7052 8940
rect 7116 8876 7117 8940
rect 7051 8875 7117 8876
rect 6870 7926 7114 7986
rect 6683 7852 6749 7853
rect 6683 7788 6684 7852
rect 6748 7788 6749 7852
rect 6683 7787 6749 7788
rect 6867 7852 6933 7853
rect 6867 7788 6868 7852
rect 6932 7788 6933 7852
rect 6867 7787 6933 7788
rect 6683 7172 6749 7173
rect 6683 7108 6684 7172
rect 6748 7108 6749 7172
rect 6683 7107 6749 7108
rect 6499 4860 6565 4861
rect 6499 4796 6500 4860
rect 6564 4796 6565 4860
rect 6499 4795 6565 4796
rect 6315 4316 6381 4317
rect 6315 4252 6316 4316
rect 6380 4252 6381 4316
rect 6315 4251 6381 4252
rect 6686 4181 6746 7107
rect 6683 4180 6749 4181
rect 6683 4116 6684 4180
rect 6748 4116 6749 4180
rect 6683 4115 6749 4116
rect 6131 3772 6197 3773
rect 6131 3708 6132 3772
rect 6196 3708 6197 3772
rect 6131 3707 6197 3708
rect 6499 3772 6565 3773
rect 6499 3708 6500 3772
rect 6564 3708 6565 3772
rect 6499 3707 6565 3708
rect 5579 3636 5645 3637
rect 5579 3572 5580 3636
rect 5644 3572 5645 3636
rect 5579 3571 5645 3572
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 6502 3093 6562 3707
rect 6870 3093 6930 7787
rect 7054 3909 7114 7926
rect 7238 4317 7298 10235
rect 7235 4316 7301 4317
rect 7235 4252 7236 4316
rect 7300 4252 7301 4316
rect 7235 4251 7301 4252
rect 7051 3908 7117 3909
rect 7051 3844 7052 3908
rect 7116 3844 7117 3908
rect 7051 3843 7117 3844
rect 7422 3093 7482 13771
rect 7606 13565 7666 16219
rect 7790 15469 7850 16491
rect 7787 15468 7853 15469
rect 7787 15404 7788 15468
rect 7852 15404 7853 15468
rect 7787 15403 7853 15404
rect 7603 13564 7669 13565
rect 7603 13500 7604 13564
rect 7668 13500 7669 13564
rect 7603 13499 7669 13500
rect 7603 13428 7669 13429
rect 7603 13364 7604 13428
rect 7668 13364 7669 13428
rect 7603 13363 7669 13364
rect 7606 10573 7666 13363
rect 7603 10572 7669 10573
rect 7603 10508 7604 10572
rect 7668 10508 7669 10572
rect 7603 10507 7669 10508
rect 7603 9756 7669 9757
rect 7603 9692 7604 9756
rect 7668 9692 7669 9756
rect 7603 9691 7669 9692
rect 7606 6221 7666 9691
rect 7790 8941 7850 15403
rect 7974 12341 8034 22747
rect 17907 22676 17973 22677
rect 17907 22612 17908 22676
rect 17972 22612 17973 22676
rect 17907 22611 17973 22612
rect 15699 22404 15765 22405
rect 15699 22340 15700 22404
rect 15764 22340 15765 22404
rect 15699 22339 15765 22340
rect 12387 22268 12453 22269
rect 12387 22204 12388 22268
rect 12452 22204 12453 22268
rect 12387 22203 12453 22204
rect 8944 21248 9264 21808
rect 10547 21588 10613 21589
rect 10547 21524 10548 21588
rect 10612 21524 10613 21588
rect 10547 21523 10613 21524
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8707 20364 8773 20365
rect 8707 20300 8708 20364
rect 8772 20300 8773 20364
rect 8707 20299 8773 20300
rect 8155 19684 8221 19685
rect 8155 19620 8156 19684
rect 8220 19620 8221 19684
rect 8155 19619 8221 19620
rect 8158 14058 8218 19619
rect 8710 19498 8770 20299
rect 8944 20160 9264 21184
rect 9811 21044 9877 21045
rect 9811 20980 9812 21044
rect 9876 20980 9877 21044
rect 9811 20979 9877 20980
rect 9627 20942 9693 20943
rect 9627 20878 9628 20942
rect 9692 20878 9693 20942
rect 9627 20877 9693 20878
rect 9630 20770 9690 20877
rect 9814 20770 9874 20979
rect 9630 20710 9874 20770
rect 10179 20772 10245 20773
rect 10179 20708 10180 20772
rect 10244 20708 10245 20772
rect 10179 20707 10245 20708
rect 10182 20178 10242 20707
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8339 18460 8405 18461
rect 8339 18396 8340 18460
rect 8404 18396 8405 18460
rect 8339 18395 8405 18396
rect 8342 14653 8402 18395
rect 8710 18325 8770 18582
rect 8707 18324 8773 18325
rect 8707 18260 8708 18324
rect 8772 18260 8773 18324
rect 8707 18259 8773 18260
rect 8523 18052 8589 18053
rect 8523 17988 8524 18052
rect 8588 17988 8589 18052
rect 8523 17987 8589 17988
rect 8339 14652 8405 14653
rect 8339 14588 8340 14652
rect 8404 14588 8405 14652
rect 8339 14587 8405 14588
rect 7971 12340 8037 12341
rect 7971 12276 7972 12340
rect 8036 12276 8037 12340
rect 7971 12275 8037 12276
rect 7971 12068 8037 12069
rect 7971 12004 7972 12068
rect 8036 12004 8037 12068
rect 7971 12003 8037 12004
rect 7787 8940 7853 8941
rect 7787 8876 7788 8940
rect 7852 8876 7853 8940
rect 7787 8875 7853 8876
rect 7787 6764 7853 6765
rect 7787 6700 7788 6764
rect 7852 6700 7853 6764
rect 7787 6699 7853 6700
rect 7603 6220 7669 6221
rect 7603 6156 7604 6220
rect 7668 6156 7669 6220
rect 7603 6155 7669 6156
rect 7790 4042 7850 6699
rect 7974 4861 8034 12003
rect 8158 4997 8218 13822
rect 8339 13564 8405 13565
rect 8339 13500 8340 13564
rect 8404 13500 8405 13564
rect 8339 13499 8405 13500
rect 8342 12749 8402 13499
rect 8526 13293 8586 17987
rect 8944 17984 9264 19008
rect 10179 18596 10245 18597
rect 10179 18532 10180 18596
rect 10244 18532 10245 18596
rect 10179 18531 10245 18532
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8707 17780 8773 17781
rect 8707 17716 8708 17780
rect 8772 17716 8773 17780
rect 8707 17715 8773 17716
rect 8523 13292 8589 13293
rect 8523 13228 8524 13292
rect 8588 13228 8589 13292
rect 8523 13227 8589 13228
rect 8339 12748 8405 12749
rect 8339 12684 8340 12748
rect 8404 12684 8405 12748
rect 8339 12683 8405 12684
rect 8342 11930 8402 12683
rect 8526 12069 8586 13227
rect 8710 12749 8770 17715
rect 8944 16896 9264 17920
rect 9627 17644 9693 17645
rect 9627 17580 9628 17644
rect 9692 17580 9693 17644
rect 9627 17579 9693 17580
rect 9443 17372 9509 17373
rect 9443 17308 9444 17372
rect 9508 17308 9509 17372
rect 9443 17307 9509 17308
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8707 12748 8773 12749
rect 8707 12684 8708 12748
rect 8772 12684 8773 12748
rect 8707 12683 8773 12684
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8523 12068 8589 12069
rect 8523 12004 8524 12068
rect 8588 12004 8589 12068
rect 8523 12003 8589 12004
rect 8342 11870 8586 11930
rect 8339 11388 8405 11389
rect 8339 11324 8340 11388
rect 8404 11324 8405 11388
rect 8339 11323 8405 11324
rect 8342 10845 8402 11323
rect 8339 10844 8405 10845
rect 8339 10780 8340 10844
rect 8404 10780 8405 10844
rect 8339 10779 8405 10780
rect 8339 10028 8405 10029
rect 8339 9964 8340 10028
rect 8404 9964 8405 10028
rect 8339 9963 8405 9964
rect 8155 4996 8221 4997
rect 8155 4932 8156 4996
rect 8220 4932 8221 4996
rect 8155 4931 8221 4932
rect 7971 4860 8037 4861
rect 7971 4796 7972 4860
rect 8036 4796 8037 4860
rect 7971 4795 8037 4796
rect 8342 4317 8402 9963
rect 8526 4317 8586 11870
rect 8944 11456 9264 12480
rect 9446 12338 9506 17307
rect 9630 12613 9690 17579
rect 10182 13973 10242 18531
rect 10550 14245 10610 21523
rect 11651 17236 11717 17237
rect 11651 17172 11652 17236
rect 11716 17172 11717 17236
rect 11651 17171 11717 17172
rect 11467 16284 11533 16285
rect 11467 16220 11468 16284
rect 11532 16220 11533 16284
rect 11467 16219 11533 16220
rect 11099 15604 11165 15605
rect 11099 15540 11100 15604
rect 11164 15540 11165 15604
rect 11099 15539 11165 15540
rect 10731 15060 10797 15061
rect 10731 14996 10732 15060
rect 10796 14996 10797 15060
rect 10731 14995 10797 14996
rect 10547 14244 10613 14245
rect 10547 14180 10548 14244
rect 10612 14180 10613 14244
rect 10547 14179 10613 14180
rect 10179 13972 10245 13973
rect 10179 13908 10180 13972
rect 10244 13908 10245 13972
rect 10179 13907 10245 13908
rect 9995 13292 10061 13293
rect 9995 13228 9996 13292
rect 10060 13228 10061 13292
rect 9995 13227 10061 13228
rect 9998 12749 10058 13227
rect 10547 13156 10613 13157
rect 10547 13092 10548 13156
rect 10612 13092 10613 13156
rect 10547 13091 10613 13092
rect 10179 13020 10245 13021
rect 10179 12956 10180 13020
rect 10244 12956 10245 13020
rect 10179 12955 10245 12956
rect 9995 12748 10061 12749
rect 9995 12684 9996 12748
rect 10060 12684 10061 12748
rect 9995 12683 10061 12684
rect 9627 12612 9693 12613
rect 9627 12548 9628 12612
rect 9692 12548 9693 12612
rect 9627 12547 9693 12548
rect 9446 12278 9874 12338
rect 9814 11794 9874 12278
rect 10182 12069 10242 12955
rect 10363 12340 10429 12341
rect 10363 12276 10364 12340
rect 10428 12276 10429 12340
rect 10363 12275 10429 12276
rect 10179 12068 10245 12069
rect 10179 12004 10180 12068
rect 10244 12004 10245 12068
rect 10179 12003 10245 12004
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8707 9892 8773 9893
rect 8707 9828 8708 9892
rect 8772 9828 8773 9892
rect 8707 9827 8773 9828
rect 8710 9621 8770 9827
rect 8707 9620 8773 9621
rect 8707 9556 8708 9620
rect 8772 9556 8773 9620
rect 8707 9555 8773 9556
rect 8944 9280 9264 10304
rect 9446 11734 9874 11794
rect 9446 10162 9506 11734
rect 9630 10162 9690 10422
rect 9446 10102 9874 10162
rect 9443 9892 9509 9893
rect 9443 9828 9444 9892
rect 9508 9890 9509 9892
rect 9630 9890 9690 10102
rect 9508 9830 9690 9890
rect 9508 9828 9509 9830
rect 9443 9827 9509 9828
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8707 8940 8773 8941
rect 8707 8876 8708 8940
rect 8772 8876 8773 8940
rect 8707 8875 8773 8876
rect 8339 4316 8405 4317
rect 8339 4252 8340 4316
rect 8404 4252 8405 4316
rect 8339 4251 8405 4252
rect 8523 4316 8589 4317
rect 8523 4252 8524 4316
rect 8588 4252 8589 4316
rect 8523 4251 8589 4252
rect 7606 3982 7850 4042
rect 6499 3092 6565 3093
rect 6499 3028 6500 3092
rect 6564 3028 6565 3092
rect 6499 3027 6565 3028
rect 6867 3092 6933 3093
rect 6867 3028 6868 3092
rect 6932 3028 6933 3092
rect 6867 3027 6933 3028
rect 7419 3092 7485 3093
rect 7419 3028 7420 3092
rect 7484 3028 7485 3092
rect 7419 3027 7485 3028
rect 6502 2277 6562 3027
rect 7606 2685 7666 3982
rect 8710 2957 8770 8875
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 9446 4181 9506 9827
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 9443 4180 9509 4181
rect 9443 4116 9444 4180
rect 9508 4116 9509 4180
rect 9443 4115 9509 4116
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8707 2956 8773 2957
rect 8707 2892 8708 2956
rect 8772 2892 8773 2956
rect 8707 2891 8773 2892
rect 8944 2752 9264 3776
rect 9630 3093 9690 9691
rect 9814 7445 9874 10102
rect 9811 7444 9877 7445
rect 9811 7380 9812 7444
rect 9876 7380 9877 7444
rect 9811 7379 9877 7380
rect 9814 4861 9874 7379
rect 9998 5813 10058 11102
rect 10179 10980 10245 10981
rect 10179 10916 10180 10980
rect 10244 10916 10245 10980
rect 10179 10915 10245 10916
rect 9995 5812 10061 5813
rect 9995 5748 9996 5812
rect 10060 5748 10061 5812
rect 9995 5747 10061 5748
rect 9998 4997 10058 5747
rect 9995 4996 10061 4997
rect 9995 4932 9996 4996
rect 10060 4932 10061 4996
rect 9995 4931 10061 4932
rect 10182 4861 10242 10915
rect 10366 9077 10426 12275
rect 10363 9076 10429 9077
rect 10363 9012 10364 9076
rect 10428 9012 10429 9076
rect 10363 9011 10429 9012
rect 10363 8940 10429 8941
rect 10363 8876 10364 8940
rect 10428 8876 10429 8940
rect 10363 8875 10429 8876
rect 10366 8258 10426 8875
rect 10550 8397 10610 13091
rect 10734 11797 10794 14995
rect 10915 12068 10981 12069
rect 10915 12004 10916 12068
rect 10980 12004 10981 12068
rect 10915 12003 10981 12004
rect 10731 11796 10797 11797
rect 10731 11732 10732 11796
rect 10796 11732 10797 11796
rect 10731 11731 10797 11732
rect 10918 9893 10978 12003
rect 11102 10029 11162 15539
rect 11283 15468 11349 15469
rect 11283 15404 11284 15468
rect 11348 15404 11349 15468
rect 11283 15403 11349 15404
rect 11286 11117 11346 15403
rect 11470 11253 11530 16219
rect 11467 11252 11533 11253
rect 11467 11188 11468 11252
rect 11532 11188 11533 11252
rect 11467 11187 11533 11188
rect 11283 11116 11349 11117
rect 11283 11052 11284 11116
rect 11348 11052 11349 11116
rect 11283 11051 11349 11052
rect 11283 10436 11349 10437
rect 11283 10372 11284 10436
rect 11348 10372 11349 10436
rect 11283 10371 11349 10372
rect 11099 10028 11165 10029
rect 11099 9964 11100 10028
rect 11164 9964 11165 10028
rect 11099 9963 11165 9964
rect 10915 9892 10981 9893
rect 10915 9828 10916 9892
rect 10980 9828 10981 9892
rect 10915 9827 10981 9828
rect 10915 9484 10981 9485
rect 10915 9420 10916 9484
rect 10980 9420 10981 9484
rect 10915 9419 10981 9420
rect 10547 8396 10613 8397
rect 10547 8332 10548 8396
rect 10612 8332 10613 8396
rect 10547 8331 10613 8332
rect 10366 8198 10610 8258
rect 10363 8124 10429 8125
rect 10363 8060 10364 8124
rect 10428 8060 10429 8124
rect 10363 8059 10429 8060
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 10179 4860 10245 4861
rect 10179 4796 10180 4860
rect 10244 4796 10245 4860
rect 10179 4795 10245 4796
rect 10366 4045 10426 8059
rect 10363 4044 10429 4045
rect 10363 3980 10364 4044
rect 10428 3980 10429 4044
rect 10363 3979 10429 3980
rect 10550 3637 10610 8198
rect 10731 5540 10797 5541
rect 10731 5476 10732 5540
rect 10796 5476 10797 5540
rect 10731 5475 10797 5476
rect 10734 4317 10794 5475
rect 10731 4316 10797 4317
rect 10731 4252 10732 4316
rect 10796 4252 10797 4316
rect 10731 4251 10797 4252
rect 10547 3636 10613 3637
rect 10547 3572 10548 3636
rect 10612 3572 10613 3636
rect 10547 3571 10613 3572
rect 10918 3501 10978 9419
rect 11286 8938 11346 10371
rect 11654 10029 11714 17171
rect 11835 16692 11901 16693
rect 11835 16628 11836 16692
rect 11900 16628 11901 16692
rect 11835 16627 11901 16628
rect 11651 10028 11717 10029
rect 11651 9964 11652 10028
rect 11716 9964 11717 10028
rect 11651 9963 11717 9964
rect 11467 9892 11533 9893
rect 11467 9828 11468 9892
rect 11532 9828 11533 9892
rect 11467 9827 11533 9828
rect 11102 8878 11346 8938
rect 11102 5541 11162 8878
rect 11283 8804 11349 8805
rect 11283 8740 11284 8804
rect 11348 8740 11349 8804
rect 11283 8739 11349 8740
rect 11099 5540 11165 5541
rect 11099 5476 11100 5540
rect 11164 5476 11165 5540
rect 11099 5475 11165 5476
rect 11286 5218 11346 8739
rect 11470 8125 11530 9827
rect 11651 9212 11717 9213
rect 11651 9148 11652 9212
rect 11716 9148 11717 9212
rect 11651 9147 11717 9148
rect 11467 8124 11533 8125
rect 11467 8060 11468 8124
rect 11532 8060 11533 8124
rect 11467 8059 11533 8060
rect 11654 5541 11714 9147
rect 11838 8261 11898 16627
rect 12019 14924 12085 14925
rect 12019 14860 12020 14924
rect 12084 14860 12085 14924
rect 12019 14859 12085 14860
rect 11835 8260 11901 8261
rect 11835 8196 11836 8260
rect 11900 8196 11901 8260
rect 11835 8195 11901 8196
rect 11835 8124 11901 8125
rect 11835 8060 11836 8124
rect 11900 8060 11901 8124
rect 11835 8059 11901 8060
rect 11651 5540 11717 5541
rect 11651 5476 11652 5540
rect 11716 5476 11717 5540
rect 11651 5475 11717 5476
rect 11838 4997 11898 8059
rect 12022 7581 12082 14859
rect 12203 14108 12269 14109
rect 12203 14044 12204 14108
rect 12268 14044 12269 14108
rect 12203 14043 12269 14044
rect 12206 9349 12266 14043
rect 12390 13973 12450 22203
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12755 20772 12821 20773
rect 12755 20708 12756 20772
rect 12820 20708 12821 20772
rect 12755 20707 12821 20708
rect 12758 18597 12818 20707
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12755 18596 12821 18597
rect 12755 18532 12756 18596
rect 12820 18532 12821 18596
rect 12755 18531 12821 18532
rect 12758 15877 12818 18531
rect 12944 18528 13264 19552
rect 13675 19412 13741 19413
rect 13675 19348 13676 19412
rect 13740 19348 13741 19412
rect 13675 19347 13741 19348
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 13678 16557 13738 19347
rect 14043 19004 14109 19005
rect 14043 18940 14044 19004
rect 14108 18940 14109 19004
rect 14043 18939 14109 18940
rect 13675 16556 13741 16557
rect 13675 16492 13676 16556
rect 13740 16492 13741 16556
rect 13675 16491 13741 16492
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12755 15876 12821 15877
rect 12755 15812 12756 15876
rect 12820 15812 12821 15876
rect 12755 15811 12821 15812
rect 12571 15196 12637 15197
rect 12571 15132 12572 15196
rect 12636 15132 12637 15196
rect 12571 15131 12637 15132
rect 12387 13972 12453 13973
rect 12387 13908 12388 13972
rect 12452 13908 12453 13972
rect 12387 13907 12453 13908
rect 12574 12477 12634 15131
rect 12571 12476 12637 12477
rect 12571 12412 12572 12476
rect 12636 12412 12637 12476
rect 12571 12411 12637 12412
rect 12571 12068 12637 12069
rect 12571 12004 12572 12068
rect 12636 12004 12637 12068
rect 12571 12003 12637 12004
rect 12574 11661 12634 12003
rect 12758 11933 12818 15811
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 13491 14788 13557 14789
rect 13491 14724 13492 14788
rect 13556 14724 13557 14788
rect 13491 14723 13557 14724
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12755 11932 12821 11933
rect 12755 11868 12756 11932
rect 12820 11868 12821 11932
rect 12755 11867 12821 11868
rect 12571 11660 12637 11661
rect 12571 11596 12572 11660
rect 12636 11596 12637 11660
rect 12571 11595 12637 11596
rect 12387 11252 12453 11253
rect 12387 11188 12388 11252
rect 12452 11188 12453 11252
rect 12387 11187 12453 11188
rect 12203 9348 12269 9349
rect 12203 9284 12204 9348
rect 12268 9284 12269 9348
rect 12203 9283 12269 9284
rect 12203 8940 12269 8941
rect 12203 8876 12204 8940
rect 12268 8876 12269 8940
rect 12203 8875 12269 8876
rect 12019 7580 12085 7581
rect 12019 7516 12020 7580
rect 12084 7516 12085 7580
rect 12019 7515 12085 7516
rect 11835 4996 11901 4997
rect 11835 4932 11836 4996
rect 11900 4932 11901 4996
rect 11835 4931 11901 4932
rect 10915 3500 10981 3501
rect 10915 3436 10916 3500
rect 10980 3436 10981 3500
rect 10915 3435 10981 3436
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 12206 2821 12266 8875
rect 12390 5405 12450 11187
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12755 10708 12821 10709
rect 12755 10644 12756 10708
rect 12820 10644 12821 10708
rect 12755 10643 12821 10644
rect 12571 10300 12637 10301
rect 12571 10236 12572 10300
rect 12636 10236 12637 10300
rect 12571 10235 12637 10236
rect 12387 5404 12453 5405
rect 12387 5340 12388 5404
rect 12452 5340 12453 5404
rect 12387 5339 12453 5340
rect 12574 4997 12634 10235
rect 12571 4996 12637 4997
rect 12571 4932 12572 4996
rect 12636 4932 12637 4996
rect 12571 4931 12637 4932
rect 12571 4588 12637 4589
rect 12571 4524 12572 4588
rect 12636 4524 12637 4588
rect 12571 4523 12637 4524
rect 12574 2821 12634 4523
rect 12758 3637 12818 10643
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 13494 7581 13554 14723
rect 14046 13973 14106 18939
rect 14595 18732 14661 18733
rect 14595 18668 14596 18732
rect 14660 18668 14661 18732
rect 14595 18667 14661 18668
rect 14227 17916 14293 17917
rect 14227 17852 14228 17916
rect 14292 17852 14293 17916
rect 14227 17851 14293 17852
rect 14043 13972 14109 13973
rect 14043 13908 14044 13972
rect 14108 13908 14109 13972
rect 14043 13907 14109 13908
rect 13675 10844 13741 10845
rect 13675 10780 13676 10844
rect 13740 10780 13741 10844
rect 13675 10779 13741 10780
rect 13678 9978 13738 10779
rect 14230 10301 14290 17851
rect 14411 16012 14477 16013
rect 14411 15948 14412 16012
rect 14476 15948 14477 16012
rect 14411 15947 14477 15948
rect 14227 10300 14293 10301
rect 14227 10236 14228 10300
rect 14292 10236 14293 10300
rect 14227 10235 14293 10236
rect 14414 9757 14474 15947
rect 14598 12477 14658 18667
rect 15331 18052 15397 18053
rect 15331 17988 15332 18052
rect 15396 17988 15397 18052
rect 15331 17987 15397 17988
rect 14963 16964 15029 16965
rect 14963 16900 14964 16964
rect 15028 16900 15029 16964
rect 14963 16899 15029 16900
rect 14779 13564 14845 13565
rect 14779 13500 14780 13564
rect 14844 13500 14845 13564
rect 14779 13499 14845 13500
rect 14595 12476 14661 12477
rect 14595 12412 14596 12476
rect 14660 12412 14661 12476
rect 14595 12411 14661 12412
rect 14782 12018 14842 13499
rect 14966 12613 15026 16899
rect 15147 14516 15213 14517
rect 15147 14452 15148 14516
rect 15212 14452 15213 14516
rect 15147 14451 15213 14452
rect 14963 12612 15029 12613
rect 14963 12548 14964 12612
rect 15028 12548 15029 12612
rect 14963 12547 15029 12548
rect 15150 11525 15210 14451
rect 15147 11524 15213 11525
rect 15147 11460 15148 11524
rect 15212 11460 15213 11524
rect 15147 11459 15213 11460
rect 15147 10980 15213 10981
rect 15147 10916 15148 10980
rect 15212 10916 15213 10980
rect 15147 10915 15213 10916
rect 14411 9756 14477 9757
rect 14411 9692 14412 9756
rect 14476 9692 14477 9756
rect 14411 9691 14477 9692
rect 13678 9558 13922 9618
rect 13678 8941 13738 9558
rect 13675 8940 13741 8941
rect 13675 8876 13676 8940
rect 13740 8876 13741 8940
rect 13675 8875 13741 8876
rect 13862 8533 13922 9558
rect 14411 8940 14477 8941
rect 14411 8876 14412 8940
rect 14476 8876 14477 8940
rect 14411 8875 14477 8876
rect 13859 8532 13925 8533
rect 13859 8468 13860 8532
rect 13924 8468 13925 8532
rect 13859 8467 13925 8468
rect 13491 7580 13557 7581
rect 13491 7516 13492 7580
rect 13556 7516 13557 7580
rect 13491 7515 13557 7516
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 14043 5132 14109 5133
rect 14043 5068 14044 5132
rect 14108 5068 14109 5132
rect 14043 5067 14109 5068
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12755 3636 12821 3637
rect 12755 3572 12756 3636
rect 12820 3572 12821 3636
rect 12755 3571 12821 3572
rect 12944 3296 13264 4320
rect 14046 3637 14106 5067
rect 14414 3858 14474 8875
rect 15150 5133 15210 10915
rect 15334 10165 15394 17987
rect 15515 14788 15581 14789
rect 15515 14724 15516 14788
rect 15580 14724 15581 14788
rect 15515 14723 15581 14724
rect 15518 13157 15578 14723
rect 15515 13156 15581 13157
rect 15515 13092 15516 13156
rect 15580 13092 15581 13156
rect 15515 13091 15581 13092
rect 15702 11661 15762 22339
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 17355 19548 17421 19549
rect 17355 19484 17356 19548
rect 17420 19484 17421 19548
rect 17355 19483 17421 19484
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 15883 18052 15949 18053
rect 15883 17988 15884 18052
rect 15948 17988 15949 18052
rect 15883 17987 15949 17988
rect 15886 13701 15946 17987
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 17358 15877 17418 19483
rect 17539 18052 17605 18053
rect 17539 17988 17540 18052
rect 17604 17988 17605 18052
rect 17539 17987 17605 17988
rect 17355 15876 17421 15877
rect 17355 15812 17356 15876
rect 17420 15812 17421 15876
rect 17355 15811 17421 15812
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16067 15196 16133 15197
rect 16067 15132 16068 15196
rect 16132 15132 16133 15196
rect 16067 15131 16133 15132
rect 15883 13700 15949 13701
rect 15883 13636 15884 13700
rect 15948 13636 15949 13700
rect 15883 13635 15949 13636
rect 15883 13292 15949 13293
rect 15883 13228 15884 13292
rect 15948 13228 15949 13292
rect 15883 13227 15949 13228
rect 15699 11660 15765 11661
rect 15699 11596 15700 11660
rect 15764 11596 15765 11660
rect 15699 11595 15765 11596
rect 15331 10164 15397 10165
rect 15331 10100 15332 10164
rect 15396 10100 15397 10164
rect 15331 10099 15397 10100
rect 15147 5132 15213 5133
rect 15147 5068 15148 5132
rect 15212 5068 15213 5132
rect 15147 5067 15213 5068
rect 14043 3636 14109 3637
rect 14043 3572 14044 3636
rect 14108 3572 14109 3636
rect 14043 3571 14109 3572
rect 13675 3500 13741 3501
rect 13675 3436 13676 3500
rect 13740 3436 13741 3500
rect 13675 3435 13741 3436
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12203 2820 12269 2821
rect 12203 2756 12204 2820
rect 12268 2756 12269 2820
rect 12203 2755 12269 2756
rect 12571 2820 12637 2821
rect 12571 2756 12572 2820
rect 12636 2756 12637 2820
rect 12571 2755 12637 2756
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 7603 2684 7669 2685
rect 7603 2620 7604 2684
rect 7668 2620 7669 2684
rect 7603 2619 7669 2620
rect 6499 2276 6565 2277
rect 6499 2212 6500 2276
rect 6564 2212 6565 2276
rect 6499 2211 6565 2212
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 2128 9264 2688
rect 4291 2004 4357 2005
rect 4291 1940 4292 2004
rect 4356 1940 4357 2004
rect 4291 1939 4357 1940
rect 12206 1818 12266 2755
rect 12944 2208 13264 3232
rect 13678 3093 13738 3435
rect 13675 3092 13741 3093
rect 13675 3028 13676 3092
rect 13740 3028 13741 3092
rect 13675 3027 13741 3028
rect 14414 2957 14474 3622
rect 15886 3229 15946 13227
rect 16070 12477 16130 15131
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16622 14245 16682 14502
rect 16251 14244 16317 14245
rect 16251 14180 16252 14244
rect 16316 14180 16317 14244
rect 16251 14179 16317 14180
rect 16619 14244 16685 14245
rect 16619 14180 16620 14244
rect 16684 14180 16685 14244
rect 16619 14179 16685 14180
rect 16067 12476 16133 12477
rect 16067 12412 16068 12476
rect 16132 12412 16133 12476
rect 16067 12411 16133 12412
rect 16254 8941 16314 14179
rect 16619 14108 16685 14109
rect 16619 14044 16620 14108
rect 16684 14044 16685 14108
rect 16619 14043 16685 14044
rect 16251 8940 16317 8941
rect 16251 8876 16252 8940
rect 16316 8876 16317 8940
rect 16251 8875 16317 8876
rect 16622 3501 16682 14043
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16803 12748 16869 12749
rect 16803 12684 16804 12748
rect 16868 12684 16869 12748
rect 16803 12683 16869 12684
rect 16806 6085 16866 12683
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16803 6084 16869 6085
rect 16803 6020 16804 6084
rect 16868 6020 16869 6084
rect 16803 6019 16869 6020
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16619 3500 16685 3501
rect 16619 3436 16620 3500
rect 16684 3436 16685 3500
rect 16619 3435 16685 3436
rect 15883 3228 15949 3229
rect 15883 3164 15884 3228
rect 15948 3164 15949 3228
rect 15883 3163 15949 3164
rect 14411 2956 14477 2957
rect 14411 2892 14412 2956
rect 14476 2892 14477 2956
rect 14411 2891 14477 2892
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 14779 2412 14845 2413
rect 14779 2348 14780 2412
rect 14844 2348 14845 2412
rect 14779 2347 14845 2348
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 14782 1818 14842 2347
rect 16944 2128 17264 2688
rect 17358 2549 17418 15811
rect 17542 6221 17602 17987
rect 17723 15196 17789 15197
rect 17723 15132 17724 15196
rect 17788 15132 17789 15196
rect 17723 15131 17789 15132
rect 17726 10301 17786 15131
rect 17910 13429 17970 22611
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 19563 20228 19629 20229
rect 19563 20164 19564 20228
rect 19628 20164 19629 20228
rect 19563 20163 19629 20164
rect 18091 13564 18157 13565
rect 18091 13500 18092 13564
rect 18156 13500 18157 13564
rect 18091 13499 18157 13500
rect 17907 13428 17973 13429
rect 17907 13364 17908 13428
rect 17972 13364 17973 13428
rect 17907 13363 17973 13364
rect 17723 10300 17789 10301
rect 17723 10236 17724 10300
rect 17788 10236 17789 10300
rect 17723 10235 17789 10236
rect 17539 6220 17605 6221
rect 17539 6156 17540 6220
rect 17604 6156 17605 6220
rect 17539 6155 17605 6156
rect 18094 5949 18154 13499
rect 18278 9213 18338 18582
rect 18459 15468 18525 15469
rect 18459 15404 18460 15468
rect 18524 15404 18525 15468
rect 18459 15403 18525 15404
rect 18462 12341 18522 15403
rect 18459 12340 18525 12341
rect 18459 12276 18460 12340
rect 18524 12276 18525 12340
rect 18459 12275 18525 12276
rect 18830 11525 18890 17902
rect 19198 14454 19396 14514
rect 19198 14245 19258 14454
rect 19195 14244 19261 14245
rect 19195 14180 19196 14244
rect 19260 14180 19261 14244
rect 19336 14242 19396 14454
rect 19336 14182 19442 14242
rect 19195 14179 19261 14180
rect 18827 11524 18893 11525
rect 18827 11460 18828 11524
rect 18892 11460 18893 11524
rect 18827 11459 18893 11460
rect 19382 9213 19442 14182
rect 19566 10437 19626 20163
rect 20118 19350 20178 19942
rect 19750 19290 20178 19350
rect 20944 19616 21264 20640
rect 23611 20228 23677 20229
rect 23611 20164 23612 20228
rect 23676 20164 23677 20228
rect 23611 20163 23677 20164
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 19563 10436 19629 10437
rect 19563 10372 19564 10436
rect 19628 10372 19629 10436
rect 19563 10371 19629 10372
rect 18275 9212 18341 9213
rect 18275 9148 18276 9212
rect 18340 9148 18341 9212
rect 18275 9147 18341 9148
rect 19379 9212 19445 9213
rect 19379 9148 19380 9212
rect 19444 9148 19445 9212
rect 19379 9147 19445 9148
rect 19563 8940 19629 8941
rect 19563 8876 19564 8940
rect 19628 8876 19629 8940
rect 19563 8875 19629 8876
rect 18459 7580 18525 7581
rect 18459 7516 18460 7580
rect 18524 7516 18525 7580
rect 18459 7515 18525 7516
rect 18091 5948 18157 5949
rect 18091 5884 18092 5948
rect 18156 5884 18157 5948
rect 18091 5883 18157 5884
rect 18462 3909 18522 7515
rect 18827 6084 18893 6085
rect 18827 6020 18828 6084
rect 18892 6020 18893 6084
rect 18827 6019 18893 6020
rect 18459 3908 18525 3909
rect 18459 3844 18460 3908
rect 18524 3844 18525 3908
rect 18459 3843 18525 3844
rect 18830 2821 18890 6019
rect 18827 2820 18893 2821
rect 18827 2756 18828 2820
rect 18892 2756 18893 2820
rect 18827 2755 18893 2756
rect 17355 2548 17421 2549
rect 17355 2484 17356 2548
rect 17420 2484 17421 2548
rect 17355 2483 17421 2484
rect 18830 1138 18890 2755
rect 19566 1189 19626 8875
rect 19750 5133 19810 19290
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 19931 18460 19997 18461
rect 19931 18396 19932 18460
rect 19996 18396 19997 18460
rect 19931 18395 19997 18396
rect 19934 15469 19994 18395
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 19931 15468 19997 15469
rect 19931 15404 19932 15468
rect 19996 15404 19997 15468
rect 19931 15403 19997 15404
rect 19934 9077 19994 15403
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20115 13292 20181 13293
rect 20115 13228 20116 13292
rect 20180 13228 20181 13292
rect 20115 13227 20181 13228
rect 19931 9076 19997 9077
rect 19931 9012 19932 9076
rect 19996 9012 19997 9076
rect 19931 9011 19997 9012
rect 19934 6357 19994 9011
rect 19931 6356 19997 6357
rect 19931 6292 19932 6356
rect 19996 6292 19997 6356
rect 19931 6291 19997 6292
rect 19747 5132 19813 5133
rect 19747 5068 19748 5132
rect 19812 5068 19813 5132
rect 19747 5067 19813 5068
rect 20118 4861 20178 13227
rect 20302 10029 20362 15182
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20667 12340 20733 12341
rect 20667 12276 20668 12340
rect 20732 12276 20733 12340
rect 20667 12275 20733 12276
rect 20299 10028 20365 10029
rect 20299 9964 20300 10028
rect 20364 9964 20365 10028
rect 20299 9963 20365 9964
rect 20299 9756 20365 9757
rect 20299 9692 20300 9756
rect 20364 9692 20365 9756
rect 20299 9691 20365 9692
rect 20115 4860 20181 4861
rect 20115 4796 20116 4860
rect 20180 4796 20181 4860
rect 20115 4795 20181 4796
rect 19931 4724 19997 4725
rect 19931 4660 19932 4724
rect 19996 4660 19997 4724
rect 19931 4659 19997 4660
rect 19934 4538 19994 4659
rect 20302 4170 20362 9691
rect 20670 6493 20730 12275
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 21958 10301 22018 13822
rect 23614 10981 23674 20163
rect 23611 10980 23677 10981
rect 23611 10916 23612 10980
rect 23676 10916 23677 10980
rect 23611 10915 23677 10916
rect 21955 10300 22021 10301
rect 21955 10236 21956 10300
rect 22020 10236 22021 10300
rect 21955 10235 22021 10236
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20667 6492 20733 6493
rect 20667 6428 20668 6492
rect 20732 6428 20733 6492
rect 20667 6427 20733 6428
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20302 4110 20730 4170
rect 19563 1188 19629 1189
rect 19563 1124 19564 1188
rect 19628 1124 19629 1188
rect 19563 1123 19629 1124
rect 20670 101 20730 4110
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 23611 3092 23677 3093
rect 23611 3028 23612 3092
rect 23676 3028 23677 3092
rect 23611 3027 23677 3028
rect 23614 2821 23674 3027
rect 23611 2820 23677 2821
rect 23611 2756 23612 2820
rect 23676 2756 23677 2820
rect 23611 2755 23677 2756
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 23611 2004 23677 2005
rect 23611 1940 23612 2004
rect 23676 1940 23677 2004
rect 23611 1939 23677 1940
rect 23614 1733 23674 1939
rect 23611 1732 23677 1733
rect 23611 1668 23612 1732
rect 23676 1668 23677 1732
rect 23611 1667 23677 1668
rect 427 100 493 101
rect 427 36 428 100
rect 492 36 493 100
rect 427 35 493 36
rect 20667 100 20733 101
rect 20667 36 20668 100
rect 20732 36 20733 100
rect 20667 35 20733 36
<< via4 >>
rect 342 19942 578 20178
rect 710 18582 946 18818
rect 2366 19262 2602 19498
rect 4574 14502 4810 14738
rect 6230 15182 6466 15418
rect 8622 19262 8858 19498
rect 9358 20092 9594 20178
rect 9358 20028 9444 20092
rect 9444 20028 9508 20092
rect 9508 20028 9594 20092
rect 9358 19942 9594 20028
rect 10094 19942 10330 20178
rect 8622 18582 8858 18818
rect 8116 13822 8352 14058
rect 9358 12068 9594 12154
rect 9358 12004 9444 12068
rect 9444 12004 9508 12068
rect 9508 12004 9594 12068
rect 9358 11918 9594 12004
rect 9910 11102 10146 11338
rect 9588 10422 9824 10658
rect 7886 3772 8122 3858
rect 7886 3708 7972 3772
rect 7972 3708 8036 3772
rect 8036 3708 8122 3772
rect 7886 3622 8122 3708
rect 9910 4452 10146 4538
rect 9910 4388 9996 4452
rect 9996 4388 10060 4452
rect 10060 4388 10146 4452
rect 9910 4302 10146 4388
rect 11198 4982 11434 5218
rect 13636 9742 13872 9978
rect 14694 11782 14930 12018
rect 14326 3622 14562 3858
rect 16534 14502 16770 14738
rect 18190 18582 18426 18818
rect 18742 17902 18978 18138
rect 18558 11252 18794 11338
rect 18558 11188 18644 11252
rect 18644 11188 18708 11252
rect 18708 11188 18794 11252
rect 18558 11102 18794 11188
rect 18558 10572 18794 10658
rect 18558 10508 18644 10572
rect 18644 10508 18708 10572
rect 18708 10508 18794 10572
rect 18558 10422 18794 10508
rect 20030 19942 20266 20178
rect 12118 1582 12354 1818
rect 14694 1582 14930 1818
rect 20214 15182 20450 15418
rect 21870 13822 22106 14058
rect 19846 4302 20082 4538
rect 21502 9892 21738 9978
rect 21502 9828 21588 9892
rect 21588 9828 21652 9892
rect 21652 9828 21738 9892
rect 21502 9742 21738 9828
rect 20582 5132 20818 5218
rect 20582 5068 20668 5132
rect 20668 5068 20732 5132
rect 20732 5068 20818 5132
rect 20582 4982 20818 5068
rect 12302 1052 12538 1138
rect 12302 988 12388 1052
rect 12388 988 12452 1052
rect 12452 988 12538 1052
rect 12302 902 12538 988
rect 18742 902 18978 1138
<< metal5 >>
rect 300 20178 9636 20220
rect 300 19942 342 20178
rect 578 19942 9358 20178
rect 9594 19942 9636 20178
rect 300 19900 9636 19942
rect 10052 20178 20308 20220
rect 10052 19942 10094 20178
rect 10330 19942 20030 20178
rect 20266 19942 20308 20178
rect 10052 19900 20308 19942
rect 2324 19498 8900 19540
rect 2324 19262 2366 19498
rect 2602 19262 8622 19498
rect 8858 19262 8900 19498
rect 2324 19220 8900 19262
rect 668 18818 4300 18860
rect 668 18582 710 18818
rect 946 18582 4300 18818
rect 668 18540 4300 18582
rect 8580 18818 18468 18860
rect 8580 18582 8622 18818
rect 8858 18582 18190 18818
rect 18426 18582 18468 18818
rect 8580 18540 18468 18582
rect 3980 18180 4300 18540
rect 3980 18138 19020 18180
rect 3980 17902 18742 18138
rect 18978 17902 19020 18138
rect 3980 17860 19020 17902
rect 6188 15418 20492 15460
rect 6188 15182 6230 15418
rect 6466 15182 20214 15418
rect 20450 15182 20492 15418
rect 6188 15140 20492 15182
rect 4532 14738 16812 14780
rect 4532 14502 4574 14738
rect 4810 14502 16534 14738
rect 16770 14502 16812 14738
rect 4532 14460 16812 14502
rect 8074 14058 22148 14100
rect 8074 13822 8116 14058
rect 8352 13822 21870 14058
rect 22106 13822 22148 14058
rect 8074 13780 22148 13822
rect 9316 12154 9636 12196
rect 9316 11918 9358 12154
rect 9594 12060 9636 12154
rect 9594 12018 14972 12060
rect 9594 11918 14694 12018
rect 9316 11782 14694 11918
rect 14930 11782 14972 12018
rect 9316 11740 14972 11782
rect 9868 11338 18836 11380
rect 9868 11102 9910 11338
rect 10146 11102 18558 11338
rect 18794 11102 18836 11338
rect 9868 11060 18836 11102
rect 9546 10658 18836 10700
rect 9546 10422 9588 10658
rect 9824 10422 18558 10658
rect 18794 10422 18836 10658
rect 9546 10380 18836 10422
rect 13594 9978 21780 10020
rect 13594 9742 13636 9978
rect 13872 9742 21502 9978
rect 21738 9742 21780 9978
rect 13594 9700 21780 9742
rect 11156 5218 20860 5260
rect 11156 4982 11198 5218
rect 11434 4982 20582 5218
rect 20818 4982 20860 5218
rect 11156 4940 20860 4982
rect 9868 4538 20124 4580
rect 9868 4302 9910 4538
rect 10146 4302 19846 4538
rect 20082 4302 20124 4538
rect 9868 4260 20124 4302
rect 7844 3858 14604 3900
rect 7844 3622 7886 3858
rect 8122 3622 14326 3858
rect 14562 3622 14604 3858
rect 7844 3580 14604 3622
rect 12076 1818 14972 1860
rect 12076 1582 12118 1818
rect 12354 1582 14694 1818
rect 14930 1582 14972 1818
rect 12076 1540 14972 1582
rect 12260 1138 19020 1180
rect 12260 902 12302 1138
rect 12538 902 18742 1138
rect 18978 902 19020 1138
rect 12260 860 19020 902
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1050 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _179_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_29 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 1050 592
use scs8hd_nor2_4  _137_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _174_
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_92 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_164 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_173
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _183_
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_conb_1  _166_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4140 0 -1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1050 592
use scs8hd_conb_1  _170_
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_116
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _171_
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_198
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 1472 0 1 3808
box -38 -48 1050 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use scs8hd_conb_1  _160_
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  _176_
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_3_41
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_155
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_221
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_225
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_or4_4  _132_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_nand2_4  _085_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 1050 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_128
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_206
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_26
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_63
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_77
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_140
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_137
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_141
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_148
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_148
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4140 0 -1 7072
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_48
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _173_
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_194
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_198
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_9
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__D
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_78
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _162_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_96
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_100
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _161_
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_10_192
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_207
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_9
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _113_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 130 592
use scs8hd_buf_2  _178_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use scs8hd_conb_1  _163_
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_26
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__C
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_54
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _175_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _177_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_157
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_161
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_14
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use scs8hd_or4_4  _076_
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_128
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_151
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_159
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_155
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_170
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_213
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_222
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_226
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _050_
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_102
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _172_
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_226
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_230
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__D
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_60
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_101
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_170
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_207
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_232
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_43
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_210
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_176
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_180
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_6
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_20
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_24
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_28
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_147
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_176
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_193
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_10
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_146
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_37
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_134
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_203
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 222 592
use scs8hd_or3_4  _057_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_207
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _164_
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _167_
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_43
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_152
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_165
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_169
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_229
timestamp 1586364061
transform 1 0 22172 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_25
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_38
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_42
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_55
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_136
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_167
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_201
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _044_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_209
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_224 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_232
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_25
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _168_
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_42
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _169_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_82
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_37
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _165_
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_166
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_or3_4  _049_
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_201 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 21160 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_222
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_230
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_232
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_55
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_140
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_232
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 406 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_49
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _054_
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_210
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_221
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_225
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_16
timestamp 1586364061
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_20
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_25
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__D
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_75
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_87
timestamp 1586364061
transform 1 0 9108 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_101
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_134
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _048_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _083_
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_180
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_195
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_232
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_12
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_16
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_52
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_60
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_70
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_100
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_104
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_116
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use scs8hd_or4_4  _051_
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_177
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_10
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_or3_4  _059_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_or4_4  _114_
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_49
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _068_
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_66
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_73
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use scs8hd_or3_4  _055_
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__C
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_136
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__D
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_180
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_197
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_203
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_219
timestamp 1586364061
transform 1 0 21252 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_231
timestamp 1586364061
transform 1 0 22356 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 1472 0 -1 21216
box -38 -48 866 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_17
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_13
timestamp 1586364061
transform 1 0 2300 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_25
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__D
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4324 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 866 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 4508 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_63
timestamp 1586364061
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 6900 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _062_
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_72
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_76
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_67
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_85
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_or3_4  _061_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__061__C
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use scs8hd_or3_4  _053_
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 866 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_106
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__C
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _052_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_136
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_142
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_150
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_170
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_180
timestamp 1586364061
transform 1 0 17664 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_204
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_197
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_209
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_212
timestamp 1586364061
transform 1 0 20608 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_226 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_232
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__C
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_6
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_10
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _065_
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use scs8hd_or4_4  _067_
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_41
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_45
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _063_
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 6624 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_52
timestamp 1586364061
transform 1 0 5888 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_72
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_76
timestamp 1586364061
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_80
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_85
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_89
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_103
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_119
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_134
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_138
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 406 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_142
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_151
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_165
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_169
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_176
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 406 592
use scs8hd_or4_4  _086_
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_182
timestamp 1586364061
transform 1 0 17848 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__D
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_200
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_207
timestamp 1586364061
transform 1 0 20148 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_221
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_225
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 2410 0 2466 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 23520 552 24000 672 6 address[1]
port 1 nsew default input
rlabel metal2 s 938 23520 994 24000 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 280 480 400 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 960 480 1080 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[5]
port 5 nsew default input
rlabel metal2 s 2778 23520 2834 24000 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 2592 480 2712 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 23520 1640 24000 1760 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal2 s 4618 23520 4674 24000 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal2 s 3422 0 3478 480 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 6458 23520 6514 24000 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 23520 2728 24000 2848 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal2 s 6458 0 6514 480 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal2 s 7470 0 7526 480 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal2 s 8298 23520 8354 24000 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 23520 3816 24000 3936 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal2 s 10138 23520 10194 24000 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 23520 4904 24000 5024 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 12438 0 12494 480 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 23520 5992 24000 6112 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 23520 7080 24000 7200 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal2 s 13450 0 13506 480 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 11432 480 11552 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal2 s 11978 23520 12034 24000 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal2 s 14462 0 14518 480 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal2 s 13818 23520 13874 24000 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal3 s 23520 8168 24000 8288 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal3 s 23520 9256 24000 9376 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal3 s 23520 10344 24000 10464 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal3 s 23520 11432 24000 11552 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 18418 0 18474 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal2 s 15658 23520 15714 24000 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 17498 23520 17554 24000 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal3 s 23520 12520 24000 12640 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal3 s 23520 13608 24000 13728 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 19338 23520 19394 24000 6 chany_top_in[0]
port 63 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chany_top_in[1]
port 64 nsew default input
rlabel metal3 s 23520 14696 24000 14816 6 chany_top_in[2]
port 65 nsew default input
rlabel metal2 s 20442 0 20498 480 6 chany_top_in[3]
port 66 nsew default input
rlabel metal3 s 23520 15784 24000 15904 6 chany_top_in[4]
port 67 nsew default input
rlabel metal3 s 23520 16872 24000 16992 6 chany_top_in[5]
port 68 nsew default input
rlabel metal3 s 0 18504 480 18624 6 chany_top_in[6]
port 69 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chany_top_in[7]
port 70 nsew default input
rlabel metal2 s 21454 0 21510 480 6 chany_top_in[8]
port 71 nsew default input
rlabel metal3 s 23520 17960 24000 18080 6 chany_top_out[0]
port 72 nsew default tristate
rlabel metal3 s 23520 19048 24000 19168 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal3 s 23520 20136 24000 20256 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 21178 23520 21234 24000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal3 s 23520 21224 24000 21344 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 data_in
port 81 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 82 nsew default input
rlabel metal3 s 0 22584 480 22704 6 left_bottom_grid_pin_12_
port 83 nsew default input
rlabel metal3 s 23520 22312 24000 22432 6 left_top_grid_pin_10_
port 84 nsew default input
rlabel metal2 s 23018 23520 23074 24000 6 right_bottom_grid_pin_12_
port 85 nsew default input
rlabel metal2 s 23478 0 23534 480 6 right_top_grid_pin_10_
port 86 nsew default input
rlabel metal3 s 0 23400 480 23520 6 top_left_grid_pin_13_
port 87 nsew default input
rlabel metal3 s 23520 23400 24000 23520 6 top_right_grid_pin_11_
port 88 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 89 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 90 nsew default input
<< end >>
