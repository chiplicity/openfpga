* NGSPICE file created from sb_2__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sb_2__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_
+ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ prog_clk_0_N_in
+ top_left_grid_pin_42_ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_
+ top_left_grid_pin_46_ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
+ top_right_grid_pin_1_ VPWR VGND
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_062_ VGND VGND VPWR VPWR _062_/HI _062_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_061_ VGND VGND VPWR VPWR _061_/HI _061_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _083_/A sky130_fd_sc_hd__buf_4
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__buf_4
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_10.mux_l2_in_0_ _042_/HI mux_top_track_10.mux_l1_in_0_/X mux_top_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_35.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__buf_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_mem_left_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_left_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_060_ VGND VGND VPWR VPWR _060_/HI _060_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_mem_left_track_1.prog_clk clkbuf_2_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_2_0_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_7.mux_l2_in_1_ _039_/HI left_bottom_grid_pin_15_ mux_left_track_7.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_22.mux_l2_in_0_ _049_/HI mux_top_track_22.mux_l1_in_0_/X mux_top_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_10.mux_l1_in_0_ chanx_left_in[15] top_left_grid_pin_43_ mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mem_left_track_1.prog_clk clkbuf_2_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_15.mux_l2_in_0_ _058_/HI mux_left_track_15.mux_l1_in_0_/X mux_left_track_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_7.mux_l1_in_1_ left_bottom_grid_pin_11_ left_bottom_grid_pin_7_ mux_left_track_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ _041_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _096_/A sky130_fd_sc_hd__buf_4
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_2_ chanx_left_in[0] top_right_grid_pin_1_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _099_/A sky130_fd_sc_hd__buf_4
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_22.mux_l1_in_0_ chanx_left_in[9] top_left_grid_pin_49_ mux_top_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_15.mux_l1_in_0_ left_bottom_grid_pin_7_ chany_top_in[13] mux_left_track_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_27.mux_l2_in_0_ _064_/HI mux_left_track_27.mux_l1_in_0_/X mux_left_track_27.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_7.mux_l1_in_0_ left_bottom_grid_pin_3_ chany_top_in[17] mux_left_track_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_21.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_27.mux_l1_in_0_ left_bottom_grid_pin_3_ chany_top_in[7] mux_left_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_27.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_39.mux_l2_in_0_ _037_/HI mux_left_track_39.mux_l1_in_0_/X ccff_tail
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _099_/A VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_27.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_39.mux_l1_in_0_ left_bottom_grid_pin_15_ chany_top_in[1] mux_left_track_39.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_098_ _098_/A VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_27.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _085_/A sky130_fd_sc_hd__buf_4
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__buf_4
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ _097_/A VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__buf_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ _066_/HI left_bottom_grid_pin_15_ mux_left_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_096_ _096_/A VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xmux_top_track_16.mux_l2_in_0_ _045_/HI mux_top_track_16.mux_l1_in_0_/X mux_top_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_079_ _079_/A VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_20.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_ _056_/HI mux_left_track_11.mux_l1_in_0_/X mux_left_track_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_2_0_mem_left_track_1.prog_clk clkbuf_3_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_2_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l1_in_1_ left_bottom_grid_pin_11_ left_bottom_grid_pin_7_ mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_095_ _095_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _101_/A sky130_fd_sc_hd__buf_4
X_078_ _078_/A VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l1_in_0_ chanx_left_in[12] top_left_grid_pin_46_ mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5_0_mem_left_track_1.prog_clk clkbuf_3_5_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ left_bottom_grid_pin_3_ chany_top_in[15] mux_left_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_23.mux_l2_in_0_ _062_/HI mux_left_track_23.mux_l1_in_0_/X mux_left_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_26.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_26.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l1_in_0_ left_bottom_grid_pin_3_ chany_top_in[19] mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_094_ _094_/A VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_19.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_077_ _077_/A VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ _053_/HI chanx_left_in[17] mux_top_track_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_26.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_23.mux_l1_in_0_ left_bottom_grid_pin_15_ chany_top_in[9] mux_left_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_093_ chanx_left_in[6] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xmux_left_track_35.mux_l2_in_0_ _035_/HI mux_left_track_35.mux_l1_in_0_/X mux_left_track_35.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_076_ _076_/A VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_31.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ VGND VGND VPWR VPWR _059_/HI _059_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _104_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ chanx_left_in[5] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_075_ _075_/A VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_29.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_35.mux_l1_in_0_ left_bottom_grid_pin_11_ chany_top_in[3] mux_left_track_35.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ VGND VGND VPWR VPWR _058_/HI _058_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_37.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _087_/A sky130_fd_sc_hd__buf_4
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ chanx_left_in[4] VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ _074_/A VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_12.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_mem_left_track_1.prog_clk clkbuf_2_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_057_ VGND VGND VPWR VPWR _057_/HI _057_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_35.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__buf_4
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ chanx_left_in[3] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_073_ _073_/A VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_056_ VGND VGND VPWR VPWR _056_/HI _056_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_18.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_12.mux_l2_in_0_ _043_/HI mux_top_track_12.mux_l1_in_0_/X mux_top_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__buf_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_27.sky130_fd_sc_hd__buf_4_0_ mux_left_track_27.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__buf_4
X_072_ _072_/A VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ _107_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_12.mux_l1_in_0_ chanx_left_in[14] top_left_grid_pin_44_ mux_top_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_23.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_071_ _071_/A VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.mux_l2_in_0_ _059_/HI mux_left_track_17.mux_l1_in_0_/X mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_1_ _050_/HI chanx_left_in[8] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_106_ _106_/A VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_1_ _040_/HI left_bottom_grid_pin_17_ mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_2.mux_l2_in_1_ _047_/HI chanx_left_in[19] mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_070_ _070_/A VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _095_/A sky130_fd_sc_hd__buf_4
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_0_ top_right_grid_pin_1_ top_left_grid_pin_42_ mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _098_/A sky130_fd_sc_hd__buf_4
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_105_ _105_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_29.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.mux_l1_in_0_ left_bottom_grid_pin_9_ chany_top_in[12] mux_left_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_29.mux_l2_in_0_ _065_/HI mux_left_track_29.mux_l1_in_0_/X mux_left_track_29.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_31.mux_l2_in_0_ _067_/HI mux_left_track_31.mux_l1_in_0_/X mux_left_track_31.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l1_in_0_ left_bottom_grid_pin_1_ chany_top_in[16] mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XFILLER_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_27.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_104_ _104_/A VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_29.mux_l1_in_0_ left_bottom_grid_pin_5_ chany_top_in[6] mux_left_track_29.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_31.mux_l1_in_0_ left_bottom_grid_pin_7_ chany_top_in[5] mux_left_track_31.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
X_103_ _103_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_3_1_0_mem_left_track_1.prog_clk clkbuf_2_0_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_102_ _102_/A VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_22.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_15.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_4_0_mem_left_track_1.prog_clk clkbuf_3_5_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_4_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _084_/A sky130_fd_sc_hd__buf_4
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_101_ _101_/A VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__buf_4
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_mem_left_track_1.prog_clk clkbuf_3_7_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__buf_4
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_13.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_5.mux_l2_in_1_ _038_/HI mux_left_track_5.mux_l1_in_2_/X mux_left_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_100_ _100_/A VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_17_ left_bottom_grid_pin_13_ mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_18.mux_l2_in_0_ _046_/HI mux_top_track_18.mux_l1_in_0_/X mux_top_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_20.mux_l2_in_0_ _048_/HI mux_top_track_20.mux_l1_in_0_/X mux_top_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_13.mux_l2_in_0_ _057_/HI mux_left_track_13.mux_l1_in_0_/X mux_left_track_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _068_/A sky130_fd_sc_hd__buf_4
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_1_ left_bottom_grid_pin_9_ left_bottom_grid_pin_5_ mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_33.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _097_/A sky130_fd_sc_hd__buf_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _100_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_18.mux_l1_in_0_ chanx_left_in[11] top_left_grid_pin_47_ mux_top_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_20.mux_l1_in_0_ chanx_left_in[10] top_left_grid_pin_48_ mux_top_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_13.mux_l1_in_0_ left_bottom_grid_pin_5_ chany_top_in[14] mux_left_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_0_ left_bottom_grid_pin_1_ chany_top_in[18] mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l1_in_1_ _063_/HI left_bottom_grid_pin_17_ mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_089_ chanx_left_in[2] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_31.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_mem_left_track_1.prog_clk clkbuf_2_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_39.mux_l1_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_0_ left_bottom_grid_pin_1_ chany_top_in[8] mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ chanx_left_in[1] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_37.mux_l2_in_0_ _036_/HI mux_left_track_37.mux_l1_in_0_/X mux_left_track_37.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_37.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _103_/A sky130_fd_sc_hd__buf_4
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l1_in_1_ _054_/HI chanx_left_in[16] mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_087_ _087_/A VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_37.mux_l1_in_0_ left_bottom_grid_pin_13_ chany_top_in[2] mux_left_track_37.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ top_right_grid_pin_1_ top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ _086_/A VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _086_/A sky130_fd_sc_hd__buf_4
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_069_ _069_/A VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_4
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_085_ _085_/A VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_068_ _068_/A VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_1_ _055_/HI mux_left_track_1.mux_l1_in_2_/X mux_left_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_17_ left_bottom_grid_pin_13_ mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_14.mux_l2_in_0_ _044_/HI mux_top_track_14.mux_l1_in_0_/X mux_top_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _070_/A sky130_fd_sc_hd__buf_4
XFILLER_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_067_ VGND VGND VPWR VPWR _067_/HI _067_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_1_ left_bottom_grid_pin_9_ left_bottom_grid_pin_5_ mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _102_/A sky130_fd_sc_hd__buf_4
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_083_ _083_/A VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_14.mux_l1_in_0_ chanx_left_in[13] top_left_grid_pin_45_ mux_top_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_26.mux_l2_in_0_ _051_/HI mux_top_track_26.mux_l1_in_0_/X mux_top_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_066_ VGND VGND VPWR VPWR _066_/HI _066_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.mux_l2_in_0_ _060_/HI mux_left_track_19.mux_l1_in_0_/X mux_left_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_21.mux_l2_in_0_ _061_/HI mux_left_track_21.mux_l1_in_0_/X mux_left_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l1_in_0_ left_bottom_grid_pin_1_ chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_082_ _082_/A VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ _052_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_065_ VGND VGND VPWR VPWR _065_/HI _065_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_26.sky130_fd_sc_hd__buf_4_0_ mux_top_track_26.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _094_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_4.mux_l1_in_2_ chanx_left_in[18] top_right_grid_pin_1_ mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_26.mux_l1_in_0_ chanx_left_in[7] top_left_grid_pin_43_ mux_top_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_11.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_2 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_19.mux_l1_in_0_ left_bottom_grid_pin_11_ chany_top_in[11] mux_left_track_19.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_mem_left_track_1.prog_clk clkbuf_2_0_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_0_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_21.mux_l1_in_0_ left_bottom_grid_pin_13_ chany_top_in[10] mux_left_track_21.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_0_ _034_/HI mux_left_track_33.mux_l1_in_0_/X mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_081_ _081_/A VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _105_/A sky130_fd_sc_hd__buf_4
X_064_ VGND VGND VPWR VPWR _064_/HI _064_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_mem_left_track_1.prog_clk clkbuf_3_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_3 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ _080_/A VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xclkbuf_3_6_0_mem_left_track_1.prog_clk clkbuf_3_7_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_6_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l1_in_0_ left_bottom_grid_pin_9_ chany_top_in[4] mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_063_ VGND VGND VPWR VPWR _063_/HI _063_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

