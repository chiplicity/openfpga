magic
tech sky130A
magscale 1 2
timestamp 1604670029
<< viali >>
rect 22661 18921 22695 18955
rect 21373 18785 21407 18819
rect 22477 18785 22511 18819
rect 21557 18649 21591 18683
rect 21465 18037 21499 18071
rect 22569 18037 22603 18071
rect 11713 10761 11747 10795
rect 11253 10693 11287 10727
rect 11069 10557 11103 10591
rect 2789 9129 2823 9163
rect 1409 8993 1443 9027
rect 1665 8993 1699 9027
rect 1593 8585 1627 8619
rect 1961 8313 1995 8347
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 10552 2465 10586 2499
rect 10977 2465 11011 2499
rect 8769 2329 8803 2363
rect 10655 2261 10689 2295
<< metal1 >>
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 22646 18952 22652 18964
rect 22607 18924 22652 18952
rect 22646 18912 22652 18924
rect 22704 18912 22710 18964
rect 21361 18819 21419 18825
rect 21361 18785 21373 18819
rect 21407 18816 21419 18819
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 21407 18788 22477 18816
rect 21407 18785 21419 18788
rect 21361 18779 21419 18785
rect 22465 18785 22477 18788
rect 22511 18816 22523 18819
rect 22554 18816 22560 18828
rect 22511 18788 22560 18816
rect 22511 18785 22523 18788
rect 22465 18779 22523 18785
rect 22554 18776 22560 18788
rect 22612 18776 22618 18828
rect 21542 18680 21548 18692
rect 21503 18652 21548 18680
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 21453 18071 21511 18077
rect 21453 18037 21465 18071
rect 21499 18068 21511 18071
rect 22554 18068 22560 18080
rect 21499 18040 22560 18068
rect 21499 18037 21511 18040
rect 21453 18031 21511 18037
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 11698 10792 11704 10804
rect 11659 10764 11704 10792
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 11238 10724 11244 10736
rect 11199 10696 11244 10724
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11698 10588 11704 10600
rect 11103 10560 11704 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 2774 9160 2780 9172
rect 2735 9132 2780 9160
rect 2774 9120 2780 9132
rect 2832 9120 2838 9172
rect 1946 9092 1952 9104
rect 1412 9064 1952 9092
rect 1412 9033 1440 9064
rect 1946 9052 1952 9064
rect 2004 9052 2010 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1486 8984 1492 9036
rect 1544 9024 1550 9036
rect 1653 9027 1711 9033
rect 1653 9024 1665 9027
rect 1544 8996 1665 9024
rect 1544 8984 1550 8996
rect 1653 8993 1665 8996
rect 1699 8993 1711 9027
rect 1653 8987 1711 8993
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 1946 8344 1952 8356
rect 1907 8316 1952 8344
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8628 2468 9137 2496
rect 8628 2456 8634 2468
rect 9125 2465 9137 2468
rect 9171 2496 9183 2499
rect 10540 2499 10598 2505
rect 10540 2496 10552 2499
rect 9171 2468 10552 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 10540 2465 10552 2468
rect 10586 2496 10598 2499
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10586 2468 10977 2496
rect 10586 2465 10598 2468
rect 10540 2459 10598 2465
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 8757 2363 8815 2369
rect 8757 2329 8769 2363
rect 8803 2360 8815 2363
rect 11146 2360 11152 2372
rect 8803 2332 11152 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 10643 2295 10701 2301
rect 10643 2261 10655 2295
rect 10689 2292 10701 2295
rect 10870 2292 10876 2304
rect 10689 2264 10876 2292
rect 10689 2261 10701 2264
rect 10643 2255 10701 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
rect 24854 1980 24860 2032
rect 24912 2020 24918 2032
rect 26142 2020 26148 2032
rect 24912 1992 26148 2020
rect 24912 1980 24918 1992
rect 26142 1980 26148 1992
rect 26200 1980 26206 2032
<< via1 >>
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 22652 18955 22704 18964
rect 22652 18921 22661 18955
rect 22661 18921 22695 18955
rect 22695 18921 22704 18955
rect 22652 18912 22704 18921
rect 22560 18776 22612 18828
rect 21548 18683 21600 18692
rect 21548 18649 21557 18683
rect 21557 18649 21591 18683
rect 21591 18649 21600 18683
rect 21548 18640 21600 18649
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 22560 18071 22612 18080
rect 22560 18037 22569 18071
rect 22569 18037 22603 18071
rect 22603 18037 22612 18071
rect 22560 18028 22612 18037
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 11244 10727 11296 10736
rect 11244 10693 11253 10727
rect 11253 10693 11287 10727
rect 11287 10693 11296 10727
rect 11244 10684 11296 10693
rect 11704 10548 11756 10600
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 1952 9052 2004 9104
rect 1492 8984 1544 9036
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1492 8576 1544 8628
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 11152 2320 11204 2372
rect 10876 2252 10928 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
rect 24860 1980 24912 2032
rect 26148 1980 26200 2032
<< metal2 >>
rect 4986 23520 5042 24000
rect 14922 23520 14978 24000
rect 24950 23520 25006 24000
rect 2778 19952 2834 19961
rect 2778 19887 2834 19896
rect 1490 11928 1546 11937
rect 1490 11863 1546 11872
rect 1504 9042 1532 11863
rect 2792 9178 2820 19887
rect 5000 18737 5028 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 14936 19281 14964 23520
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 24964 19417 24992 23520
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 22650 19408 22706 19417
rect 22650 19343 22706 19352
rect 24950 19408 25006 19417
rect 24950 19343 25006 19352
rect 11702 19272 11758 19281
rect 11702 19207 11758 19216
rect 14922 19272 14978 19281
rect 14922 19207 14978 19216
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 4986 18728 5042 18737
rect 4986 18663 5042 18672
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 11716 10810 11744 19207
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 22664 18970 22692 19343
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 21546 18728 21602 18737
rect 21546 18663 21548 18672
rect 21600 18663 21602 18672
rect 21548 18634 21600 18640
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 22572 18086 22600 18770
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 22560 18080 22612 18086
rect 22558 18048 22560 18057
rect 22612 18048 22614 18057
rect 20956 17980 21252 18000
rect 22558 17983 22614 17992
rect 24858 18048 24914 18057
rect 24858 17983 24914 17992
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 10577 11284 10678
rect 11716 10606 11744 10746
rect 11704 10600 11756 10606
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 11242 10568 11298 10577
rect 11704 10542 11756 10548
rect 11242 10503 11298 10512
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1504 8634 1532 8978
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1964 8362 1992 9046
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1964 4049 1992 8298
rect 1950 4040 2006 4049
rect 1950 3975 2006 3984
rect 2792 2553 2820 9114
rect 2778 2544 2834 2553
rect 2778 2479 2834 2488
rect 4080 626 4108 10503
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 8574 2544 8630 2553
rect 8574 2479 8576 2488
rect 8628 2479 8630 2488
rect 8576 2450 8628 2456
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 10888 1465 10916 2246
rect 10874 1456 10930 1465
rect 10874 1391 10930 1400
rect 3712 598 4108 626
rect 3712 480 3740 598
rect 11164 480 11192 2314
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 24872 2038 24900 17983
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 26148 2032 26200 2038
rect 26148 1974 26200 1980
rect 18694 1456 18750 1465
rect 18694 1391 18750 1400
rect 18708 480 18736 1391
rect 26160 480 26188 1974
rect 3698 0 3754 480
rect 11150 0 11206 480
rect 18694 0 18750 480
rect 26146 0 26202 480
<< via2 >>
rect 2778 19896 2834 19952
rect 1490 11872 1546 11928
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 22650 19352 22706 19408
rect 24950 19352 25006 19408
rect 11702 19216 11758 19272
rect 14922 19216 14978 19272
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 4986 18672 5042 18728
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 21546 18692 21602 18728
rect 21546 18672 21548 18692
rect 21548 18672 21600 18692
rect 21600 18672 21602 18692
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 22558 18028 22560 18048
rect 22560 18028 22612 18048
rect 22612 18028 22614 18048
rect 22558 17992 22614 18028
rect 24858 17992 24914 18048
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 4066 10512 4122 10568
rect 11242 10512 11298 10568
rect 1950 3984 2006 4040
rect 2778 2488 2834 2544
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 8574 2508 8630 2544
rect 8574 2488 8576 2508
rect 8576 2488 8628 2508
rect 8628 2488 8630 2508
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 10874 1400 10930 1456
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 18694 1400 18750 1456
<< metal3 >>
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 10944 20160 11264 20161
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 0 19954 480 19984
rect 2773 19954 2839 19957
rect 0 19952 2839 19954
rect 0 19896 2778 19952
rect 2834 19896 2839 19952
rect 0 19894 2839 19896
rect 0 19864 480 19894
rect 2773 19891 2839 19894
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 22645 19410 22711 19413
rect 24945 19410 25011 19413
rect 22645 19408 25011 19410
rect 22645 19352 22650 19408
rect 22706 19352 24950 19408
rect 25006 19352 25011 19408
rect 22645 19350 25011 19352
rect 22645 19347 22711 19350
rect 24945 19347 25011 19350
rect 11697 19274 11763 19277
rect 14917 19274 14983 19277
rect 11697 19272 14983 19274
rect 11697 19216 11702 19272
rect 11758 19216 14922 19272
rect 14978 19216 14983 19272
rect 11697 19214 14983 19216
rect 11697 19211 11763 19214
rect 14917 19211 14983 19214
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 4981 18730 5047 18733
rect 21541 18730 21607 18733
rect 4981 18728 21607 18730
rect 4981 18672 4986 18728
rect 5042 18672 21546 18728
rect 21602 18672 21607 18728
rect 4981 18670 21607 18672
rect 4981 18667 5047 18670
rect 21541 18667 21607 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 22553 18050 22619 18053
rect 24853 18050 24919 18053
rect 22553 18048 24919 18050
rect 22553 17992 22558 18048
rect 22614 17992 24858 18048
rect 24914 17992 24919 18048
rect 22553 17990 24919 17992
rect 22553 17987 22619 17990
rect 24853 17987 24919 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 15743 21264 15744
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 15199 26264 15200
rect 10944 14720 11264 14721
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 5944 14176 6264 14177
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 5944 12000 6264 12001
rect 0 11930 480 11960
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 1485 11930 1551 11933
rect 0 11928 1551 11930
rect 0 11872 1490 11928
rect 1546 11872 1551 11928
rect 0 11870 1551 11872
rect 0 11840 480 11870
rect 1485 11867 1551 11870
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 4061 10570 4127 10573
rect 11237 10570 11303 10573
rect 4061 10568 11303 10570
rect 4061 10512 4066 10568
rect 4122 10512 11242 10568
rect 11298 10512 11303 10568
rect 4061 10510 11303 10512
rect 4061 10507 4127 10510
rect 11237 10507 11303 10510
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 10303 21264 10304
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 9759 26264 9760
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 9215 21264 9216
rect 5944 8736 6264 8737
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 10944 8192 11264 8193
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 4319 26264 4320
rect 0 4042 480 4072
rect 1945 4042 2011 4045
rect 0 4040 2011 4042
rect 0 3984 1950 4040
rect 2006 3984 2011 4040
rect 0 3982 2011 3984
rect 0 3952 480 3982
rect 1945 3979 2011 3982
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 3775 21264 3776
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 3231 26264 3232
rect 10944 2752 11264 2753
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 2773 2546 2839 2549
rect 8569 2546 8635 2549
rect 2773 2544 8635 2546
rect 2773 2488 2778 2544
rect 2834 2488 8574 2544
rect 8630 2488 8635 2544
rect 2773 2486 8635 2488
rect 2773 2483 2839 2486
rect 8569 2483 8635 2486
rect 5944 2208 6264 2209
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 10869 1458 10935 1461
rect 18689 1458 18755 1461
rect 10869 1456 18755 1458
rect 10869 1400 10874 1456
rect 10930 1400 18694 1456
rect 18750 1400 18755 1456
rect 10869 1398 18755 1400
rect 10869 1395 10935 1398
rect 18689 1395 18755 1398
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604666999
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604666999
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75
timestamp 1604666999
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604666999
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604666999
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1604666999
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604666999
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.ie_oe_inv tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 10488 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.ie_oe_inv_A
timestamp 1604666999
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1604666999
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_109
timestamp 1604666999
transform 1 0 11132 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1604666999
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604666999
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604666999
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604666999
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604666999
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604666999
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604666999
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604666999
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604666999
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604666999
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604666999
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604666999
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604666999
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604666999
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1604666999
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_292
timestamp 1604666999
transform 1 0 27968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1604666999
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1604666999
transform 1 0 28060 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 28520 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604666999
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604666999
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604666999
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604666999
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604666999
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604666999
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604666999
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604666999
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_288
timestamp 1604666999
transform 1 0 27600 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp 1604666999
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604666999
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604666999
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604666999
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604666999
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604666999
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604666999
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1604666999
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1604666999
transform 1 0 28060 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604666999
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604666999
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604666999
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604666999
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604666999
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604666999
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604666999
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_288
timestamp 1604666999
transform 1 0 27600 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_296
timestamp 1604666999
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604666999
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604666999
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604666999
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604666999
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604666999
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604666999
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604666999
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604666999
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604666999
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1604666999
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1604666999
transform 1 0 28060 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604666999
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604666999
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604666999
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604666999
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604666999
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604666999
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604666999
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604666999
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604666999
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604666999
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604666999
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604666999
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604666999
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604666999
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604666999
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604666999
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604666999
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604666999
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1604666999
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_288
timestamp 1604666999
transform 1 0 27600 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_296
timestamp 1604666999
transform 1 0 28336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1604666999
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1604666999
transform 1 0 28060 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604666999
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604666999
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604666999
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604666999
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604666999
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604666999
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604666999
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604666999
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604666999
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604666999
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604666999
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_288
timestamp 1604666999
transform 1 0 27600 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_296
timestamp 1604666999
transform 1 0 28336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604666999
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604666999
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604666999
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604666999
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604666999
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604666999
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604666999
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604666999
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604666999
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604666999
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604666999
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604666999
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1604666999
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1604666999
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1604666999
transform 1 0 28060 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604666999
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604666999
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604666999
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604666999
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604666999
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604666999
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604666999
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604666999
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604666999
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604666999
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_288
timestamp 1604666999
transform 1 0 27600 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_296
timestamp 1604666999
transform 1 0 28336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604666999
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_11
timestamp 1604666999
transform 1 0 2116 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_23
timestamp 1604666999
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_35
timestamp 1604666999
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_47
timestamp 1604666999
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604666999
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604666999
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604666999
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604666999
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604666999
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604666999
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604666999
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604666999
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604666999
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604666999
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1604666999
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1604666999
transform 1 0 28060 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1604666999
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604666999
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604666999
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604666999
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604666999
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604666999
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604666999
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604666999
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604666999
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604666999
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604666999
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604666999
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604666999
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604666999
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604666999
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604666999
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604666999
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_288
timestamp 1604666999
transform 1 0 27600 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1604666999
transform 1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604666999
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604666999
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604666999
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604666999
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604666999
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604666999
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604666999
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604666999
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604666999
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604666999
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604666999
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604666999
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604666999
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1604666999
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604666999
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604666999
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604666999
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604666999
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604666999
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604666999
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604666999
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604666999
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604666999
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604666999
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604666999
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604666999
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604666999
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604666999
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1604666999
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604666999
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1604666999
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1604666999
transform 1 0 28060 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_288
timestamp 1604666999
transform 1 0 27600 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_296
timestamp 1604666999
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604666999
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604666999
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604666999
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604666999
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604666999
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604666999
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0_
timestamp 1604666999
transform 1 0 11040 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0__A
timestamp 1604666999
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1604666999
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1604666999
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_116
timestamp 1604666999
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1604666999
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1604666999
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1604666999
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1604666999
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604666999
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604666999
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604666999
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604666999
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604666999
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1604666999
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1604666999
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1604666999
transform 1 0 28060 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604666999
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604666999
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604666999
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604666999
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604666999
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604666999
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604666999
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604666999
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1604666999
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604666999
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1604666999
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1604666999
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1604666999
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604666999
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604666999
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604666999
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604666999
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_288
timestamp 1604666999
transform 1 0 27600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_296
timestamp 1604666999
transform 1 0 28336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604666999
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604666999
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604666999
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604666999
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604666999
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604666999
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604666999
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604666999
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1604666999
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1604666999
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1604666999
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604666999
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604666999
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1604666999
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1604666999
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604666999
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_269
timestamp 1604666999
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1604666999
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1604666999
transform 1 0 28060 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604666999
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604666999
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604666999
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604666999
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604666999
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604666999
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604666999
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604666999
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604666999
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604666999
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604666999
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604666999
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604666999
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604666999
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604666999
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604666999
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_288
timestamp 1604666999
transform 1 0 27600 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1604666999
transform 1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604666999
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604666999
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604666999
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604666999
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604666999
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604666999
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604666999
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604666999
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604666999
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604666999
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604666999
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604666999
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604666999
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604666999
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604666999
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604666999
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604666999
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1604666999
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1604666999
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604666999
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604666999
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604666999
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604666999
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604666999
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604666999
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604666999
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604666999
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604666999
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604666999
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604666999
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604666999
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1604666999
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604666999
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1604666999
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1604666999
transform 1 0 28060 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604666999
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604666999
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604666999
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604666999
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604666999
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604666999
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604666999
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604666999
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604666999
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604666999
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604666999
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604666999
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604666999
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604666999
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604666999
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604666999
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604666999
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1604666999
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1604666999
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1604666999
transform 1 0 28060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604666999
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604666999
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604666999
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604666999
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604666999
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604666999
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604666999
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604666999
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604666999
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604666999
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604666999
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604666999
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604666999
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604666999
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604666999
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604666999
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604666999
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604666999
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604666999
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604666999
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604666999
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604666999
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604666999
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604666999
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604666999
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604666999
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604666999
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604666999
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604666999
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604666999
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604666999
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604666999
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604666999
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1604666999
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1604666999
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1604666999
transform 1 0 28060 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604666999
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604666999
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604666999
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604666999
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604666999
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604666999
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604666999
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604666999
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604666999
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604666999
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604666999
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604666999
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604666999
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604666999
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604666999
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604666999
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604666999
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp 1604666999
transform 1 0 27600 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1604666999
transform 1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604666999
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604666999
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604666999
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604666999
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604666999
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604666999
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604666999
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604666999
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604666999
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604666999
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604666999
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604666999
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604666999
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604666999
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1604666999
transform 1 0 25852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1604666999
transform 1 0 26956 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1604666999
transform 1 0 28060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604666999
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604666999
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604666999
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604666999
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604666999
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604666999
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604666999
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604666999
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604666999
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604666999
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604666999
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604666999
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604666999
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604666999
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604666999
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604666999
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604666999
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604666999
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604666999
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604666999
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604666999
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604666999
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604666999
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604666999
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604666999
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604666999
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604666999
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604666999
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604666999
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1604666999
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604666999
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1604666999
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1604666999
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1604666999
transform 1 0 28060 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604666999
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604666999
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604666999
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604666999
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604666999
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604666999
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604666999
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604666999
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604666999
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604666999
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604666999
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604666999
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604666999
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604666999
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604666999
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604666999
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604666999
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604666999
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604666999
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604666999
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604666999
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604666999
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604666999
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604666999
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604666999
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604666999
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__3__A
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2__A
timestamp 1604666999
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_222
timestamp 1604666999
transform 1 0 21528 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_230
timestamp 1604666999
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_234
timestamp 1604666999
transform 1 0 22632 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_242
timestamp 1604666999
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604666999
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1604666999
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1604666999
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1604666999
transform 1 0 28060 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604666999
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604666999
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604666999
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604666999
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604666999
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604666999
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604666999
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604666999
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604666999
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604666999
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2_
timestamp 1604666999
transform 1 0 22448 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _3_
timestamp 1604666999
transform 1 0 21344 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1604666999
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_224
timestamp 1604666999
transform 1 0 21712 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_236
timestamp 1604666999
transform 1 0 22816 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_248
timestamp 1604666999
transform 1 0 23920 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_260
timestamp 1604666999
transform 1 0 25024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1604666999
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604666999
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604666999
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604666999
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604666999
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604666999
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604666999
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604666999
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604666999
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604666999
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604666999
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604666999
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604666999
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604666999
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604666999
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1604666999
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1604666999
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1604666999
transform 1 0 28060 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604666999
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604666999
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604666999
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604666999
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604666999
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604666999
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604666999
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604666999
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604666999
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604666999
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604666999
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604666999
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604666999
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604666999
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604666999
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1604666999
transform 1 0 27600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604666999
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604666999
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604666999
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604666999
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604666999
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604666999
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604666999
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604666999
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604666999
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604666999
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604666999
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604666999
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604666999
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604666999
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604666999
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604666999
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604666999
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604666999
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604666999
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604666999
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604666999
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604666999
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604666999
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604666999
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1604666999
transform 1 0 25852 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604666999
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1604666999
transform 1 0 26956 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1604666999
transform 1 0 28060 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604666999
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604666999
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604666999
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604666999
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604666999
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604666999
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604666999
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604666999
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604666999
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604666999
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604666999
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604666999
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604666999
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604666999
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604666999
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604666999
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604666999
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604666999
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604666999
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604666999
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604666999
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604666999
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604666999
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604666999
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604666999
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604666999
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604666999
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 11840 480 11960 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 19864 480 19984 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 gfpga_pad_GPIO_A
port 2 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 gfpga_pad_GPIO_IE
port 3 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 gfpga_pad_GPIO_OE
port 4 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 gfpga_pad_GPIO_Y
port 5 nsew default bidirectional
rlabel metal3 s 0 3952 480 4072 6 prog_clk
port 6 nsew default input
rlabel metal2 s 14922 23520 14978 24000 6 top_width_0_height_0__pin_0_
port 7 nsew default input
rlabel metal2 s 24950 23520 25006 24000 6 top_width_0_height_0__pin_1_lower
port 8 nsew default tristate
rlabel metal2 s 4986 23520 5042 24000 6 top_width_0_height_0__pin_1_upper
port 9 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 10 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 11 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28926 24000
<< end >>
