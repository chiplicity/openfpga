* NGSPICE file created from grid_io_left.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_1 abstract view
.subckt scs8hd_ebufn_1 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and4_4 abstract view
.subckt scs8hd_and4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt grid_io_left address[0] address[1] address[2] address[3] data_in enable gfpga_pad_GPIO_PAD[0]
+ gfpga_pad_GPIO_PAD[1] gfpga_pad_GPIO_PAD[2] gfpga_pad_GPIO_PAD[3] gfpga_pad_GPIO_PAD[4]
+ gfpga_pad_GPIO_PAD[5] gfpga_pad_GPIO_PAD[6] gfpga_pad_GPIO_PAD[7] right_width_0_height_0__pin_0_
+ right_width_0_height_0__pin_10_ right_width_0_height_0__pin_11_ right_width_0_height_0__pin_12_
+ right_width_0_height_0__pin_13_ right_width_0_height_0__pin_14_ right_width_0_height_0__pin_15_
+ right_width_0_height_0__pin_1_ right_width_0_height_0__pin_2_ right_width_0_height_0__pin_3_
+ right_width_0_height_0__pin_4_ right_width_0_height_0__pin_5_ right_width_0_height_0__pin_6_
+ right_width_0_height_0__pin_7_ right_width_0_height_0__pin_8_ right_width_0_height_0__pin_9_
+ vpwr vgnd
XFILLER_77_15 vgnd vpwr scs8hd_decap_12
XFILLER_77_59 vpwr vgnd scs8hd_fill_2
XFILLER_172_3 vgnd vpwr scs8hd_decap_12
XFILLER_133_98 vgnd vpwr scs8hd_decap_12
XFILLER_158_105 vgnd vpwr scs8hd_decap_12
XFILLER_190_93 vgnd vpwr scs8hd_decap_12
XFILLER_179_39 vgnd vpwr scs8hd_decap_12
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_128_32 vgnd vpwr scs8hd_decap_12
XFILLER_92_117 vgnd vpwr scs8hd_decap_8
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_78_80 vgnd vpwr scs8hd_decap_12
XFILLER_114_56 vgnd vpwr scs8hd_decap_12
XFILLER_74_27 vgnd vpwr scs8hd_decap_4
XFILLER_74_117 vgnd vpwr scs8hd_decap_8
XPHY_768 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_757 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_746 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_735 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_724 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_713 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_702 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_44 vgnd vpwr scs8hd_decap_12
XFILLER_90_15 vgnd vpwr scs8hd_decap_12
XFILLER_139_86 vgnd vpwr scs8hd_decap_12
XFILLER_135_3 vgnd vpwr scs8hd_decap_12
XFILLER_155_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_121 vgnd vpwr scs8hd_decap_4
XFILLER_171_62 vgnd vpwr scs8hd_decap_12
XFILLER_171_51 vgnd vpwr scs8hd_decap_8
XFILLER_64_93 vgnd vpwr scs8hd_decap_12
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_117 vgnd vpwr scs8hd_decap_8
XFILLER_69_27 vgnd vpwr scs8hd_decap_12
XFILLER_85_15 vgnd vpwr scs8hd_decap_12
XFILLER_85_59 vpwr vgnd scs8hd_fill_2
XFILLER_141_98 vgnd vpwr scs8hd_decap_12
XPHY_598 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_587 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_576 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_565 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_38_117 vgnd vpwr scs8hd_decap_8
XFILLER_98_3 vgnd vpwr scs8hd_decap_12
XFILLER_187_39 vgnd vpwr scs8hd_decap_12
XFILLER_71_39 vgnd vpwr scs8hd_decap_12
XFILLER_136_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_4
XFILLER_45_51 vgnd vpwr scs8hd_decap_8
XFILLER_45_62 vgnd vpwr scs8hd_decap_12
XPHY_373 vgnd vpwr scs8hd_decap_3
XPHY_362 vgnd vpwr scs8hd_decap_3
XPHY_351 vgnd vpwr scs8hd_decap_3
XPHY_340 vgnd vpwr scs8hd_decap_3
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_86_80 vgnd vpwr scs8hd_decap_12
XFILLER_106_68 vgnd vpwr scs8hd_decap_12
XFILLER_103_114 vpwr vgnd scs8hd_fill_2
XFILLER_122_56 vgnd vpwr scs8hd_decap_12
XFILLER_82_27 vgnd vpwr scs8hd_decap_4
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
XFILLER_147_86 vgnd vpwr scs8hd_decap_12
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XFILLER_163_74 vgnd vpwr scs8hd_decap_12
XFILLER_176_117 vgnd vpwr scs8hd_decap_8
XFILLER_31_123 vpwr vgnd scs8hd_fill_2
XFILLER_72_93 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_decap_3
XFILLER_188_93 vgnd vpwr scs8hd_decap_12
XPHY_192 vgnd vpwr scs8hd_decap_3
XPHY_181 vgnd vpwr scs8hd_decap_3
XFILLER_100_117 vgnd vpwr scs8hd_decap_8
XFILLER_89_123 vpwr vgnd scs8hd_fill_2
XFILLER_77_27 vgnd vpwr scs8hd_decap_12
XFILLER_93_15 vgnd vpwr scs8hd_decap_12
XFILLER_165_3 vgnd vpwr scs8hd_decap_12
XFILLER_158_117 vgnd vpwr scs8hd_decap_8
XFILLER_93_59 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_80_3 vgnd vpwr scs8hd_decap_12
XFILLER_128_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_144_32 vgnd vpwr scs8hd_decap_12
XFILLER_77_115 vgnd vpwr scs8hd_decap_6
XFILLER_88_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_169_62 vgnd vpwr scs8hd_decap_12
XFILLER_169_51 vgnd vpwr scs8hd_decap_8
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_94_80 vgnd vpwr scs8hd_decap_12
XFILLER_114_68 vgnd vpwr scs8hd_decap_12
XPHY_769 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_758 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_747 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_736 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_725 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_714 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_703 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_56 vgnd vpwr scs8hd_decap_12
XFILLER_90_27 vgnd vpwr scs8hd_decap_4
XFILLER_151_123 vpwr vgnd scs8hd_fill_2
XFILLER_139_98 vgnd vpwr scs8hd_decap_12
XFILLER_128_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_98 vpwr vgnd scs8hd_fill_2
XFILLER_155_86 vgnd vpwr scs8hd_decap_12
XFILLER_171_74 vgnd vpwr scs8hd_decap_12
XFILLER_80_93 vgnd vpwr scs8hd_decap_12
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_100_15 vgnd vpwr scs8hd_decap_12
XFILLER_133_123 vpwr vgnd scs8hd_fill_2
XFILLER_69_39 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _10_/X vgnd vpwr scs8hd_diode_2
XFILLER_85_27 vgnd vpwr scs8hd_decap_12
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_599 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_588 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_577 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_566 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
XFILLER_115_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_118 vgnd vpwr scs8hd_decap_4
XFILLER_136_44 vgnd vpwr scs8hd_decap_12
XFILLER_96_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_152_32 vgnd vpwr scs8hd_decap_12
XPHY_352 vgnd vpwr scs8hd_decap_3
XPHY_341 vgnd vpwr scs8hd_decap_3
XPHY_330 vgnd vpwr scs8hd_decap_3
XFILLER_43_110 vgnd vpwr scs8hd_decap_12
XFILLER_45_74 vgnd vpwr scs8hd_decap_12
XPHY_374 vgnd vpwr scs8hd_decap_3
XPHY_363 vgnd vpwr scs8hd_decap_3
XFILLER_177_62 vgnd vpwr scs8hd_decap_12
XFILLER_177_51 vgnd vpwr scs8hd_decap_8
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_122_68 vgnd vpwr scs8hd_decap_12
XFILLER_25_110 vgnd vpwr scs8hd_decap_12
XFILLER_110_3 vgnd vpwr scs8hd_decap_12
XFILLER_147_98 vgnd vpwr scs8hd_decap_12
XFILLER_163_86 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_decap_3
XPHY_182 vgnd vpwr scs8hd_decap_3
XPHY_160 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_decap_3
XFILLER_22_102 vpwr vgnd scs8hd_fill_2
XFILLER_22_124 vgnd vpwr scs8hd_fill_1
XFILLER_77_39 vgnd vpwr scs8hd_decap_12
XFILLER_93_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_158_3 vgnd vpwr scs8hd_decap_12
XFILLER_181_110 vgnd vpwr scs8hd_decap_12
XFILLER_73_3 vgnd vpwr scs8hd_decap_12
XFILLER_86_105 vgnd vpwr scs8hd_decap_12
XFILLER_103_15 vgnd vpwr scs8hd_decap_12
XFILLER_103_59 vpwr vgnd scs8hd_fill_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_163_110 vgnd vpwr scs8hd_decap_12
XFILLER_128_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_88_27 vgnd vpwr scs8hd_decap_4
XFILLER_144_44 vgnd vpwr scs8hd_decap_12
XFILLER_160_32 vgnd vpwr scs8hd_decap_12
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_169_74 vgnd vpwr scs8hd_decap_12
XFILLER_53_74 vgnd vpwr scs8hd_decap_12
XFILLER_185_62 vgnd vpwr scs8hd_decap_12
XFILLER_185_51 vgnd vpwr scs8hd_decap_8
XFILLER_68_105 vgnd vpwr scs8hd_fill_1
XFILLER_78_93 vgnd vpwr scs8hd_decap_12
XFILLER_145_110 vgnd vpwr scs8hd_decap_12
XPHY_759 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_748 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_737 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_726 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_715 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_704 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_66 vgnd vpwr scs8hd_fill_1
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_99_59 vpwr vgnd scs8hd_fill_2
XFILLER_99_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_171_86 vgnd vpwr scs8hd_decap_12
XFILLER_155_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_104_80 vgnd vpwr scs8hd_decap_12
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_100_27 vgnd vpwr scs8hd_decap_4
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_85_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_140_3 vgnd vpwr scs8hd_decap_12
XFILLER_109_110 vgnd vpwr scs8hd_decap_12
XPHY_589 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_578 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_567 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_130_105 vgnd vpwr scs8hd_decap_12
XFILLER_111_59 vpwr vgnd scs8hd_fill_2
XFILLER_111_15 vgnd vpwr scs8hd_decap_12
XFILLER_136_56 vgnd vpwr scs8hd_decap_12
XFILLER_96_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_188_3 vgnd vpwr scs8hd_decap_12
XFILLER_152_44 vgnd vpwr scs8hd_decap_12
XFILLER_188_105 vgnd vpwr scs8hd_decap_12
XPHY_375 vgnd vpwr scs8hd_decap_3
XPHY_364 vgnd vpwr scs8hd_decap_3
XPHY_353 vgnd vpwr scs8hd_decap_3
XPHY_342 vgnd vpwr scs8hd_decap_3
XPHY_331 vgnd vpwr scs8hd_decap_3
XPHY_320 vgnd vpwr scs8hd_decap_3
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_45_86 vgnd vpwr scs8hd_decap_12
XFILLER_177_74 vgnd vpwr scs8hd_decap_12
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XFILLER_112_105 vgnd vpwr scs8hd_decap_12
XFILLER_86_93 vgnd vpwr scs8hd_decap_12
XFILLER_106_15 vgnd vpwr scs8hd_decap_12
XANTENNA__04__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_163_98 vgnd vpwr scs8hd_decap_12
XFILLER_103_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_111 vgnd vpwr scs8hd_decap_12
XFILLER_112_80 vgnd vpwr scs8hd_decap_12
XPHY_194 vgnd vpwr scs8hd_decap_3
XPHY_183 vgnd vpwr scs8hd_decap_3
XPHY_150 vgnd vpwr scs8hd_decap_3
XPHY_161 vgnd vpwr scs8hd_decap_3
XPHY_172 vgnd vpwr scs8hd_decap_3
XFILLER_93_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_158_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vgnd vpwr scs8hd_decap_4
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_67_51 vgnd vpwr scs8hd_decap_8
XFILLER_67_62 vgnd vpwr scs8hd_decap_12
XFILLER_66_3 vgnd vpwr scs8hd_decap_12
XFILLER_86_117 vgnd vpwr scs8hd_decap_8
XFILLER_103_27 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_8
XFILLER_128_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_144_56 vgnd vpwr scs8hd_decap_12
XFILLER_170_3 vgnd vpwr scs8hd_decap_12
XFILLER_160_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_169_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_53_86 vgnd vpwr scs8hd_decap_12
XFILLER_185_74 vgnd vpwr scs8hd_decap_12
XFILLER_94_93 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_8_ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_ebufn_1
XFILLER_114_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XPHY_727 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_716 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_705 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_749 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_738 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_99_27 vgnd vpwr scs8hd_decap_12
XANTENNA__12__A _12_/A vgnd vpwr scs8hd_diode_2
XFILLER_171_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_120_80 vgnd vpwr scs8hd_decap_12
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_109_59 vpwr vgnd scs8hd_fill_2
XFILLER_109_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XPHY_568 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__07__A _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_32 vgnd vpwr scs8hd_decap_12
XFILLER_133_3 vgnd vpwr scs8hd_decap_12
XPHY_579 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
XFILLER_59_74 vgnd vpwr scs8hd_decap_12
XFILLER_61_123 vpwr vgnd scs8hd_fill_2
XFILLER_75_51 vgnd vpwr scs8hd_decap_8
XFILLER_75_62 vgnd vpwr scs8hd_decap_12
XFILLER_130_117 vgnd vpwr scs8hd_decap_8
XFILLER_111_27 vgnd vpwr scs8hd_decap_12
XFILLER_136_68 vgnd vpwr scs8hd_decap_12
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_152_56 vgnd vpwr scs8hd_decap_12
XFILLER_43_123 vpwr vgnd scs8hd_fill_2
XFILLER_188_117 vgnd vpwr scs8hd_decap_8
XPHY_376 vgnd vpwr scs8hd_decap_3
XPHY_365 vgnd vpwr scs8hd_decap_3
XPHY_354 vgnd vpwr scs8hd_decap_3
XPHY_343 vgnd vpwr scs8hd_decap_3
XPHY_332 vgnd vpwr scs8hd_decap_3
XPHY_321 vgnd vpwr scs8hd_decap_3
XPHY_310 vgnd vpwr scs8hd_decap_3
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_45_98 vgnd vpwr scs8hd_decap_6
XFILLER_61_86 vgnd vpwr scs8hd_decap_12
XFILLER_177_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_112_117 vgnd vpwr scs8hd_decap_8
XFILLER_96_3 vgnd vpwr scs8hd_decap_12
XFILLER_106_27 vgnd vpwr scs8hd_decap_4
XFILLER_122_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_101 vgnd vpwr scs8hd_decap_3
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XANTENNA__20__A gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_123 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_decap_3
XPHY_184 vgnd vpwr scs8hd_decap_3
XPHY_140 vgnd vpwr scs8hd_decap_3
XPHY_151 vgnd vpwr scs8hd_decap_3
XPHY_162 vgnd vpwr scs8hd_decap_3
XPHY_173 vgnd vpwr scs8hd_decap_3
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_117_15 vgnd vpwr scs8hd_decap_12
XFILLER_117_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_158_44 vgnd vpwr scs8hd_decap_12
XANTENNA__15__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_181_123 vpwr vgnd scs8hd_fill_2
XFILLER_174_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_67_74 vgnd vpwr scs8hd_decap_12
XFILLER_83_51 vgnd vpwr scs8hd_decap_8
XFILLER_83_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XFILLER_103_39 vgnd vpwr scs8hd_decap_12
XFILLER_163_123 vpwr vgnd scs8hd_fill_2
XFILLER_144_68 vgnd vpwr scs8hd_decap_12
XFILLER_163_3 vgnd vpwr scs8hd_decap_12
XFILLER_160_56 vgnd vpwr scs8hd_decap_12
XFILLER_169_98 vgnd vpwr scs8hd_decap_8
XFILLER_53_98 vgnd vpwr scs8hd_decap_12
XFILLER_185_86 vgnd vpwr scs8hd_decap_12
XFILLER_118_80 vgnd vpwr scs8hd_decap_12
XFILLER_91_110 vgnd vpwr scs8hd_decap_12
XFILLER_145_123 vpwr vgnd scs8hd_fill_2
XFILLER_114_27 vgnd vpwr scs8hd_decap_4
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _12_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_739 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_728 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_717 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_706 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_15 vgnd vpwr scs8hd_decap_12
XFILLER_99_39 vgnd vpwr scs8hd_decap_12
XANTENNA__12__B _13_/B vgnd vpwr scs8hd_diode_2
XFILLER_151_115 vgnd vpwr scs8hd_decap_6
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
XFILLER_104_93 vgnd vpwr scs8hd_decap_12
XFILLER_73_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_127_123 vpwr vgnd scs8hd_fill_2
XFILLER_109_27 vgnd vpwr scs8hd_decap_12
XFILLER_125_59 vpwr vgnd scs8hd_fill_2
XFILLER_125_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_55_110 vgnd vpwr scs8hd_decap_12
XPHY_569 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__07__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_44 vgnd vpwr scs8hd_decap_12
XFILLER_126_3 vgnd vpwr scs8hd_decap_12
XFILLER_109_123 vpwr vgnd scs8hd_fill_2
XANTENNA__23__A gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_diode_2
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XFILLER_182_32 vgnd vpwr scs8hd_decap_12
XFILLER_59_86 vgnd vpwr scs8hd_decap_12
XFILLER_91_51 vgnd vpwr scs8hd_decap_8
XFILLER_75_74 vgnd vpwr scs8hd_decap_12
XFILLER_91_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_111_39 vgnd vpwr scs8hd_decap_12
XANTENNA__18__A gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_diode_2
XFILLER_152_68 vgnd vpwr scs8hd_decap_12
XPHY_300 vgnd vpwr scs8hd_decap_3
XFILLER_28_121 vgnd vpwr scs8hd_decap_4
XPHY_377 vgnd vpwr scs8hd_decap_3
XPHY_366 vgnd vpwr scs8hd_decap_3
XPHY_355 vgnd vpwr scs8hd_decap_3
XPHY_344 vgnd vpwr scs8hd_decap_3
XPHY_333 vgnd vpwr scs8hd_decap_3
XPHY_322 vgnd vpwr scs8hd_decap_3
XPHY_311 vgnd vpwr scs8hd_decap_3
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XFILLER_177_98 vgnd vpwr scs8hd_decap_12
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_126_80 vgnd vpwr scs8hd_decap_12
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_89_3 vgnd vpwr scs8hd_decap_12
XFILLER_103_118 vgnd vpwr scs8hd_decap_4
XFILLER_122_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_112_93 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_decap_3
XPHY_141 vgnd vpwr scs8hd_decap_3
XPHY_152 vgnd vpwr scs8hd_decap_3
XPHY_196 vgnd vpwr scs8hd_decap_3
XPHY_185 vgnd vpwr scs8hd_decap_3
XPHY_163 vgnd vpwr scs8hd_decap_3
XPHY_174 vgnd vpwr scs8hd_decap_3
XFILLER_98_105 vgnd vpwr scs8hd_decap_12
XFILLER_117_27 vgnd vpwr scs8hd_decap_12
XFILLER_133_59 vpwr vgnd scs8hd_fill_2
XFILLER_133_15 vgnd vpwr scs8hd_decap_12
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_158_56 vgnd vpwr scs8hd_decap_12
XANTENNA__15__B _13_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XFILLER_174_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_190_32 vgnd vpwr scs8hd_decap_12
XFILLER_67_86 vgnd vpwr scs8hd_decap_12
XFILLER_157_110 vgnd vpwr scs8hd_decap_12
XFILLER_83_74 vgnd vpwr scs8hd_decap_12
XFILLER_128_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_160_68 vgnd vpwr scs8hd_decap_12
XFILLER_156_3 vgnd vpwr scs8hd_decap_12
XFILLER_139_110 vgnd vpwr scs8hd_decap_12
XFILLER_185_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_134_80 vgnd vpwr scs8hd_decap_12
XFILLER_68_108 vgnd vpwr scs8hd_decap_12
XFILLER_71_3 vgnd vpwr scs8hd_decap_12
XFILLER_160_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XPHY_729 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_718 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_707 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_27 vgnd vpwr scs8hd_decap_4
XFILLER_23_69 vpwr vgnd scs8hd_fill_2
XANTENNA__12__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_120_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_142_105 vgnd vpwr scs8hd_decap_12
XFILLER_89_62 vgnd vpwr scs8hd_decap_12
XFILLER_89_51 vgnd vpwr scs8hd_decap_8
XFILLER_109_39 vgnd vpwr scs8hd_decap_12
XFILLER_125_27 vgnd vpwr scs8hd_decap_12
XFILLER_141_59 vpwr vgnd scs8hd_fill_2
XFILLER_141_15 vgnd vpwr scs8hd_decap_12
XANTENNA__07__C _12_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_56 vgnd vpwr scs8hd_decap_12
XFILLER_124_105 vgnd vpwr scs8hd_decap_12
XFILLER_119_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_182_44 vgnd vpwr scs8hd_decap_12
XFILLER_59_98 vgnd vpwr scs8hd_decap_12
XFILLER_91_74 vgnd vpwr scs8hd_decap_12
XFILLER_75_86 vgnd vpwr scs8hd_decap_12
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_136_15 vgnd vpwr scs8hd_decap_12
XFILLER_106_105 vgnd vpwr scs8hd_decap_12
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XPHY_334 vgnd vpwr scs8hd_decap_3
XPHY_323 vgnd vpwr scs8hd_decap_3
XPHY_312 vgnd vpwr scs8hd_decap_3
XPHY_301 vgnd vpwr scs8hd_decap_3
XFILLER_101_51 vgnd vpwr scs8hd_decap_8
XPHY_378 vgnd vpwr scs8hd_decap_3
XPHY_367 vgnd vpwr scs8hd_decap_3
XPHY_356 vgnd vpwr scs8hd_decap_3
XPHY_345 vgnd vpwr scs8hd_decap_3
XFILLER_101_62 vgnd vpwr scs8hd_decap_12
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_142_80 vgnd vpwr scs8hd_decap_12
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_117 vgnd vpwr scs8hd_decap_8
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_186_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XFILLER_188_32 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_131 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_decap_3
XFILLER_72_32 vgnd vpwr scs8hd_decap_12
XPHY_153 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_decap_3
XPHY_175 vgnd vpwr scs8hd_decap_3
XPHY_197 vgnd vpwr scs8hd_decap_3
XPHY_186 vgnd vpwr scs8hd_decap_3
XFILLER_98_117 vgnd vpwr scs8hd_decap_8
XFILLER_97_62 vgnd vpwr scs8hd_decap_12
XFILLER_97_51 vgnd vpwr scs8hd_decap_8
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_106 vgnd vpwr scs8hd_decap_12
XFILLER_117_39 vgnd vpwr scs8hd_decap_12
XFILLER_133_27 vgnd vpwr scs8hd_decap_12
XANTENNA__15__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_158_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
XFILLER_174_56 vgnd vpwr scs8hd_decap_12
XFILLER_101_3 vgnd vpwr scs8hd_decap_12
XFILLER_190_44 vgnd vpwr scs8hd_decap_12
XFILLER_67_98 vgnd vpwr scs8hd_decap_12
XFILLER_83_86 vgnd vpwr scs8hd_decap_12
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XFILLER_16_80 vgnd vpwr scs8hd_decap_3
XFILLER_128_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_144_15 vgnd vpwr scs8hd_decap_12
XFILLER_149_3 vgnd vpwr scs8hd_decap_12
XFILLER_118_93 vgnd vpwr scs8hd_decap_12
XFILLER_150_80 vgnd vpwr scs8hd_decap_12
XFILLER_91_123 vpwr vgnd scs8hd_fill_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_160_117 vgnd vpwr scs8hd_decap_8
XPHY_719 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_708 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_139_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_139_59 vpwr vgnd scs8hd_fill_2
XANTENNA__12__D _13_/D vgnd vpwr scs8hd_diode_2
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_73_123 vpwr vgnd scs8hd_fill_2
XFILLER_127_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_80_32 vgnd vpwr scs8hd_decap_12
XFILLER_142_117 vgnd vpwr scs8hd_decap_8
XFILLER_89_74 vgnd vpwr scs8hd_decap_12
XFILLER_125_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_141_27 vgnd vpwr scs8hd_decap_12
XANTENNA__07__D enable vgnd vpwr scs8hd_diode_2
XFILLER_55_123 vpwr vgnd scs8hd_fill_2
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_68 vgnd vpwr scs8hd_decap_12
XFILLER_124_117 vgnd vpwr scs8hd_decap_8
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XFILLER_182_56 vgnd vpwr scs8hd_decap_12
XFILLER_75_98 vgnd vpwr scs8hd_decap_12
XFILLER_91_86 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vpwr vgnd scs8hd_fill_2
XFILLER_136_27 vgnd vpwr scs8hd_decap_4
XFILLER_106_117 vgnd vpwr scs8hd_decap_8
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_152_15 vgnd vpwr scs8hd_decap_12
XPHY_368 vgnd vpwr scs8hd_decap_3
XPHY_357 vgnd vpwr scs8hd_decap_3
XPHY_346 vgnd vpwr scs8hd_decap_3
XPHY_335 vgnd vpwr scs8hd_decap_3
XPHY_324 vgnd vpwr scs8hd_decap_3
XPHY_313 vgnd vpwr scs8hd_decap_3
XPHY_302 vgnd vpwr scs8hd_decap_3
XFILLER_101_74 vgnd vpwr scs8hd_decap_12
XPHY_379 vgnd vpwr scs8hd_decap_3
XFILLER_131_3 vgnd vpwr scs8hd_decap_12
XFILLER_126_93 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
X_09_ address[1] enable address[3] _13_/D _09_/X vgnd vpwr scs8hd_and4_4
XFILLER_147_59 vpwr vgnd scs8hd_fill_2
XFILLER_147_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_179_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
XFILLER_188_44 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_decap_3
XPHY_187 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_132 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_decap_3
XFILLER_72_44 vgnd vpwr scs8hd_decap_12
XPHY_154 vgnd vpwr scs8hd_decap_3
XPHY_165 vgnd vpwr scs8hd_decap_3
XPHY_176 vgnd vpwr scs8hd_decap_3
XFILLER_97_74 vgnd vpwr scs8hd_decap_12
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_118 vgnd vpwr scs8hd_decap_6
XFILLER_175_123 vpwr vgnd scs8hd_fill_2
XFILLER_94_3 vgnd vpwr scs8hd_decap_12
XFILLER_133_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA__15__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_190_56 vgnd vpwr scs8hd_decap_12
XFILLER_174_68 vgnd vpwr scs8hd_decap_12
XFILLER_107_62 vgnd vpwr scs8hd_decap_12
XFILLER_107_51 vgnd vpwr scs8hd_decap_8
XFILLER_83_98 vgnd vpwr scs8hd_decap_12
XFILLER_157_123 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_148_80 vgnd vpwr scs8hd_decap_12
XFILLER_144_27 vgnd vpwr scs8hd_decap_4
XFILLER_85_110 vgnd vpwr scs8hd_decap_12
XFILLER_160_15 vgnd vpwr scs8hd_decap_12
XFILLER_139_123 vpwr vgnd scs8hd_fill_2
XFILLER_78_32 vgnd vpwr scs8hd_decap_12
XFILLER_134_93 vgnd vpwr scs8hd_decap_12
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_67_110 vgnd vpwr scs8hd_decap_12
XPHY_709 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_139_27 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_155_59 vpwr vgnd scs8hd_fill_2
XFILLER_155_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
XFILLER_161_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_56 vgnd vpwr scs8hd_decap_12
XFILLER_80_44 vgnd vpwr scs8hd_decap_12
XFILLER_89_86 vgnd vpwr scs8hd_decap_12
XFILLER_49_110 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_141_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_105 vgnd vpwr scs8hd_decap_12
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_182_68 vgnd vpwr scs8hd_decap_12
XFILLER_115_62 vgnd vpwr scs8hd_decap_12
XFILLER_115_51 vgnd vpwr scs8hd_decap_8
XFILLER_91_98 vgnd vpwr scs8hd_decap_12
XFILLER_156_80 vgnd vpwr scs8hd_decap_12
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vgnd vpwr scs8hd_fill_1
XFILLER_52_105 vgnd vpwr scs8hd_decap_12
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_152_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XPHY_369 vgnd vpwr scs8hd_decap_3
XPHY_358 vgnd vpwr scs8hd_decap_3
XPHY_347 vgnd vpwr scs8hd_decap_3
XPHY_336 vgnd vpwr scs8hd_decap_3
XPHY_325 vgnd vpwr scs8hd_decap_3
XPHY_314 vgnd vpwr scs8hd_decap_3
XPHY_303 vgnd vpwr scs8hd_decap_3
XFILLER_101_86 vgnd vpwr scs8hd_decap_12
XFILLER_124_3 vgnd vpwr scs8hd_decap_12
XFILLER_86_32 vgnd vpwr scs8hd_decap_12
XFILLER_142_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_187_110 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_10_ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_ebufn_1
XFILLER_111_110 vgnd vpwr scs8hd_decap_12
X_08_ address[2] _13_/D vgnd vpwr scs8hd_inv_8
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_147_27 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_163_59 vpwr vgnd scs8hd_fill_2
XFILLER_163_15 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XFILLER_188_56 vgnd vpwr scs8hd_decap_12
XFILLER_169_121 vgnd vpwr scs8hd_fill_1
XPHY_199 vgnd vpwr scs8hd_decap_3
XPHY_188 vgnd vpwr scs8hd_decap_3
XFILLER_31_119 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_133 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_decap_3
XFILLER_72_56 vgnd vpwr scs8hd_decap_12
XPHY_155 vgnd vpwr scs8hd_decap_3
XPHY_166 vgnd vpwr scs8hd_decap_3
XPHY_177 vgnd vpwr scs8hd_decap_3
XFILLER_97_86 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_190_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_87_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_158_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_191_3 vgnd vpwr scs8hd_decap_12
XFILLER_190_68 vgnd vpwr scs8hd_decap_12
XFILLER_123_62 vgnd vpwr scs8hd_decap_12
XFILLER_123_51 vgnd vpwr scs8hd_decap_8
XFILLER_107_74 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_6
XFILLER_172_105 vgnd vpwr scs8hd_decap_12
XFILLER_164_80 vgnd vpwr scs8hd_decap_12
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_160_27 vgnd vpwr scs8hd_decap_4
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_154_105 vgnd vpwr scs8hd_decap_12
XFILLER_78_44 vgnd vpwr scs8hd_decap_12
XFILLER_94_32 vgnd vpwr scs8hd_decap_12
XFILLER_150_93 vgnd vpwr scs8hd_decap_12
XFILLER_139_39 vgnd vpwr scs8hd_decap_12
XFILLER_136_105 vgnd vpwr scs8hd_decap_12
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_155_27 vgnd vpwr scs8hd_decap_12
XFILLER_171_59 vpwr vgnd scs8hd_fill_2
XFILLER_171_15 vgnd vpwr scs8hd_decap_12
XFILLER_154_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_68 vgnd vpwr scs8hd_decap_12
XFILLER_80_56 vgnd vpwr scs8hd_decap_12
XFILLER_89_98 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_118_105 vgnd vpwr scs8hd_decap_4
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_117 vgnd vpwr scs8hd_decap_8
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_15 vgnd vpwr scs8hd_decap_12
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_131_62 vgnd vpwr scs8hd_decap_12
XFILLER_131_51 vgnd vpwr scs8hd_decap_8
XFILLER_115_74 vgnd vpwr scs8hd_decap_12
XFILLER_172_80 vgnd vpwr scs8hd_decap_12
XFILLER_52_117 vgnd vpwr scs8hd_decap_8
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
XPHY_359 vgnd vpwr scs8hd_decap_3
XPHY_348 vgnd vpwr scs8hd_decap_3
XPHY_337 vgnd vpwr scs8hd_decap_3
XPHY_326 vgnd vpwr scs8hd_decap_3
XPHY_315 vgnd vpwr scs8hd_decap_3
XPHY_304 vgnd vpwr scs8hd_decap_3
XFILLER_101_98 vgnd vpwr scs8hd_decap_12
XFILLER_117_3 vgnd vpwr scs8hd_decap_12
XFILLER_86_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_117 vgnd vpwr scs8hd_decap_8
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
X_07_ _13_/C address[2] _12_/A enable _07_/X vgnd vpwr scs8hd_and4_4
XFILLER_25_106 vpwr vgnd scs8hd_fill_2
XFILLER_147_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_163_27 vgnd vpwr scs8hd_decap_12
XFILLER_169_111 vpwr vgnd scs8hd_fill_2
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_decap_3
XFILLER_72_68 vgnd vpwr scs8hd_decap_12
XFILLER_188_68 vgnd vpwr scs8hd_decap_12
XPHY_189 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_decap_3
XPHY_156 vgnd vpwr scs8hd_decap_3
XPHY_167 vgnd vpwr scs8hd_decap_3
XPHY_178 vgnd vpwr scs8hd_decap_3
XFILLER_97_98 vgnd vpwr scs8hd_decap_12
XFILLER_175_114 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_46_80 vgnd vpwr scs8hd_decap_12
XFILLER_190_117 vgnd vpwr scs8hd_decap_8
XPHY_690 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XFILLER_158_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_174_15 vgnd vpwr scs8hd_decap_12
XFILLER_184_3 vgnd vpwr scs8hd_decap_12
XFILLER_123_74 vgnd vpwr scs8hd_decap_12
XFILLER_107_86 vgnd vpwr scs8hd_decap_12
XFILLER_172_117 vgnd vpwr scs8hd_decap_8
XFILLER_148_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_180_80 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_85_123 vpwr vgnd scs8hd_fill_2
XFILLER_169_59 vpwr vgnd scs8hd_fill_2
XFILLER_169_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_154_117 vgnd vpwr scs8hd_decap_8
XFILLER_78_56 vgnd vpwr scs8hd_decap_12
XFILLER_94_44 vgnd vpwr scs8hd_decap_12
XFILLER_67_123 vpwr vgnd scs8hd_fill_2
XFILLER_136_117 vgnd vpwr scs8hd_decap_8
XFILLER_171_27 vgnd vpwr scs8hd_decap_12
XFILLER_155_39 vgnd vpwr scs8hd_decap_12
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_104_32 vgnd vpwr scs8hd_decap_12
XFILLER_147_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_80_68 vgnd vpwr scs8hd_decap_12
XFILLER_129_62 vgnd vpwr scs8hd_decap_12
XFILLER_129_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_49_123 vpwr vgnd scs8hd_fill_2
XFILLER_54_80 vgnd vpwr scs8hd_decap_12
XFILLER_118_117 vgnd vpwr scs8hd_decap_8
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_27 vgnd vpwr scs8hd_decap_4
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XFILLER_182_15 vgnd vpwr scs8hd_decap_12
XFILLER_115_86 vgnd vpwr scs8hd_decap_12
XFILLER_131_74 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
XFILLER_156_93 vgnd vpwr scs8hd_decap_12
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_23_ gfpga_pad_GPIO_PAD[4] right_width_0_height_0__pin_9_ vgnd vpwr scs8hd_buf_2
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _12_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XPHY_316 vgnd vpwr scs8hd_decap_3
XPHY_305 vgnd vpwr scs8hd_decap_3
XFILLER_45_27 vgnd vpwr scs8hd_decap_12
XFILLER_177_59 vpwr vgnd scs8hd_fill_2
XFILLER_177_15 vgnd vpwr scs8hd_decap_12
XPHY_349 vgnd vpwr scs8hd_decap_3
XPHY_338 vgnd vpwr scs8hd_decap_3
XPHY_327 vgnd vpwr scs8hd_decap_3
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vgnd vpwr scs8hd_decap_6
XFILLER_86_56 vgnd vpwr scs8hd_decap_12
XFILLER_187_123 vpwr vgnd scs8hd_fill_2
XFILLER_111_123 vpwr vgnd scs8hd_fill_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_06_ address[1] _12_/A vgnd vpwr scs8hd_inv_8
XFILLER_163_39 vgnd vpwr scs8hd_decap_12
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XFILLER_169_123 vpwr vgnd scs8hd_fill_2
XFILLER_112_32 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_135 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_decap_3
XPHY_157 vgnd vpwr scs8hd_decap_3
XPHY_179 vgnd vpwr scs8hd_decap_3
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XPHY_168 vgnd vpwr scs8hd_decap_3
XFILLER_137_62 vgnd vpwr scs8hd_decap_12
XFILLER_137_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XFILLER_178_80 vgnd vpwr scs8hd_decap_12
XPHY_691 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_680 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_97_110 vgnd vpwr scs8hd_decap_12
XFILLER_190_15 vgnd vpwr scs8hd_decap_12
XFILLER_174_27 vgnd vpwr scs8hd_decap_4
XFILLER_107_98 vgnd vpwr scs8hd_decap_12
XFILLER_177_3 vgnd vpwr scs8hd_decap_12
XFILLER_123_86 vgnd vpwr scs8hd_decap_12
XFILLER_164_93 vgnd vpwr scs8hd_decap_12
XFILLER_79_110 vgnd vpwr scs8hd_decap_12
XFILLER_92_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_169_27 vgnd vpwr scs8hd_decap_12
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
XFILLER_185_59 vpwr vgnd scs8hd_fill_2
XFILLER_185_15 vgnd vpwr scs8hd_decap_12
XFILLER_78_68 vgnd vpwr scs8hd_decap_12
XFILLER_94_56 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_82_105 vgnd vpwr scs8hd_decap_12
XFILLER_2_109 vgnd vpwr scs8hd_decap_12
XFILLER_171_39 vgnd vpwr scs8hd_decap_12
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XFILLER_120_32 vgnd vpwr scs8hd_decap_12
XFILLER_104_44 vgnd vpwr scs8hd_decap_12
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XFILLER_127_118 vgnd vpwr scs8hd_decap_4
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_145_62 vgnd vpwr scs8hd_decap_12
XFILLER_145_51 vgnd vpwr scs8hd_decap_8
XFILLER_129_74 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_64_105 vgnd vpwr scs8hd_decap_12
XFILLER_186_80 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _05_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XFILLER_70_80 vgnd vpwr scs8hd_decap_12
XFILLER_141_110 vgnd vpwr scs8hd_decap_12
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_182_27 vgnd vpwr scs8hd_decap_4
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_115_98 vgnd vpwr scs8hd_decap_12
XFILLER_46_105 vgnd vpwr scs8hd_decap_12
XFILLER_131_86 vgnd vpwr scs8hd_decap_12
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_123_110 vgnd vpwr scs8hd_decap_12
XFILLER_172_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
X_22_ gfpga_pad_GPIO_PAD[3] right_width_0_height_0__pin_7_ vgnd vpwr scs8hd_buf_2
XPHY_339 vgnd vpwr scs8hd_decap_3
XPHY_328 vgnd vpwr scs8hd_decap_3
XPHY_317 vgnd vpwr scs8hd_decap_3
XPHY_306 vgnd vpwr scs8hd_decap_3
XFILLER_45_39 vgnd vpwr scs8hd_decap_12
XFILLER_177_27 vgnd vpwr scs8hd_decap_12
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_105_110 vgnd vpwr scs8hd_decap_12
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_86_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
X_05_ _13_/C address[2] address[1] enable _05_/X vgnd vpwr scs8hd_and4_4
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_188_15 vgnd vpwr scs8hd_decap_12
XFILLER_184_105 vgnd vpwr scs8hd_decap_12
XFILLER_112_44 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_136 vgnd vpwr scs8hd_decap_3
XFILLER_72_15 vgnd vpwr scs8hd_decap_12
XPHY_147 vgnd vpwr scs8hd_decap_3
XPHY_158 vgnd vpwr scs8hd_decap_3
XPHY_169 vgnd vpwr scs8hd_decap_3
XFILLER_137_74 vgnd vpwr scs8hd_decap_12
XFILLER_122_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_74 vgnd vpwr scs8hd_fill_1
XFILLER_153_62 vgnd vpwr scs8hd_decap_12
XFILLER_153_51 vgnd vpwr scs8hd_decap_8
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_46_93 vgnd vpwr scs8hd_decap_12
XPHY_692 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_681 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_670 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_166_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_111 vgnd vpwr scs8hd_decap_8
XFILLER_190_27 vgnd vpwr scs8hd_decap_4
XFILLER_67_15 vgnd vpwr scs8hd_decap_12
XFILLER_67_59 vpwr vgnd scs8hd_fill_2
XFILLER_123_98 vgnd vpwr scs8hd_decap_12
XFILLER_16_85 vgnd vpwr scs8hd_decap_6
XFILLER_180_93 vgnd vpwr scs8hd_decap_12
XFILLER_148_105 vgnd vpwr scs8hd_decap_12
XFILLER_85_3 vgnd vpwr scs8hd_decap_12
XFILLER_169_39 vgnd vpwr scs8hd_decap_12
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
XFILLER_185_27 vgnd vpwr scs8hd_decap_12
XFILLER_118_32 vgnd vpwr scs8hd_decap_12
XFILLER_94_68 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_68_80 vgnd vpwr scs8hd_decap_12
XFILLER_82_117 vgnd vpwr scs8hd_decap_8
XFILLER_120_44 vgnd vpwr scs8hd_decap_12
XFILLER_104_56 vgnd vpwr scs8hd_decap_12
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_80_15 vgnd vpwr scs8hd_decap_12
XFILLER_145_74 vgnd vpwr scs8hd_decap_12
XFILLER_129_86 vgnd vpwr scs8hd_decap_12
XFILLER_161_62 vgnd vpwr scs8hd_decap_12
XFILLER_161_51 vgnd vpwr scs8hd_decap_8
XFILLER_64_117 vgnd vpwr scs8hd_decap_8
XFILLER_54_93 vgnd vpwr scs8hd_decap_12
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XFILLER_46_117 vgnd vpwr scs8hd_decap_8
XFILLER_75_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_59 vpwr vgnd scs8hd_fill_2
XFILLER_152_3 vgnd vpwr scs8hd_decap_12
XFILLER_131_98 vgnd vpwr scs8hd_decap_12
XFILLER_24_74 vgnd vpwr scs8hd_fill_1
X_21_ gfpga_pad_GPIO_PAD[2] right_width_0_height_0__pin_5_ vgnd vpwr scs8hd_buf_2
XPHY_329 vgnd vpwr scs8hd_decap_3
XPHY_318 vgnd vpwr scs8hd_decap_3
XPHY_307 vgnd vpwr scs8hd_decap_3
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_177_39 vgnd vpwr scs8hd_decap_12
XFILLER_126_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_85 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _13_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_04_ address[3] _13_/C vgnd vpwr scs8hd_buf_1
XFILLER_76_80 vgnd vpwr scs8hd_decap_12
XFILLER_112_56 vgnd vpwr scs8hd_decap_12
XFILLER_188_27 vgnd vpwr scs8hd_decap_4
XFILLER_184_117 vgnd vpwr scs8hd_decap_8
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_137 vgnd vpwr scs8hd_decap_3
XFILLER_72_27 vgnd vpwr scs8hd_decap_4
XPHY_148 vgnd vpwr scs8hd_decap_3
XPHY_159 vgnd vpwr scs8hd_decap_3
XFILLER_137_86 vgnd vpwr scs8hd_decap_12
XFILLER_115_3 vgnd vpwr scs8hd_decap_12
XFILLER_153_74 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_178_93 vgnd vpwr scs8hd_decap_12
XPHY_693 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_682 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_671 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_660 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_123 vpwr vgnd scs8hd_fill_2
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XFILLER_97_123 vpwr vgnd scs8hd_fill_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_166_117 vgnd vpwr scs8hd_decap_8
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_67_27 vgnd vpwr scs8hd_decap_12
XFILLER_83_15 vgnd vpwr scs8hd_decap_12
XFILLER_83_59 vpwr vgnd scs8hd_fill_2
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_79_123 vpwr vgnd scs8hd_fill_2
XFILLER_148_117 vgnd vpwr scs8hd_decap_8
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_78_3 vgnd vpwr scs8hd_decap_12
XFILLER_185_39 vgnd vpwr scs8hd_decap_12
XFILLER_118_44 vgnd vpwr scs8hd_decap_12
XFILLER_78_15 vgnd vpwr scs8hd_decap_12
XFILLER_182_3 vgnd vpwr scs8hd_decap_12
XFILLER_134_32 vgnd vpwr scs8hd_decap_12
XFILLER_27_74 vpwr vgnd scs8hd_fill_2
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XFILLER_159_62 vgnd vpwr scs8hd_decap_12
XFILLER_159_51 vgnd vpwr scs8hd_decap_8
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_12_ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_ebufn_1
XFILLER_84_80 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_104_68 vgnd vpwr scs8hd_decap_12
XFILLER_120_56 vgnd vpwr scs8hd_decap_12
XFILLER_80_27 vgnd vpwr scs8hd_decap_4
XFILLER_129_98 vgnd vpwr scs8hd_decap_12
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_145_86 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_161_74 vgnd vpwr scs8hd_decap_12
XFILLER_186_93 vgnd vpwr scs8hd_decap_12
XFILLER_141_123 vpwr vgnd scs8hd_fill_2
XFILLER_70_93 vgnd vpwr scs8hd_decap_12
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
XFILLER_91_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_27 vgnd vpwr scs8hd_decap_12
XFILLER_145_3 vgnd vpwr scs8hd_decap_12
XFILLER_91_59 vpwr vgnd scs8hd_fill_2
XFILLER_123_123 vpwr vgnd scs8hd_fill_2
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_20_ gfpga_pad_GPIO_PAD[1] right_width_0_height_0__pin_3_ vgnd vpwr scs8hd_buf_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XPHY_319 vgnd vpwr scs8hd_decap_3
XPHY_308 vgnd vpwr scs8hd_decap_3
XFILLER_51_110 vgnd vpwr scs8hd_decap_12
XFILLER_105_123 vpwr vgnd scs8hd_fill_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_142_32 vgnd vpwr scs8hd_decap_12
XFILLER_126_44 vgnd vpwr scs8hd_decap_12
XFILLER_86_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_97 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_167_62 vgnd vpwr scs8hd_decap_12
XFILLER_167_51 vgnd vpwr scs8hd_decap_8
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
XFILLER_92_80 vgnd vpwr scs8hd_decap_12
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XFILLER_169_115 vgnd vpwr scs8hd_decap_6
XFILLER_112_68 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_decap_3
XPHY_116 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_138 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_decap_3
XFILLER_137_98 vgnd vpwr scs8hd_decap_12
XFILLER_108_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_87 vgnd vpwr scs8hd_decap_6
XFILLER_153_86 vgnd vpwr scs8hd_decap_12
XPHY_661 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_650 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XFILLER_175_118 vgnd vpwr scs8hd_decap_4
XPHY_694 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_683 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_672 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _05_/X vgnd vpwr scs8hd_diode_2
XFILLER_67_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_83_27 vgnd vpwr scs8hd_decap_12
XFILLER_8_117 vgnd vpwr scs8hd_decap_8
XFILLER_94_105 vgnd vpwr scs8hd_decap_4
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_171_110 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_134_44 vgnd vpwr scs8hd_decap_12
XFILLER_118_56 vgnd vpwr scs8hd_decap_12
XFILLER_76_105 vgnd vpwr scs8hd_decap_12
XFILLER_78_27 vgnd vpwr scs8hd_decap_4
XFILLER_175_3 vgnd vpwr scs8hd_decap_12
XFILLER_150_32 vgnd vpwr scs8hd_decap_12
XFILLER_94_15 vgnd vpwr scs8hd_decap_12
XFILLER_159_74 vgnd vpwr scs8hd_decap_12
XFILLER_43_74 vgnd vpwr scs8hd_decap_12
XFILLER_175_62 vgnd vpwr scs8hd_decap_12
XFILLER_175_51 vgnd vpwr scs8hd_decap_8
XFILLER_153_110 vgnd vpwr scs8hd_decap_12
XFILLER_191_94 vgnd vpwr scs8hd_decap_12
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_68_93 vgnd vpwr scs8hd_decap_12
XFILLER_90_3 vgnd vpwr scs8hd_decap_12
XFILLER_58_105 vgnd vpwr scs8hd_decap_12
XFILLER_120_68 vgnd vpwr scs8hd_decap_12
XFILLER_135_110 vgnd vpwr scs8hd_decap_12
XFILLER_89_15 vgnd vpwr scs8hd_decap_12
XFILLER_89_59 vpwr vgnd scs8hd_fill_2
XFILLER_145_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_123 vpwr vgnd scs8hd_fill_2
XFILLER_161_86 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_117_121 vgnd vpwr scs8hd_fill_1
XFILLER_91_27 vgnd vpwr scs8hd_decap_12
XFILLER_75_39 vgnd vpwr scs8hd_decap_12
XFILLER_138_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XFILLER_101_15 vgnd vpwr scs8hd_decap_12
XPHY_309 vgnd vpwr scs8hd_decap_3
XFILLER_101_59 vpwr vgnd scs8hd_fill_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_142_44 vgnd vpwr scs8hd_decap_12
XFILLER_126_56 vgnd vpwr scs8hd_decap_12
XFILLER_120_105 vgnd vpwr scs8hd_decap_12
XFILLER_86_27 vgnd vpwr scs8hd_decap_4
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_167_74 vgnd vpwr scs8hd_decap_12
XFILLER_51_74 vgnd vpwr scs8hd_decap_12
XFILLER_183_62 vgnd vpwr scs8hd_decap_12
XFILLER_183_51 vgnd vpwr scs8hd_decap_8
XFILLER_76_93 vgnd vpwr scs8hd_decap_12
XFILLER_178_105 vgnd vpwr scs8hd_decap_12
XFILLER_102_105 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_decap_3
XFILLER_97_59 vpwr vgnd scs8hd_fill_2
XFILLER_97_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_77 vgnd vpwr scs8hd_decap_8
XFILLER_21_99 vgnd vpwr scs8hd_decap_12
XFILLER_153_98 vgnd vpwr scs8hd_decap_12
XPHY_695 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_684 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_673 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_662 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_651 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_640 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_80 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_83_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_99 vgnd vpwr scs8hd_fill_1
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_148_32 vgnd vpwr scs8hd_decap_12
XFILLER_120_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_94_117 vgnd vpwr scs8hd_decap_8
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_98_80 vgnd vpwr scs8hd_decap_12
XFILLER_134_56 vgnd vpwr scs8hd_decap_12
XFILLER_118_68 vgnd vpwr scs8hd_decap_12
XFILLER_94_27 vgnd vpwr scs8hd_decap_4
XFILLER_76_117 vgnd vpwr scs8hd_decap_8
XFILLER_168_3 vgnd vpwr scs8hd_decap_12
XFILLER_150_44 vgnd vpwr scs8hd_decap_12
XFILLER_159_86 vgnd vpwr scs8hd_decap_12
XFILLER_43_86 vgnd vpwr scs8hd_decap_12
XFILLER_175_74 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_84_93 vgnd vpwr scs8hd_decap_12
XFILLER_83_3 vgnd vpwr scs8hd_decap_12
XFILLER_58_117 vgnd vpwr scs8hd_decap_8
XFILLER_104_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_102 vpwr vgnd scs8hd_fill_2
XFILLER_89_27 vgnd vpwr scs8hd_decap_12
XFILLER_161_98 vgnd vpwr scs8hd_decap_12
XFILLER_110_80 vgnd vpwr scs8hd_decap_12
XFILLER_117_111 vpwr vgnd scs8hd_fill_2
XFILLER_91_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_156_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_49_74 vgnd vpwr scs8hd_decap_12
XFILLER_65_51 vgnd vpwr scs8hd_decap_8
XFILLER_65_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_109 vgnd vpwr scs8hd_decap_12
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_101_27 vgnd vpwr scs8hd_decap_12
XFILLER_51_123 vpwr vgnd scs8hd_fill_2
XFILLER_126_68 vgnd vpwr scs8hd_decap_12
XFILLER_120_117 vgnd vpwr scs8hd_decap_8
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_142_56 vgnd vpwr scs8hd_decap_12
XFILLER_150_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_167_86 vgnd vpwr scs8hd_decap_12
XFILLER_51_86 vgnd vpwr scs8hd_decap_12
XFILLER_183_74 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
XFILLER_178_117 vgnd vpwr scs8hd_decap_8
XFILLER_92_93 vgnd vpwr scs8hd_decap_12
XFILLER_102_117 vgnd vpwr scs8hd_decap_8
XFILLER_112_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_80 vgnd vpwr scs8hd_fill_1
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XFILLER_169_106 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_129 vgnd vpwr scs8hd_decap_3
XFILLER_97_27 vgnd vpwr scs8hd_decap_12
XANTENNA__10__A _12_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XPHY_696 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_685 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_674 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_663 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_652 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_641 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_630 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_115 vgnd vpwr scs8hd_decap_8
XFILLER_107_59 vpwr vgnd scs8hd_fill_2
XFILLER_107_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XANTENNA__05__A _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_164_32 vgnd vpwr scs8hd_decap_12
XFILLER_148_44 vgnd vpwr scs8hd_decap_12
XFILLER_113_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_74 vgnd vpwr scs8hd_decap_12
XFILLER_189_62 vgnd vpwr scs8hd_decap_12
XFILLER_189_51 vgnd vpwr scs8hd_decap_8
XFILLER_73_51 vgnd vpwr scs8hd_decap_8
XFILLER_73_62 vgnd vpwr scs8hd_decap_12
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_171_123 vpwr vgnd scs8hd_fill_2
XFILLER_134_68 vgnd vpwr scs8hd_decap_12
XFILLER_150_56 vgnd vpwr scs8hd_decap_12
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XFILLER_159_98 vgnd vpwr scs8hd_decap_12
XFILLER_43_98 vgnd vpwr scs8hd_decap_12
XFILLER_175_86 vgnd vpwr scs8hd_decap_12
XFILLER_153_123 vpwr vgnd scs8hd_fill_2
XFILLER_108_80 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_191_63 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_decap_3
XFILLER_76_3 vgnd vpwr scs8hd_decap_12
XFILLER_104_27 vgnd vpwr scs8hd_decap_4
XFILLER_120_15 vgnd vpwr scs8hd_decap_12
XFILLER_81_110 vgnd vpwr scs8hd_decap_12
XFILLER_135_123 vpwr vgnd scs8hd_fill_2
XFILLER_89_39 vgnd vpwr scs8hd_decap_12
XFILLER_180_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XFILLER_117_123 vpwr vgnd scs8hd_fill_2
XFILLER_115_59 vpwr vgnd scs8hd_fill_2
XFILLER_115_15 vgnd vpwr scs8hd_decap_12
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_156_44 vgnd vpwr scs8hd_decap_12
XANTENNA__13__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_172_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XFILLER_65_74 vgnd vpwr scs8hd_decap_12
XFILLER_81_51 vgnd vpwr scs8hd_decap_8
XFILLER_81_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_101_39 vgnd vpwr scs8hd_decap_12
XFILLER_142_68 vgnd vpwr scs8hd_decap_12
XANTENNA__08__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_143_3 vgnd vpwr scs8hd_decap_12
XFILLER_167_98 vgnd vpwr scs8hd_decap_12
XFILLER_51_98 vgnd vpwr scs8hd_decap_12
XFILLER_183_86 vgnd vpwr scs8hd_decap_12
XFILLER_116_80 vgnd vpwr scs8hd_decap_12
XFILLER_112_27 vgnd vpwr scs8hd_decap_4
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XFILLER_24_124 vgnd vpwr scs8hd_fill_1
XPHY_108 vgnd vpwr scs8hd_decap_3
XPHY_119 vgnd vpwr scs8hd_decap_3
XFILLER_97_39 vgnd vpwr scs8hd_decap_12
XANTENNA__10__B enable vgnd vpwr scs8hd_diode_2
XPHY_620 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_102 vpwr vgnd scs8hd_fill_2
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XFILLER_183_110 vgnd vpwr scs8hd_decap_12
XPHY_697 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_686 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_675 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_664 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_653 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_642 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_631 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_123_15 vgnd vpwr scs8hd_decap_12
XFILLER_107_27 vgnd vpwr scs8hd_decap_12
XFILLER_88_105 vgnd vpwr scs8hd_decap_12
XFILLER_123_59 vpwr vgnd scs8hd_fill_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_165_110 vgnd vpwr scs8hd_decap_12
XFILLER_148_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XANTENNA__05__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_164_44 vgnd vpwr scs8hd_decap_12
XFILLER_106_3 vgnd vpwr scs8hd_decap_12
XANTENNA__21__A gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_diode_2
XFILLER_180_32 vgnd vpwr scs8hd_decap_12
XFILLER_57_86 vgnd vpwr scs8hd_decap_12
XFILLER_189_74 vgnd vpwr scs8hd_decap_12
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_73_74 vgnd vpwr scs8hd_decap_12
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_98_93 vgnd vpwr scs8hd_decap_12
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_147_110 vgnd vpwr scs8hd_decap_12
XFILLER_118_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_150_68 vgnd vpwr scs8hd_decap_12
XANTENNA__16__A gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_78 vpwr vgnd scs8hd_fill_2
XFILLER_175_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_191_75 vgnd vpwr scs8hd_decap_12
XFILLER_124_80 vgnd vpwr scs8hd_decap_12
XPHY_291 vgnd vpwr scs8hd_decap_3
XPHY_280 vgnd vpwr scs8hd_decap_3
XFILLER_129_110 vgnd vpwr scs8hd_decap_12
XFILLER_69_3 vgnd vpwr scs8hd_decap_12
XFILLER_120_27 vgnd vpwr scs8hd_decap_4
XFILLER_150_105 vgnd vpwr scs8hd_decap_12
XFILLER_173_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XFILLER_110_93 vgnd vpwr scs8hd_decap_12
XFILLER_79_51 vgnd vpwr scs8hd_decap_8
XFILLER_79_62 vgnd vpwr scs8hd_decap_12
XFILLER_132_105 vgnd vpwr scs8hd_decap_12
XFILLER_115_27 vgnd vpwr scs8hd_decap_12
XFILLER_131_15 vgnd vpwr scs8hd_decap_12
XFILLER_131_59 vpwr vgnd scs8hd_fill_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_6
XFILLER_156_56 vgnd vpwr scs8hd_decap_12
XANTENNA__13__B _13_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_172_44 vgnd vpwr scs8hd_decap_12
XFILLER_49_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_65_86 vgnd vpwr scs8hd_decap_12
XFILLER_81_74 vgnd vpwr scs8hd_decap_12
XFILLER_114_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_126_15 vgnd vpwr scs8hd_decap_12
XFILLER_136_3 vgnd vpwr scs8hd_decap_12
XFILLER_183_98 vgnd vpwr scs8hd_decap_12
XFILLER_132_80 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_14_ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_ebufn_1
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_93 vgnd vpwr scs8hd_decap_4
XPHY_109 vgnd vpwr scs8hd_decap_3
XANTENNA__10__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__19__A gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_diode_2
XPHY_643 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_632 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_621 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_610 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_178_32 vgnd vpwr scs8hd_decap_12
XPHY_698 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_687 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_676 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_665 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_654 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XFILLER_87_51 vgnd vpwr scs8hd_decap_8
XFILLER_87_62 vgnd vpwr scs8hd_decap_12
XFILLER_99_3 vgnd vpwr scs8hd_decap_12
XFILLER_107_39 vgnd vpwr scs8hd_decap_12
XFILLER_123_27 vgnd vpwr scs8hd_decap_12
XFILLER_88_117 vgnd vpwr scs8hd_decap_8
XFILLER_12_117 vgnd vpwr scs8hd_decap_8
XFILLER_148_68 vgnd vpwr scs8hd_decap_12
XANTENNA__05__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_164_56 vgnd vpwr scs8hd_decap_12
XFILLER_180_44 vgnd vpwr scs8hd_decap_12
XFILLER_57_98 vgnd vpwr scs8hd_decap_12
XFILLER_189_86 vgnd vpwr scs8hd_decap_12
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_73_86 vgnd vpwr scs8hd_decap_12
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_134_15 vgnd vpwr scs8hd_decap_12
XFILLER_118_27 vgnd vpwr scs8hd_decap_4
XFILLER_191_87 vgnd vpwr scs8hd_decap_6
XFILLER_191_32 vgnd vpwr scs8hd_decap_12
XFILLER_108_93 vgnd vpwr scs8hd_decap_12
XPHY_292 vgnd vpwr scs8hd_decap_3
XPHY_281 vgnd vpwr scs8hd_decap_3
XFILLER_140_80 vgnd vpwr scs8hd_decap_12
XPHY_270 vgnd vpwr scs8hd_decap_3
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_81_123 vpwr vgnd scs8hd_fill_2
XFILLER_129_59 vpwr vgnd scs8hd_fill_2
XFILLER_129_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_150_117 vgnd vpwr scs8hd_decap_8
XFILLER_166_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XFILLER_186_32 vgnd vpwr scs8hd_decap_12
XFILLER_70_32 vgnd vpwr scs8hd_decap_12
XFILLER_79_74 vgnd vpwr scs8hd_decap_12
XFILLER_95_62 vgnd vpwr scs8hd_decap_12
XFILLER_95_51 vgnd vpwr scs8hd_decap_8
XFILLER_63_123 vpwr vgnd scs8hd_fill_2
XFILLER_81_3 vgnd vpwr scs8hd_decap_12
XFILLER_132_117 vgnd vpwr scs8hd_decap_8
XFILLER_115_39 vgnd vpwr scs8hd_decap_12
XFILLER_131_27 vgnd vpwr scs8hd_decap_12
XFILLER_156_68 vgnd vpwr scs8hd_decap_12
XANTENNA__13__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_172_56 vgnd vpwr scs8hd_decap_12
XFILLER_45_123 vpwr vgnd scs8hd_fill_2
XFILLER_65_98 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_81_86 vgnd vpwr scs8hd_decap_12
XFILLER_114_117 vgnd vpwr scs8hd_decap_8
XFILLER_30_90 vpwr vgnd scs8hd_fill_2
XFILLER_126_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_142_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vpwr vgnd scs8hd_fill_2
XFILLER_129_3 vgnd vpwr scs8hd_decap_12
XFILLER_116_93 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _13_/Y vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_83 vgnd vpwr scs8hd_decap_8
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_137_59 vpwr vgnd scs8hd_fill_2
XFILLER_137_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XANTENNA__10__D _13_/D vgnd vpwr scs8hd_diode_2
XFILLER_46_56 vgnd vpwr scs8hd_decap_12
XFILLER_178_44 vgnd vpwr scs8hd_decap_12
XPHY_677 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_666 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_655 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_644 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_633 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_622 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_611 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_600 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _07_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_183_123 vpwr vgnd scs8hd_fill_2
XPHY_699 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_688 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_87_74 vgnd vpwr scs8hd_decap_12
XFILLER_123_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA__05__D enable vgnd vpwr scs8hd_diode_2
XFILLER_165_123 vpwr vgnd scs8hd_fill_2
XFILLER_164_68 vgnd vpwr scs8hd_decap_12
XFILLER_180_56 vgnd vpwr scs8hd_decap_12
XFILLER_189_98 vgnd vpwr scs8hd_decap_12
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_73_98 vgnd vpwr scs8hd_decap_12
XFILLER_138_80 vgnd vpwr scs8hd_decap_12
XFILLER_93_121 vgnd vpwr scs8hd_fill_1
XFILLER_147_123 vpwr vgnd scs8hd_fill_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_134_27 vgnd vpwr scs8hd_decap_4
XFILLER_150_15 vgnd vpwr scs8hd_decap_12
XFILLER_111_3 vgnd vpwr scs8hd_decap_12
XFILLER_191_44 vgnd vpwr scs8hd_decap_12
XFILLER_68_32 vgnd vpwr scs8hd_decap_12
XFILLER_75_110 vgnd vpwr scs8hd_decap_12
XFILLER_124_93 vgnd vpwr scs8hd_decap_12
XPHY_293 vgnd vpwr scs8hd_decap_3
XPHY_282 vgnd vpwr scs8hd_decap_3
XPHY_271 vgnd vpwr scs8hd_decap_3
XPHY_260 vgnd vpwr scs8hd_decap_3
XFILLER_129_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_145_15 vgnd vpwr scs8hd_decap_12
XFILLER_129_27 vgnd vpwr scs8hd_decap_12
XFILLER_1_106 vgnd vpwr scs8hd_decap_12
XFILLER_145_59 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_57_110 vgnd vpwr scs8hd_decap_12
XFILLER_159_3 vgnd vpwr scs8hd_decap_12
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
XFILLER_186_44 vgnd vpwr scs8hd_decap_12
XFILLER_70_44 vgnd vpwr scs8hd_decap_12
XFILLER_79_86 vgnd vpwr scs8hd_decap_12
XFILLER_95_74 vgnd vpwr scs8hd_decap_12
XFILLER_117_115 vgnd vpwr scs8hd_decap_6
XFILLER_74_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_131_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA__13__D _13_/D vgnd vpwr scs8hd_diode_2
XFILLER_172_68 vgnd vpwr scs8hd_decap_12
XFILLER_105_62 vgnd vpwr scs8hd_decap_12
XFILLER_105_51 vgnd vpwr scs8hd_decap_8
XFILLER_60_105 vgnd vpwr scs8hd_decap_12
XFILLER_81_98 vgnd vpwr scs8hd_decap_12
XFILLER_146_80 vgnd vpwr scs8hd_decap_12
XFILLER_142_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_76_32 vgnd vpwr scs8hd_decap_12
XFILLER_132_93 vgnd vpwr scs8hd_decap_12
XFILLER_25_80 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_decap_3
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_177_110 vgnd vpwr scs8hd_decap_12
XFILLER_137_27 vgnd vpwr scs8hd_decap_12
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XFILLER_153_15 vgnd vpwr scs8hd_decap_12
XFILLER_101_110 vgnd vpwr scs8hd_decap_12
XFILLER_153_59 vpwr vgnd scs8hd_fill_2
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XFILLER_178_56 vgnd vpwr scs8hd_decap_12
XPHY_689 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_678 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_141_3 vgnd vpwr scs8hd_decap_12
XPHY_667 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_656 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_645 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_634 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_623 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_612 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_601 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XFILLER_87_86 vgnd vpwr scs8hd_decap_12
XFILLER_159_110 vgnd vpwr scs8hd_decap_12
XFILLER_21_119 vgnd vpwr scs8hd_decap_3
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_180_105 vgnd vpwr scs8hd_decap_12
XFILLER_148_15 vgnd vpwr scs8hd_decap_12
XFILLER_189_3 vgnd vpwr scs8hd_decap_12
XFILLER_180_68 vgnd vpwr scs8hd_decap_12
XFILLER_113_62 vgnd vpwr scs8hd_decap_12
XFILLER_113_51 vgnd vpwr scs8hd_decap_8
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_154_80 vgnd vpwr scs8hd_decap_12
XFILLER_93_111 vpwr vgnd scs8hd_fill_2
XFILLER_162_105 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _14_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_150_27 vgnd vpwr scs8hd_decap_4
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_104_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_44 vgnd vpwr scs8hd_decap_12
XFILLER_191_56 vgnd vpwr scs8hd_decap_6
XFILLER_84_32 vgnd vpwr scs8hd_decap_12
XFILLER_140_93 vgnd vpwr scs8hd_decap_12
XPHY_261 vgnd vpwr scs8hd_decap_3
XPHY_250 vgnd vpwr scs8hd_decap_3
XPHY_294 vgnd vpwr scs8hd_decap_3
XFILLER_144_105 vgnd vpwr scs8hd_decap_4
XPHY_283 vgnd vpwr scs8hd_decap_3
XPHY_272 vgnd vpwr scs8hd_decap_3
XFILLER_129_39 vgnd vpwr scs8hd_decap_12
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_145_27 vgnd vpwr scs8hd_decap_12
XFILLER_1_118 vgnd vpwr scs8hd_decap_4
XFILLER_161_59 vpwr vgnd scs8hd_fill_2
XFILLER_161_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
XFILLER_186_56 vgnd vpwr scs8hd_decap_12
XFILLER_126_105 vgnd vpwr scs8hd_decap_12
XFILLER_70_56 vgnd vpwr scs8hd_decap_12
XFILLER_79_98 vgnd vpwr scs8hd_decap_12
XFILLER_95_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_80 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_67_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_156_15 vgnd vpwr scs8hd_decap_12
XFILLER_108_105 vgnd vpwr scs8hd_decap_12
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_171_3 vgnd vpwr scs8hd_decap_12
XFILLER_105_74 vgnd vpwr scs8hd_decap_12
XFILLER_45_114 vgnd vpwr scs8hd_decap_8
XFILLER_121_62 vgnd vpwr scs8hd_decap_12
XFILLER_121_51 vgnd vpwr scs8hd_decap_8
XFILLER_60_117 vgnd vpwr scs8hd_decap_8
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_162_80 vgnd vpwr scs8hd_decap_12
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_103 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_117 vgnd vpwr scs8hd_decap_8
XFILLER_76_44 vgnd vpwr scs8hd_decap_12
XFILLER_92_32 vgnd vpwr scs8hd_decap_12
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_decap_3
XFILLER_24_106 vgnd vpwr scs8hd_decap_12
XFILLER_137_39 vgnd vpwr scs8hd_decap_12
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XFILLER_153_27 vgnd vpwr scs8hd_decap_12
XPHY_602 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_106 vgnd vpwr scs8hd_decap_12
XFILLER_178_68 vgnd vpwr scs8hd_decap_12
XPHY_679 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_668 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_657 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_134_3 vgnd vpwr scs8hd_decap_12
XPHY_646 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_635 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_624 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_613 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
XFILLER_87_98 vgnd vpwr scs8hd_decap_12
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_148_27 vgnd vpwr scs8hd_decap_4
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_180_117 vgnd vpwr scs8hd_decap_8
XFILLER_164_15 vgnd vpwr scs8hd_decap_12
XFILLER_113_74 vgnd vpwr scs8hd_decap_12
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_138_93 vgnd vpwr scs8hd_decap_12
XFILLER_170_80 vgnd vpwr scs8hd_decap_12
XFILLER_93_123 vpwr vgnd scs8hd_fill_2
XFILLER_97_3 vgnd vpwr scs8hd_decap_12
XFILLER_162_117 vgnd vpwr scs8hd_decap_8
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_159_59 vpwr vgnd scs8hd_fill_2
XFILLER_159_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XFILLER_68_56 vgnd vpwr scs8hd_decap_12
XFILLER_75_123 vpwr vgnd scs8hd_fill_2
XFILLER_84_44 vgnd vpwr scs8hd_decap_12
XPHY_295 vgnd vpwr scs8hd_decap_3
XPHY_284 vgnd vpwr scs8hd_decap_3
XPHY_273 vgnd vpwr scs8hd_decap_3
XPHY_262 vgnd vpwr scs8hd_decap_3
XPHY_251 vgnd vpwr scs8hd_decap_3
XPHY_240 vgnd vpwr scs8hd_decap_3
XFILLER_144_117 vgnd vpwr scs8hd_decap_8
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_145_39 vgnd vpwr scs8hd_decap_12
XFILLER_161_27 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_123 vpwr vgnd scs8hd_fill_2
XFILLER_186_68 vgnd vpwr scs8hd_decap_12
XFILLER_126_117 vgnd vpwr scs8hd_decap_8
XFILLER_119_62 vgnd vpwr scs8hd_decap_12
XFILLER_119_51 vgnd vpwr scs8hd_decap_8
XFILLER_70_68 vgnd vpwr scs8hd_decap_12
XFILLER_95_98 vgnd vpwr scs8hd_decap_12
XFILLER_117_106 vgnd vpwr scs8hd_decap_3
XFILLER_44_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vpwr vgnd scs8hd_fill_2
XFILLER_156_27 vgnd vpwr scs8hd_decap_4
XFILLER_108_117 vgnd vpwr scs8hd_decap_8
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_172_15 vgnd vpwr scs8hd_decap_12
XFILLER_164_3 vgnd vpwr scs8hd_decap_12
XFILLER_105_86 vgnd vpwr scs8hd_decap_12
XFILLER_121_74 vgnd vpwr scs8hd_decap_12
XFILLER_146_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_82 vgnd vpwr scs8hd_decap_8
XFILLER_30_93 vgnd vpwr scs8hd_decap_6
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_167_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_167_59 vpwr vgnd scs8hd_fill_2
XFILLER_76_56 vgnd vpwr scs8hd_decap_12
XFILLER_92_44 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_2_97 vgnd vpwr scs8hd_fill_1
XFILLER_177_123 vpwr vgnd scs8hd_fill_2
XFILLER_24_118 vgnd vpwr scs8hd_decap_6
XFILLER_153_39 vgnd vpwr scs8hd_decap_12
XFILLER_101_123 vpwr vgnd scs8hd_fill_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
XPHY_625 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_614 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_603 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_32 vgnd vpwr scs8hd_decap_12
XFILLER_15_118 vgnd vpwr scs8hd_decap_4
XPHY_669 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_658 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_647 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_127_3 vgnd vpwr scs8hd_decap_12
XPHY_636 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_127_62 vgnd vpwr scs8hd_decap_12
XFILLER_127_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_159_123 vpwr vgnd scs8hd_fill_2
XFILLER_168_80 vgnd vpwr scs8hd_decap_12
XFILLER_52_80 vgnd vpwr scs8hd_decap_12
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_164_27 vgnd vpwr scs8hd_decap_4
XFILLER_87_110 vgnd vpwr scs8hd_decap_12
XFILLER_180_15 vgnd vpwr scs8hd_decap_12
XFILLER_113_86 vgnd vpwr scs8hd_decap_12
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_98_32 vgnd vpwr scs8hd_decap_12
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_154_93 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_0_ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_ebufn_1
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _07_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_159_27 vgnd vpwr scs8hd_decap_12
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XFILLER_175_59 vpwr vgnd scs8hd_fill_2
XFILLER_175_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_8
XFILLER_68_68 vgnd vpwr scs8hd_decap_12
XFILLER_90_105 vgnd vpwr scs8hd_decap_12
XFILLER_84_56 vgnd vpwr scs8hd_decap_12
XPHY_296 vgnd vpwr scs8hd_decap_3
XPHY_285 vgnd vpwr scs8hd_decap_3
XPHY_274 vgnd vpwr scs8hd_decap_3
XPHY_263 vgnd vpwr scs8hd_decap_3
XPHY_252 vgnd vpwr scs8hd_decap_3
XPHY_241 vgnd vpwr scs8hd_decap_3
XPHY_230 vgnd vpwr scs8hd_decap_3
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_161_39 vgnd vpwr scs8hd_decap_12
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_72_105 vgnd vpwr scs8hd_decap_12
XFILLER_110_32 vgnd vpwr scs8hd_decap_12
XFILLER_119_74 vgnd vpwr scs8hd_decap_12
XFILLER_135_62 vgnd vpwr scs8hd_decap_12
XFILLER_135_51 vgnd vpwr scs8hd_decap_8
XFILLER_28_93 vgnd vpwr scs8hd_decap_4
XFILLER_60_80 vgnd vpwr scs8hd_decap_12
XFILLER_176_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_54_105 vgnd vpwr scs8hd_decap_12
XFILLER_172_27 vgnd vpwr scs8hd_decap_4
XFILLER_131_110 vgnd vpwr scs8hd_decap_12
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XFILLER_157_3 vgnd vpwr scs8hd_decap_12
XFILLER_121_86 vgnd vpwr scs8hd_decap_12
XFILLER_105_98 vgnd vpwr scs8hd_decap_12
XFILLER_162_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XFILLER_189_110 vgnd vpwr scs8hd_decap_12
XFILLER_72_3 vgnd vpwr scs8hd_decap_12
XFILLER_113_110 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_167_27 vgnd vpwr scs8hd_decap_12
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XFILLER_183_59 vpwr vgnd scs8hd_fill_2
XFILLER_183_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XFILLER_76_68 vgnd vpwr scs8hd_decap_12
XFILLER_92_56 vgnd vpwr scs8hd_decap_12
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_decap_3
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_178_15 vgnd vpwr scs8hd_decap_12
XPHY_659 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_648 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_637 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_626 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_615 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_604 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_44 vgnd vpwr scs8hd_decap_12
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_127_74 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_143_62 vgnd vpwr scs8hd_decap_12
XFILLER_143_51 vgnd vpwr scs8hd_decap_8
XFILLER_174_105 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_184_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_180_27 vgnd vpwr scs8hd_decap_4
XFILLER_113_98 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XFILLER_156_105 vgnd vpwr scs8hd_decap_12
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_98_44 vgnd vpwr scs8hd_decap_12
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_170_93 vgnd vpwr scs8hd_decap_12
XFILLER_159_39 vgnd vpwr scs8hd_decap_12
XFILLER_138_105 vgnd vpwr scs8hd_decap_12
XFILLER_43_39 vgnd vpwr scs8hd_decap_12
XFILLER_175_27 vgnd vpwr scs8hd_decap_12
XFILLER_108_32 vgnd vpwr scs8hd_decap_12
XFILLER_191_15 vgnd vpwr scs8hd_decap_12
XFILLER_187_3 vgnd vpwr scs8hd_decap_12
XFILLER_90_117 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_84_68 vgnd vpwr scs8hd_decap_12
XPHY_297 vgnd vpwr scs8hd_decap_3
XPHY_286 vgnd vpwr scs8hd_decap_3
XPHY_275 vgnd vpwr scs8hd_decap_3
XPHY_264 vgnd vpwr scs8hd_decap_3
XPHY_253 vgnd vpwr scs8hd_decap_3
XPHY_242 vgnd vpwr scs8hd_decap_3
XPHY_231 vgnd vpwr scs8hd_decap_3
XPHY_220 vgnd vpwr scs8hd_decap_3
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XFILLER_72_117 vgnd vpwr scs8hd_decap_8
XFILLER_186_15 vgnd vpwr scs8hd_decap_12
XFILLER_110_44 vgnd vpwr scs8hd_decap_12
XFILLER_70_15 vgnd vpwr scs8hd_decap_12
XFILLER_119_86 vgnd vpwr scs8hd_decap_12
XFILLER_102_3 vgnd vpwr scs8hd_decap_12
XFILLER_151_51 vgnd vpwr scs8hd_decap_8
XFILLER_135_74 vgnd vpwr scs8hd_decap_12
XFILLER_151_62 vgnd vpwr scs8hd_decap_12
XFILLER_44_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_54_117 vgnd vpwr scs8hd_decap_8
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XFILLER_65_15 vgnd vpwr scs8hd_decap_12
XFILLER_121_98 vgnd vpwr scs8hd_decap_12
XFILLER_65_59 vpwr vgnd scs8hd_fill_2
XFILLER_36_117 vgnd vpwr scs8hd_decap_8
XFILLER_65_3 vgnd vpwr scs8hd_decap_12
XFILLER_167_39 vgnd vpwr scs8hd_decap_12
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
XFILLER_183_27 vgnd vpwr scs8hd_decap_12
XFILLER_116_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_117 vgnd vpwr scs8hd_decap_8
XFILLER_92_68 vgnd vpwr scs8hd_decap_12
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_decap_3
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_66_80 vgnd vpwr scs8hd_decap_12
XFILLER_178_27 vgnd vpwr scs8hd_decap_4
XPHY_649 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_638 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_627 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_616 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_605 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_56 vgnd vpwr scs8hd_decap_12
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XFILLER_127_86 vgnd vpwr scs8hd_decap_12
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XFILLER_143_74 vgnd vpwr scs8hd_decap_12
XFILLER_174_117 vgnd vpwr scs8hd_decap_8
XFILLER_168_93 vgnd vpwr scs8hd_decap_12
XFILLER_52_93 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XFILLER_87_123 vpwr vgnd scs8hd_fill_2
XFILLER_189_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_59 vpwr vgnd scs8hd_fill_2
XFILLER_189_59 vpwr vgnd scs8hd_fill_2
XFILLER_156_117 vgnd vpwr scs8hd_decap_8
XFILLER_132_3 vgnd vpwr scs8hd_decap_12
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_98_56 vgnd vpwr scs8hd_decap_12
XFILLER_22_74 vgnd vpwr scs8hd_fill_1
XFILLER_93_115 vgnd vpwr scs8hd_decap_6
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_69_123 vpwr vgnd scs8hd_fill_2
X_19_ gfpga_pad_GPIO_PAD[0] right_width_0_height_0__pin_1_ vgnd vpwr scs8hd_buf_2
XFILLER_138_117 vgnd vpwr scs8hd_decap_8
XFILLER_175_39 vgnd vpwr scs8hd_decap_12
XFILLER_108_44 vgnd vpwr scs8hd_decap_12
XFILLER_68_15 vgnd vpwr scs8hd_decap_12
XFILLER_191_27 vgnd vpwr scs8hd_decap_4
XFILLER_124_32 vgnd vpwr scs8hd_decap_12
XPHY_243 vgnd vpwr scs8hd_decap_3
XPHY_232 vgnd vpwr scs8hd_decap_3
XPHY_221 vgnd vpwr scs8hd_decap_3
XPHY_210 vgnd vpwr scs8hd_decap_3
XFILLER_17_74 vgnd vpwr scs8hd_decap_3
XFILLER_149_62 vgnd vpwr scs8hd_decap_12
XFILLER_149_51 vgnd vpwr scs8hd_decap_8
XPHY_298 vgnd vpwr scs8hd_decap_3
XPHY_287 vgnd vpwr scs8hd_decap_3
XPHY_276 vgnd vpwr scs8hd_decap_3
XPHY_265 vgnd vpwr scs8hd_decap_3
XPHY_254 vgnd vpwr scs8hd_decap_3
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_95_3 vgnd vpwr scs8hd_decap_12
XFILLER_74_80 vgnd vpwr scs8hd_decap_12
XFILLER_186_27 vgnd vpwr scs8hd_decap_4
XFILLER_110_56 vgnd vpwr scs8hd_decap_12
XFILLER_70_27 vgnd vpwr scs8hd_decap_4
XFILLER_119_98 vgnd vpwr scs8hd_decap_12
XFILLER_151_74 vgnd vpwr scs8hd_decap_12
XFILLER_135_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XFILLER_176_93 vgnd vpwr scs8hd_decap_12
XFILLER_60_93 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_131_123 vpwr vgnd scs8hd_fill_2
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
XFILLER_65_27 vgnd vpwr scs8hd_decap_12
XFILLER_81_15 vgnd vpwr scs8hd_decap_12
XFILLER_81_59 vpwr vgnd scs8hd_fill_2
XFILLER_189_123 vpwr vgnd scs8hd_fill_2
XFILLER_113_123 vpwr vgnd scs8hd_fill_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_27_107 vgnd vpwr scs8hd_decap_3
XFILLER_27_118 vgnd vpwr scs8hd_decap_4
XFILLER_183_39 vgnd vpwr scs8hd_decap_12
XFILLER_116_44 vgnd vpwr scs8hd_decap_12
XFILLER_76_15 vgnd vpwr scs8hd_decap_12
XFILLER_162_3 vgnd vpwr scs8hd_decap_12
XFILLER_132_32 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XFILLER_157_62 vgnd vpwr scs8hd_decap_12
XFILLER_157_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_82_80 vgnd vpwr scs8hd_decap_12
XFILLER_99_110 vgnd vpwr scs8hd_decap_12
XPHY_639 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_628 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_617 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_606 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_121 vgnd vpwr scs8hd_fill_1
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_143_86 vgnd vpwr scs8hd_decap_12
XFILLER_127_98 vgnd vpwr scs8hd_decap_12
XFILLER_184_93 vgnd vpwr scs8hd_decap_12
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
XFILLER_189_27 vgnd vpwr scs8hd_decap_12
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_73_27 vgnd vpwr scs8hd_decap_12
XFILLER_125_3 vgnd vpwr scs8hd_decap_12
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_98_68 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_84_105 vgnd vpwr scs8hd_decap_12
X_18_ gfpga_pad_GPIO_PAD[7] right_width_0_height_0__pin_15_ vgnd vpwr scs8hd_buf_2
XFILLER_161_110 vgnd vpwr scs8hd_decap_12
XFILLER_108_56 vgnd vpwr scs8hd_decap_12
XFILLER_68_27 vgnd vpwr scs8hd_decap_4
XFILLER_124_44 vgnd vpwr scs8hd_decap_12
XFILLER_84_15 vgnd vpwr scs8hd_decap_12
XFILLER_140_32 vgnd vpwr scs8hd_decap_12
XPHY_277 vgnd vpwr scs8hd_decap_3
XPHY_266 vgnd vpwr scs8hd_decap_3
XPHY_255 vgnd vpwr scs8hd_decap_3
XPHY_244 vgnd vpwr scs8hd_decap_3
XPHY_233 vgnd vpwr scs8hd_decap_3
XPHY_222 vgnd vpwr scs8hd_decap_3
XPHY_211 vgnd vpwr scs8hd_decap_3
XPHY_200 vgnd vpwr scs8hd_decap_3
XPHY_299 vgnd vpwr scs8hd_decap_3
XFILLER_149_74 vgnd vpwr scs8hd_decap_12
XPHY_288 vgnd vpwr scs8hd_decap_3
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_165_62 vgnd vpwr scs8hd_decap_12
XFILLER_165_51 vgnd vpwr scs8hd_decap_8
XFILLER_66_105 vgnd vpwr scs8hd_decap_12
XFILLER_58_93 vgnd vpwr scs8hd_decap_12
XFILLER_90_80 vgnd vpwr scs8hd_decap_12
XFILLER_88_3 vgnd vpwr scs8hd_decap_12
XFILLER_143_121 vgnd vpwr scs8hd_fill_1
XFILLER_110_68 vgnd vpwr scs8hd_decap_12
XFILLER_79_15 vgnd vpwr scs8hd_decap_12
XFILLER_135_98 vgnd vpwr scs8hd_decap_12
XFILLER_48_105 vgnd vpwr scs8hd_decap_12
XFILLER_79_59 vpwr vgnd scs8hd_fill_2
XFILLER_151_86 vgnd vpwr scs8hd_decap_12
XFILLER_125_110 vgnd vpwr scs8hd_decap_12
XFILLER_65_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_81_27 vgnd vpwr scs8hd_decap_12
XFILLER_107_110 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_116_56 vgnd vpwr scs8hd_decap_12
XFILLER_76_27 vgnd vpwr scs8hd_decap_4
XFILLER_155_3 vgnd vpwr scs8hd_decap_12
XFILLER_132_44 vgnd vpwr scs8hd_decap_12
XFILLER_92_15 vgnd vpwr scs8hd_decap_12
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XFILLER_186_105 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_86 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XFILLER_173_62 vgnd vpwr scs8hd_decap_12
XFILLER_173_51 vgnd vpwr scs8hd_decap_8
XFILLER_157_74 vgnd vpwr scs8hd_decap_12
XFILLER_110_105 vgnd vpwr scs8hd_decap_12
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_66_93 vgnd vpwr scs8hd_decap_12
XFILLER_70_3 vgnd vpwr scs8hd_decap_12
XPHY_607 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_111 vpwr vgnd scs8hd_fill_2
XFILLER_168_105 vgnd vpwr scs8hd_decap_12
XPHY_629 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_618 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_87_15 vgnd vpwr scs8hd_decap_12
XFILLER_87_59 vpwr vgnd scs8hd_fill_2
XFILLER_143_98 vgnd vpwr scs8hd_decap_8
XFILLER_189_39 vgnd vpwr scs8hd_decap_12
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_73_39 vgnd vpwr scs8hd_decap_12
XFILLER_138_32 vgnd vpwr scs8hd_decap_12
XFILLER_118_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_93_106 vgnd vpwr scs8hd_decap_3
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_114 vgnd vpwr scs8hd_decap_8
XFILLER_84_117 vgnd vpwr scs8hd_decap_8
XFILLER_88_80 vgnd vpwr scs8hd_decap_12
X_17_ gfpga_pad_GPIO_PAD[6] right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_buf_2
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_108_68 vgnd vpwr scs8hd_decap_12
XFILLER_124_56 vgnd vpwr scs8hd_decap_12
XFILLER_84_27 vgnd vpwr scs8hd_decap_4
XPHY_289 vgnd vpwr scs8hd_decap_3
XFILLER_140_44 vgnd vpwr scs8hd_decap_12
XPHY_278 vgnd vpwr scs8hd_decap_3
XPHY_267 vgnd vpwr scs8hd_decap_3
XPHY_256 vgnd vpwr scs8hd_decap_3
XPHY_245 vgnd vpwr scs8hd_decap_3
XPHY_234 vgnd vpwr scs8hd_decap_3
XPHY_223 vgnd vpwr scs8hd_decap_3
XPHY_212 vgnd vpwr scs8hd_decap_3
XPHY_201 vgnd vpwr scs8hd_decap_3
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_149_86 vgnd vpwr scs8hd_decap_12
XFILLER_181_62 vgnd vpwr scs8hd_decap_12
XFILLER_181_51 vgnd vpwr scs8hd_decap_8
XFILLER_165_74 vgnd vpwr scs8hd_decap_12
XFILLER_66_117 vgnd vpwr scs8hd_decap_8
XFILLER_74_93 vgnd vpwr scs8hd_decap_12
XFILLER_143_111 vpwr vgnd scs8hd_fill_2
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _09_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_79_27 vgnd vpwr scs8hd_decap_12
XFILLER_95_59 vpwr vgnd scs8hd_fill_2
XFILLER_95_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_117 vgnd vpwr scs8hd_decap_8
XFILLER_185_3 vgnd vpwr scs8hd_decap_12
XFILLER_151_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_97 vgnd vpwr scs8hd_fill_1
XFILLER_100_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_81_39 vgnd vpwr scs8hd_decap_12
XFILLER_146_32 vgnd vpwr scs8hd_decap_12
XFILLER_100_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_44_120 vgnd vpwr scs8hd_decap_4
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_96_80 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_2_ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_ebufn_1
XFILLER_116_68 vgnd vpwr scs8hd_decap_12
XFILLER_186_117 vgnd vpwr scs8hd_decap_8
XFILLER_148_3 vgnd vpwr scs8hd_decap_12
XFILLER_132_56 vgnd vpwr scs8hd_decap_12
XFILLER_92_27 vgnd vpwr scs8hd_decap_4
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_76 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vpwr vgnd scs8hd_fill_2
XPHY_87 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XFILLER_173_74 vgnd vpwr scs8hd_decap_12
XFILLER_157_86 vgnd vpwr scs8hd_decap_12
XFILLER_110_117 vgnd vpwr scs8hd_decap_8
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XFILLER_82_93 vgnd vpwr scs8hd_decap_12
XFILLER_99_123 vpwr vgnd scs8hd_fill_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_168_117 vgnd vpwr scs8hd_decap_8
XPHY_619 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_608 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_87_27 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _14_/Y vgnd vpwr scs8hd_diode_2
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_138_44 vgnd vpwr scs8hd_decap_12
XFILLER_98_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_154_32 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XFILLER_47_74 vgnd vpwr scs8hd_decap_12
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_179_62 vgnd vpwr scs8hd_decap_12
XFILLER_179_51 vgnd vpwr scs8hd_decap_8
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
X_16_ gfpga_pad_GPIO_PAD[5] right_width_0_height_0__pin_11_ vgnd vpwr scs8hd_buf_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_161_123 vpwr vgnd scs8hd_fill_2
XFILLER_140_56 vgnd vpwr scs8hd_decap_12
XFILLER_124_68 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_decap_3
XPHY_268 vgnd vpwr scs8hd_decap_3
XFILLER_130_3 vgnd vpwr scs8hd_decap_12
XPHY_257 vgnd vpwr scs8hd_decap_3
XPHY_246 vgnd vpwr scs8hd_decap_3
XPHY_235 vgnd vpwr scs8hd_decap_3
XPHY_224 vgnd vpwr scs8hd_decap_3
XPHY_213 vgnd vpwr scs8hd_decap_3
XPHY_202 vgnd vpwr scs8hd_decap_3
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_165_86 vgnd vpwr scs8hd_decap_12
XFILLER_149_98 vgnd vpwr scs8hd_decap_12
XFILLER_181_74 vgnd vpwr scs8hd_decap_12
XFILLER_143_123 vpwr vgnd scs8hd_fill_2
XFILLER_90_93 vgnd vpwr scs8hd_decap_12
XFILLER_110_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_91 vpwr vgnd scs8hd_fill_2
XFILLER_79_39 vgnd vpwr scs8hd_decap_12
XFILLER_95_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_178_3 vgnd vpwr scs8hd_decap_12
XFILLER_71_110 vgnd vpwr scs8hd_decap_12
XFILLER_125_123 vpwr vgnd scs8hd_fill_2
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_93_3 vgnd vpwr scs8hd_decap_12
XFILLER_105_59 vpwr vgnd scs8hd_fill_2
XFILLER_105_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_146_44 vgnd vpwr scs8hd_decap_12
XFILLER_107_123 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_99 vgnd vpwr scs8hd_fill_1
XFILLER_162_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_55_74 vgnd vpwr scs8hd_decap_12
XFILLER_71_51 vgnd vpwr scs8hd_decap_8
XFILLER_71_62 vgnd vpwr scs8hd_decap_12
XFILLER_187_62 vgnd vpwr scs8hd_decap_12
XFILLER_187_51 vgnd vpwr scs8hd_decap_8
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _15_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_132_68 vgnd vpwr scs8hd_decap_12
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_decap_3
XFILLER_157_98 vgnd vpwr scs8hd_decap_12
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_173_86 vgnd vpwr scs8hd_decap_12
XFILLER_106_80 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
XPHY_609 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_102_27 vgnd vpwr scs8hd_decap_4
XFILLER_87_39 vgnd vpwr scs8hd_decap_12
XFILLER_160_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_96_105 vgnd vpwr scs8hd_decap_12
XFILLER_20_105 vgnd vpwr scs8hd_decap_4
XFILLER_173_110 vgnd vpwr scs8hd_decap_12
XFILLER_113_59 vpwr vgnd scs8hd_fill_2
XFILLER_113_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_138_56 vgnd vpwr scs8hd_decap_12
XFILLER_98_27 vgnd vpwr scs8hd_decap_4
XANTENNA__11__A enable vgnd vpwr scs8hd_diode_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XFILLER_170_32 vgnd vpwr scs8hd_decap_12
XFILLER_154_44 vgnd vpwr scs8hd_decap_12
XFILLER_78_105 vgnd vpwr scs8hd_decap_8
XFILLER_47_86 vgnd vpwr scs8hd_decap_12
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_179_74 vgnd vpwr scs8hd_decap_12
XFILLER_155_110 vgnd vpwr scs8hd_decap_12
XFILLER_88_93 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
X_15_ address[1] _13_/B _13_/C address[2] _15_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_108_15 vgnd vpwr scs8hd_decap_12
XFILLER_140_68 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_decap_3
XPHY_214 vgnd vpwr scs8hd_decap_3
XPHY_203 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
XFILLER_137_110 vgnd vpwr scs8hd_decap_12
XPHY_269 vgnd vpwr scs8hd_decap_3
XPHY_258 vgnd vpwr scs8hd_decap_3
XPHY_247 vgnd vpwr scs8hd_decap_3
XFILLER_123_3 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_decap_3
XANTENNA__06__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_165_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_123 vpwr vgnd scs8hd_fill_2
XFILLER_181_86 vgnd vpwr scs8hd_decap_12
XFILLER_114_80 vgnd vpwr scs8hd_decap_12
XPHY_770 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_119_110 vgnd vpwr scs8hd_decap_12
XFILLER_110_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_104 vpwr vgnd scs8hd_fill_2
XFILLER_95_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_44_32 vgnd vpwr scs8hd_decap_12
XFILLER_100_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_140_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_69_51 vgnd vpwr scs8hd_decap_8
XFILLER_69_62 vgnd vpwr scs8hd_decap_12
XFILLER_86_3 vgnd vpwr scs8hd_decap_12
XFILLER_105_27 vgnd vpwr scs8hd_decap_12
XFILLER_121_59 vpwr vgnd scs8hd_fill_2
XFILLER_121_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_162_44 vgnd vpwr scs8hd_decap_12
XFILLER_146_56 vgnd vpwr scs8hd_decap_12
XFILLER_122_105 vgnd vpwr scs8hd_decap_12
XFILLER_190_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_55_86 vgnd vpwr scs8hd_decap_12
XFILLER_187_74 vgnd vpwr scs8hd_decap_12
XFILLER_71_74 vgnd vpwr scs8hd_decap_12
XFILLER_96_93 vgnd vpwr scs8hd_decap_12
XFILLER_116_15 vgnd vpwr scs8hd_decap_12
XFILLER_104_105 vgnd vpwr scs8hd_decap_12
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XANTENNA__14__A _12_/A vgnd vpwr scs8hd_diode_2
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_173_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_122_80 vgnd vpwr scs8hd_decap_12
XFILLER_17_100 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XFILLER_153_3 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_168_32 vgnd vpwr scs8hd_decap_12
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
XFILLER_96_117 vgnd vpwr scs8hd_decap_8
XFILLER_77_51 vgnd vpwr scs8hd_decap_8
XFILLER_77_62 vgnd vpwr scs8hd_decap_12
XFILLER_20_117 vgnd vpwr scs8hd_decap_8
XFILLER_113_27 vgnd vpwr scs8hd_decap_12
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_138_68 vgnd vpwr scs8hd_decap_12
XFILLER_22_68 vgnd vpwr scs8hd_decap_6
XFILLER_78_117 vgnd vpwr scs8hd_decap_8
XFILLER_170_44 vgnd vpwr scs8hd_decap_12
XFILLER_154_56 vgnd vpwr scs8hd_decap_12
XFILLER_47_98 vgnd vpwr scs8hd_decap_12
XFILLER_179_86 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
X_14_ _12_/A _13_/B _13_/C address[2] _14_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_108_27 vgnd vpwr scs8hd_decap_4
XFILLER_124_15 vgnd vpwr scs8hd_decap_12
XPHY_259 vgnd vpwr scs8hd_decap_3
XPHY_248 vgnd vpwr scs8hd_decap_3
XPHY_237 vgnd vpwr scs8hd_decap_3
XPHY_226 vgnd vpwr scs8hd_decap_3
XPHY_215 vgnd vpwr scs8hd_decap_3
XPHY_204 vgnd vpwr scs8hd_decap_3
XFILLER_17_79 vpwr vgnd scs8hd_fill_2
XFILLER_116_3 vgnd vpwr scs8hd_decap_12
XANTENNA__22__A gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_diode_2
XFILLER_181_98 vgnd vpwr scs8hd_decap_12
XPHY_771 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_760 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_80 vgnd vpwr scs8hd_decap_12
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_119_59 vpwr vgnd scs8hd_fill_2
XFILLER_119_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_116 vgnd vpwr scs8hd_decap_8
XANTENNA__17__A gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_71_123 vpwr vgnd scs8hd_fill_2
XFILLER_44_44 vgnd vpwr scs8hd_decap_12
XFILLER_176_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_140_117 vgnd vpwr scs8hd_decap_8
XFILLER_69_74 vgnd vpwr scs8hd_decap_12
XFILLER_85_51 vgnd vpwr scs8hd_decap_8
XFILLER_85_62 vgnd vpwr scs8hd_decap_12
XPHY_590 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_79_3 vgnd vpwr scs8hd_decap_12
XFILLER_105_39 vgnd vpwr scs8hd_decap_12
XFILLER_53_123 vpwr vgnd scs8hd_fill_2
XFILLER_121_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_162_56 vgnd vpwr scs8hd_decap_12
XFILLER_146_68 vgnd vpwr scs8hd_decap_12
XFILLER_122_117 vgnd vpwr scs8hd_decap_8
XFILLER_183_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_98 vgnd vpwr scs8hd_decap_12
XFILLER_187_86 vgnd vpwr scs8hd_decap_12
XFILLER_71_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vpwr vgnd scs8hd_fill_2
XFILLER_116_27 vgnd vpwr scs8hd_decap_4
XFILLER_104_117 vgnd vpwr scs8hd_decap_8
XFILLER_132_15 vgnd vpwr scs8hd_decap_12
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_26_101 vgnd vpwr scs8hd_decap_3
XFILLER_26_123 vpwr vgnd scs8hd_fill_2
XANTENNA__14__B _13_/B vgnd vpwr scs8hd_diode_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_106_93 vgnd vpwr scs8hd_decap_12
XFILLER_17_112 vgnd vpwr scs8hd_decap_8
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_115 vgnd vpwr scs8hd_decap_6
XFILLER_127_59 vpwr vgnd scs8hd_fill_2
XFILLER_127_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XANTENNA__09__B enable vgnd vpwr scs8hd_diode_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_168_44 vgnd vpwr scs8hd_decap_12
XFILLER_146_3 vgnd vpwr scs8hd_decap_12
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XFILLER_184_32 vgnd vpwr scs8hd_decap_12
XFILLER_93_62 vgnd vpwr scs8hd_decap_12
XFILLER_93_51 vgnd vpwr scs8hd_decap_8
XFILLER_77_74 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_173_123 vpwr vgnd scs8hd_fill_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XFILLER_113_39 vgnd vpwr scs8hd_decap_12
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_154_68 vgnd vpwr scs8hd_decap_12
XFILLER_170_56 vgnd vpwr scs8hd_decap_12
XFILLER_179_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_155_123 vpwr vgnd scs8hd_fill_2
XFILLER_128_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
X_13_ address[1] _13_/B _13_/C _13_/D _13_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_140_15 vgnd vpwr scs8hd_decap_12
XFILLER_124_27 vgnd vpwr scs8hd_decap_4
XFILLER_83_110 vgnd vpwr scs8hd_decap_12
XPHY_249 vgnd vpwr scs8hd_decap_3
XPHY_238 vgnd vpwr scs8hd_decap_3
XPHY_227 vgnd vpwr scs8hd_decap_3
XPHY_216 vgnd vpwr scs8hd_decap_3
XPHY_205 vgnd vpwr scs8hd_decap_3
XFILLER_137_123 vpwr vgnd scs8hd_fill_2
XFILLER_109_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
XFILLER_114_93 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _09_/X vgnd vpwr scs8hd_diode_2
XPHY_761 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_750 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_143_115 vgnd vpwr scs8hd_decap_6
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_65_110 vgnd vpwr scs8hd_decap_12
XFILLER_0_83 vgnd vpwr scs8hd_decap_8
XFILLER_0_94 vgnd vpwr scs8hd_decap_8
XFILLER_119_123 vpwr vgnd scs8hd_fill_2
XFILLER_119_27 vgnd vpwr scs8hd_decap_12
XFILLER_135_59 vpwr vgnd scs8hd_fill_2
XFILLER_135_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_44_56 vgnd vpwr scs8hd_decap_12
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XFILLER_176_44 vgnd vpwr scs8hd_decap_12
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_47_110 vgnd vpwr scs8hd_decap_12
XFILLER_69_86 vgnd vpwr scs8hd_decap_12
XFILLER_85_74 vgnd vpwr scs8hd_decap_12
XPHY_591 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_580 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_121_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_162_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_110 vpwr vgnd scs8hd_fill_2
XFILLER_176_3 vgnd vpwr scs8hd_decap_12
XFILLER_44_124 vgnd vpwr scs8hd_fill_1
XFILLER_187_98 vgnd vpwr scs8hd_decap_12
XFILLER_71_98 vgnd vpwr scs8hd_decap_12
XFILLER_136_80 vgnd vpwr scs8hd_decap_12
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XFILLER_91_3 vgnd vpwr scs8hd_decap_12
XFILLER_50_105 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XFILLER_132_27 vgnd vpwr scs8hd_decap_4
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XANTENNA__14__C _13_/C vgnd vpwr scs8hd_diode_2
XFILLER_66_32 vgnd vpwr scs8hd_decap_12
XFILLER_185_110 vgnd vpwr scs8hd_decap_12
XFILLER_122_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_127_27 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XFILLER_143_59 vpwr vgnd scs8hd_fill_2
XFILLER_143_15 vgnd vpwr scs8hd_decap_12
XANTENNA__09__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_167_110 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XFILLER_184_44 vgnd vpwr scs8hd_decap_12
XFILLER_168_56 vgnd vpwr scs8hd_decap_12
XFILLER_139_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_86 vgnd vpwr scs8hd_decap_12
XFILLER_93_74 vgnd vpwr scs8hd_decap_12
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XFILLER_149_110 vgnd vpwr scs8hd_decap_12
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_138_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_170_68 vgnd vpwr scs8hd_decap_12
XFILLER_103_62 vgnd vpwr scs8hd_decap_12
XFILLER_103_51 vgnd vpwr scs8hd_decap_8
XFILLER_170_105 vgnd vpwr scs8hd_decap_4
XFILLER_144_80 vgnd vpwr scs8hd_decap_12
X_12_ _12_/A _13_/B _13_/C _13_/D _12_/Y vgnd vpwr scs8hd_nor4_4
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_4_ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_ebufn_1
XFILLER_140_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XPHY_239 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_decap_3
XPHY_217 vgnd vpwr scs8hd_decap_3
XPHY_206 vgnd vpwr scs8hd_decap_3
XFILLER_152_105 vgnd vpwr scs8hd_decap_8
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
XFILLER_74_32 vgnd vpwr scs8hd_decap_12
XPHY_762 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_751 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_740 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_93 vgnd vpwr scs8hd_decap_12
XFILLER_99_62 vgnd vpwr scs8hd_decap_12
XFILLER_99_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_134_105 vgnd vpwr scs8hd_decap_12
XFILLER_119_39 vgnd vpwr scs8hd_decap_12
XFILLER_151_15 vgnd vpwr scs8hd_decap_12
XFILLER_135_27 vgnd vpwr scs8hd_decap_12
XFILLER_151_59 vpwr vgnd scs8hd_fill_2
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_176_56 vgnd vpwr scs8hd_decap_12
XFILLER_121_3 vgnd vpwr scs8hd_decap_12
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XFILLER_69_98 vgnd vpwr scs8hd_decap_6
XFILLER_18_80 vgnd vpwr scs8hd_decap_3
XFILLER_85_86 vgnd vpwr scs8hd_decap_12
XPHY_570 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_116_105 vgnd vpwr scs8hd_decap_12
XPHY_592 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_581 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_53_114 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_146_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_169_3 vgnd vpwr scs8hd_decap_12
XFILLER_111_62 vgnd vpwr scs8hd_decap_12
XFILLER_111_51 vgnd vpwr scs8hd_decap_8
XFILLER_152_80 vgnd vpwr scs8hd_decap_12
XFILLER_50_117 vgnd vpwr scs8hd_decap_8
XFILLER_84_3 vgnd vpwr scs8hd_decap_12
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA__14__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_66_44 vgnd vpwr scs8hd_decap_12
XFILLER_82_32 vgnd vpwr scs8hd_decap_12
XFILLER_32_117 vgnd vpwr scs8hd_decap_8
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_143_27 vgnd vpwr scs8hd_decap_12
XFILLER_127_39 vgnd vpwr scs8hd_decap_12
XANTENNA__09__D _13_/D vgnd vpwr scs8hd_diode_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_8
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
XFILLER_184_56 vgnd vpwr scs8hd_decap_12
XFILLER_168_68 vgnd vpwr scs8hd_decap_12
XFILLER_77_98 vgnd vpwr scs8hd_decap_12
XFILLER_93_86 vgnd vpwr scs8hd_decap_12
XFILLER_26_80 vpwr vgnd scs8hd_fill_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_95 vgnd vpwr scs8hd_decap_12
XFILLER_138_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_154_15 vgnd vpwr scs8hd_decap_12
XFILLER_151_3 vgnd vpwr scs8hd_decap_12
XFILLER_103_74 vgnd vpwr scs8hd_decap_12
XFILLER_170_117 vgnd vpwr scs8hd_decap_8
XFILLER_128_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
X_11_ enable _13_/B vgnd vpwr scs8hd_inv_8
XFILLER_160_80 vgnd vpwr scs8hd_decap_12
XFILLER_68_120 vgnd vpwr scs8hd_decap_4
XPHY_207 vgnd vpwr scs8hd_decap_3
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_83_123 vpwr vgnd scs8hd_fill_2
XFILLER_149_59 vpwr vgnd scs8hd_fill_2
XFILLER_149_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_decap_3
XPHY_218 vgnd vpwr scs8hd_decap_3
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_152_117 vgnd vpwr scs8hd_decap_8
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
XPHY_763 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_752 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_741 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_730 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_90_32 vgnd vpwr scs8hd_decap_12
XFILLER_74_44 vgnd vpwr scs8hd_decap_12
XFILLER_143_106 vgnd vpwr scs8hd_decap_3
XFILLER_99_74 vgnd vpwr scs8hd_decap_12
XFILLER_23_81 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_65_123 vpwr vgnd scs8hd_fill_2
XFILLER_134_117 vgnd vpwr scs8hd_decap_8
XFILLER_151_27 vgnd vpwr scs8hd_decap_12
XFILLER_135_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_176_68 vgnd vpwr scs8hd_decap_12
XFILLER_114_3 vgnd vpwr scs8hd_decap_12
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XFILLER_109_62 vgnd vpwr scs8hd_decap_12
XFILLER_109_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_123 vpwr vgnd scs8hd_fill_2
XFILLER_85_98 vgnd vpwr scs8hd_decap_12
XPHY_593 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_582 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_571 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_116_117 vgnd vpwr scs8hd_decap_8
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_162_15 vgnd vpwr scs8hd_decap_12
XFILLER_146_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_123 vpwr vgnd scs8hd_fill_2
XFILLER_111_74 vgnd vpwr scs8hd_decap_12
XFILLER_136_93 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XFILLER_29_91 vpwr vgnd scs8hd_fill_2
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_77_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_115 vgnd vpwr scs8hd_decap_8
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XFILLER_157_59 vpwr vgnd scs8hd_fill_2
XFILLER_157_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_181_3 vgnd vpwr scs8hd_decap_12
XFILLER_66_56 vgnd vpwr scs8hd_decap_12
XFILLER_82_44 vgnd vpwr scs8hd_decap_12
XFILLER_185_123 vpwr vgnd scs8hd_fill_2
XFILLER_143_39 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_167_123 vpwr vgnd scs8hd_fill_2
XFILLER_184_68 vgnd vpwr scs8hd_decap_12
XFILLER_117_62 vgnd vpwr scs8hd_decap_12
XFILLER_117_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_93_98 vgnd vpwr scs8hd_decap_8
XFILLER_158_80 vgnd vpwr scs8hd_decap_12
XFILLER_42_80 vgnd vpwr scs8hd_decap_12
XFILLER_95_110 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_149_123 vpwr vgnd scs8hd_fill_2
XFILLER_154_27 vgnd vpwr scs8hd_decap_4
XFILLER_170_15 vgnd vpwr scs8hd_decap_12
XFILLER_103_86 vgnd vpwr scs8hd_decap_12
XFILLER_144_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_110 vgnd vpwr scs8hd_decap_3
XFILLER_77_121 vgnd vpwr scs8hd_fill_1
XFILLER_88_32 vgnd vpwr scs8hd_decap_12
XFILLER_144_93 vgnd vpwr scs8hd_decap_12
X_10_ _12_/A enable address[3] _13_/D _10_/X vgnd vpwr scs8hd_and4_4
XPHY_219 vgnd vpwr scs8hd_decap_3
XPHY_208 vgnd vpwr scs8hd_decap_3
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_149_27 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_165_59 vpwr vgnd scs8hd_fill_2
XFILLER_165_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_110 vgnd vpwr scs8hd_decap_12
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XFILLER_74_56 vgnd vpwr scs8hd_decap_12
XPHY_764 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_753 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_742 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_731 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_720 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_90_44 vgnd vpwr scs8hd_decap_12
XFILLER_99_86 vgnd vpwr scs8hd_decap_12
XFILLER_0_75 vgnd vpwr scs8hd_decap_6
XFILLER_80_105 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_151_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_100_32 vgnd vpwr scs8hd_decap_12
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XFILLER_109_74 vgnd vpwr scs8hd_decap_12
XFILLER_107_3 vgnd vpwr scs8hd_decap_12
XFILLER_125_62 vgnd vpwr scs8hd_decap_12
XFILLER_125_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XPHY_594 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_583 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_572 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_80 vgnd vpwr scs8hd_decap_12
XFILLER_50_80 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_162_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_44_105 vgnd vpwr scs8hd_fill_1
XFILLER_111_86 vgnd vpwr scs8hd_decap_12
XFILLER_121_110 vgnd vpwr scs8hd_decap_12
XFILLER_96_32 vgnd vpwr scs8hd_decap_12
XFILLER_152_93 vgnd vpwr scs8hd_decap_12
XPHY_380 vgnd vpwr scs8hd_decap_3
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XFILLER_179_110 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_173_15 vgnd vpwr scs8hd_decap_12
XFILLER_157_27 vgnd vpwr scs8hd_decap_12
XFILLER_173_59 vpwr vgnd scs8hd_fill_2
XFILLER_66_68 vgnd vpwr scs8hd_decap_12
XFILLER_174_3 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _10_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_82_56 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_182_105 vgnd vpwr scs8hd_decap_12
XFILLER_168_15 vgnd vpwr scs8hd_decap_12
XFILLER_117_74 vgnd vpwr scs8hd_decap_12
XFILLER_133_62 vgnd vpwr scs8hd_decap_12
XFILLER_133_51 vgnd vpwr scs8hd_decap_8
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_8
XFILLER_174_80 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vpwr vgnd scs8hd_fill_2
XFILLER_164_105 vgnd vpwr scs8hd_decap_12
XFILLER_170_27 vgnd vpwr scs8hd_decap_4
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XFILLER_103_98 vgnd vpwr scs8hd_decap_12
XFILLER_137_3 vgnd vpwr scs8hd_decap_12
XFILLER_88_44 vgnd vpwr scs8hd_decap_12
XFILLER_160_93 vgnd vpwr scs8hd_decap_12
XFILLER_146_105 vgnd vpwr scs8hd_decap_12
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_decap_3
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XFILLER_165_27 vgnd vpwr scs8hd_decap_12
XFILLER_149_39 vgnd vpwr scs8hd_decap_12
XFILLER_3_107 vgnd vpwr scs8hd_decap_3
XFILLER_181_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_118 vgnd vpwr scs8hd_decap_4
XFILLER_181_59 vpwr vgnd scs8hd_fill_2
XFILLER_74_68 vgnd vpwr scs8hd_decap_12
XPHY_765 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_754 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_743 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_732 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_721 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_710 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_128_105 vgnd vpwr scs8hd_decap_12
XFILLER_90_56 vgnd vpwr scs8hd_decap_12
XFILLER_99_98 vgnd vpwr scs8hd_decap_12
XFILLER_23_94 vpwr vgnd scs8hd_fill_2
XFILLER_48_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_80_117 vgnd vpwr scs8hd_decap_8
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_100_44 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_176_15 vgnd vpwr scs8hd_decap_12
XFILLER_109_86 vgnd vpwr scs8hd_decap_12
XFILLER_125_74 vgnd vpwr scs8hd_decap_12
XFILLER_141_62 vgnd vpwr scs8hd_decap_12
XFILLER_141_51 vgnd vpwr scs8hd_decap_8
XFILLER_62_117 vgnd vpwr scs8hd_decap_8
XPHY_595 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_584 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_573 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_182_80 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_111_98 vgnd vpwr scs8hd_decap_12
XFILLER_96_44 vgnd vpwr scs8hd_decap_12
XPHY_370 vgnd vpwr scs8hd_decap_3
XPHY_381 vgnd vpwr scs8hd_decap_3
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_157_39 vgnd vpwr scs8hd_decap_12
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_173_27 vgnd vpwr scs8hd_decap_12
XFILLER_106_32 vgnd vpwr scs8hd_decap_12
XFILLER_167_3 vgnd vpwr scs8hd_decap_12
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_82_68 vgnd vpwr scs8hd_decap_12
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
XFILLER_191_106 vgnd vpwr scs8hd_decap_12
XFILLER_82_3 vgnd vpwr scs8hd_decap_12
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_184_15 vgnd vpwr scs8hd_decap_12
XFILLER_182_117 vgnd vpwr scs8hd_decap_8
XFILLER_168_27 vgnd vpwr scs8hd_decap_4
XFILLER_117_86 vgnd vpwr scs8hd_decap_12
XFILLER_133_74 vgnd vpwr scs8hd_decap_12
XFILLER_158_93 vgnd vpwr scs8hd_decap_12
XFILLER_42_93 vgnd vpwr scs8hd_decap_12
XFILLER_190_80 vgnd vpwr scs8hd_decap_12
XFILLER_95_123 vpwr vgnd scs8hd_fill_2
XFILLER_164_117 vgnd vpwr scs8hd_decap_8
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _15_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_179_59 vpwr vgnd scs8hd_fill_2
XFILLER_179_15 vgnd vpwr scs8hd_decap_12
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_77_123 vpwr vgnd scs8hd_fill_2
XFILLER_88_56 vgnd vpwr scs8hd_decap_12
XFILLER_146_117 vgnd vpwr scs8hd_decap_8
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
XFILLER_165_39 vgnd vpwr scs8hd_decap_12
XFILLER_181_27 vgnd vpwr scs8hd_decap_12
XFILLER_114_32 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_123 vpwr vgnd scs8hd_fill_2
XPHY_711 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_700 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_766 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_755 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_744 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_733 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_722 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_139_62 vgnd vpwr scs8hd_decap_12
XFILLER_139_51 vgnd vpwr scs8hd_decap_8
XFILLER_128_117 vgnd vpwr scs8hd_decap_8
XFILLER_90_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_64_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_176_27 vgnd vpwr scs8hd_decap_4
XFILLER_100_56 vgnd vpwr scs8hd_decap_12
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_109_98 vgnd vpwr scs8hd_decap_12
XFILLER_125_86 vgnd vpwr scs8hd_decap_12
XFILLER_141_74 vgnd vpwr scs8hd_decap_12
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_596 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_585 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_574 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_93 vgnd vpwr scs8hd_decap_12
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_166_93 vgnd vpwr scs8hd_decap_12
XFILLER_53_118 vgnd vpwr scs8hd_decap_4
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
XFILLER_71_15 vgnd vpwr scs8hd_decap_12
XFILLER_187_59 vpwr vgnd scs8hd_fill_2
XFILLER_187_15 vgnd vpwr scs8hd_decap_12
XFILLER_112_3 vgnd vpwr scs8hd_decap_12
XFILLER_71_59 vpwr vgnd scs8hd_fill_2
XFILLER_121_123 vpwr vgnd scs8hd_fill_2
XFILLER_96_56 vgnd vpwr scs8hd_decap_12
XPHY_382 vgnd vpwr scs8hd_decap_3
XPHY_371 vgnd vpwr scs8hd_decap_3
XPHY_360 vgnd vpwr scs8hd_decap_3
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_6_ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_ebufn_1
XFILLER_179_123 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_173_39 vgnd vpwr scs8hd_decap_12
XFILLER_106_44 vgnd vpwr scs8hd_decap_12
XFILLER_103_123 vpwr vgnd scs8hd_fill_2
XFILLER_122_32 vgnd vpwr scs8hd_decap_12
XFILLER_66_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_147_62 vgnd vpwr scs8hd_decap_12
XFILLER_147_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_191_118 vgnd vpwr scs8hd_decap_6
XFILLER_188_80 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_decap_3
XFILLER_72_80 vgnd vpwr scs8hd_decap_12
XFILLER_75_3 vgnd vpwr scs8hd_decap_12
XFILLER_184_27 vgnd vpwr scs8hd_decap_4
XFILLER_117_98 vgnd vpwr scs8hd_decap_8
XFILLER_89_110 vgnd vpwr scs8hd_decap_12
XFILLER_133_86 vgnd vpwr scs8hd_decap_12
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XFILLER_174_93 vgnd vpwr scs8hd_decap_12
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_179_27 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_8
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_88_68 vgnd vpwr scs8hd_decap_12
XFILLER_92_105 vgnd vpwr scs8hd_decap_12
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_124 vgnd vpwr scs8hd_fill_1
XFILLER_181_39 vgnd vpwr scs8hd_decap_12
XFILLER_114_44 vgnd vpwr scs8hd_decap_12
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XFILLER_74_15 vgnd vpwr scs8hd_decap_12
XFILLER_74_105 vgnd vpwr scs8hd_decap_12
XPHY_745 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_734 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_723 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_712 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_701 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_130_32 vgnd vpwr scs8hd_decap_12
XPHY_767 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_756 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_142_3 vgnd vpwr scs8hd_decap_12
XFILLER_139_74 vgnd vpwr scs8hd_decap_12
XFILLER_155_62 vgnd vpwr scs8hd_decap_12
XFILLER_155_51 vgnd vpwr scs8hd_decap_8
XFILLER_151_121 vgnd vpwr scs8hd_fill_1
XFILLER_151_110 vgnd vpwr scs8hd_decap_3
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_48_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XFILLER_80_80 vgnd vpwr scs8hd_decap_12
XFILLER_56_105 vgnd vpwr scs8hd_decap_12
XFILLER_100_68 vgnd vpwr scs8hd_decap_12
XFILLER_133_110 vgnd vpwr scs8hd_decap_12
XFILLER_69_15 vgnd vpwr scs8hd_decap_12
XFILLER_69_59 vpwr vgnd scs8hd_fill_2
XFILLER_125_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
XFILLER_141_86 vgnd vpwr scs8hd_decap_12
XPHY_586 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_575 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_597 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_182_93 vgnd vpwr scs8hd_decap_12
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_115_110 vgnd vpwr scs8hd_decap_12
XFILLER_44_108 vgnd vpwr scs8hd_decap_12
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
XFILLER_187_27 vgnd vpwr scs8hd_decap_12
XFILLER_71_27 vgnd vpwr scs8hd_decap_12
XFILLER_105_3 vgnd vpwr scs8hd_decap_12
XFILLER_96_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XPHY_383 vgnd vpwr scs8hd_decap_3
XPHY_372 vgnd vpwr scs8hd_decap_3
XPHY_361 vgnd vpwr scs8hd_decap_3
XPHY_350 vgnd vpwr scs8hd_decap_3
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_106_56 vgnd vpwr scs8hd_decap_12
XFILLER_66_27 vgnd vpwr scs8hd_decap_4
XFILLER_122_44 vgnd vpwr scs8hd_decap_12
XFILLER_82_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_147_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_163_62 vgnd vpwr scs8hd_decap_12
XFILLER_163_51 vgnd vpwr scs8hd_decap_8
XFILLER_176_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_111 vgnd vpwr scs8hd_decap_8
XFILLER_56_93 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_decap_3
XPHY_180 vgnd vpwr scs8hd_decap_3
XFILLER_68_3 vgnd vpwr scs8hd_decap_12
XFILLER_100_105 vgnd vpwr scs8hd_decap_12
.ends

