* NGSPICE file created from sb_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_1__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable left_bottom_grid_pin_12_ left_top_grid_pin_10_ right_bottom_grid_pin_12_
+ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_ vpwr vgnd
XFILLER_39_211 vpwr vgnd scs8hd_fill_2
XFILLER_36_19 vgnd vpwr scs8hd_decap_12
XFILLER_22_144 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__203__B _205_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_111 vgnd vpwr scs8hd_decap_6
XFILLER_9_104 vpwr vgnd scs8hd_fill_2
XFILLER_9_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_6_.latch data_in mem_left_track_1.LATCH_6_.latch/Q _190_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _215_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__214__A _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_3
XFILLER_18_247 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__B _220_/A vgnd vpwr scs8hd_diode_2
X_277_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A _099_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XFILLER_5_195 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _241_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__209__A _208_/X vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _205_/B _200_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
X_131_ _130_/X _123_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_33 vpwr vgnd scs8hd_fill_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _229_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _274_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__211__B _211_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_97 vpwr vgnd scs8hd_fill_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_7_213 vgnd vpwr scs8hd_decap_3
XFILLER_11_220 vgnd vpwr scs8hd_decap_3
X_114_ _114_/A _114_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_7 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_37_161 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_43 vgnd vpwr scs8hd_decap_8
XFILLER_20_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_249 vgnd vpwr scs8hd_fill_1
XANTENNA__206__B _198_/X vgnd vpwr scs8hd_diode_2
XANTENNA__222__A _114_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_109 vgnd vpwr scs8hd_decap_4
XFILLER_28_183 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _132_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_186 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _161_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_101 vpwr vgnd scs8hd_fill_2
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_15_21 vpwr vgnd scs8hd_fill_2
XANTENNA__217__A _217_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_53 vgnd vpwr scs8hd_decap_4
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XFILLER_31_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _203_/Y vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _241_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_64 vgnd vpwr scs8hd_decap_4
XFILLER_9_116 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vpwr vgnd scs8hd_fill_2
XFILLER_13_178 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_6_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_193 vpwr vgnd scs8hd_fill_2
XFILLER_27_226 vpwr vgnd scs8hd_fill_2
XFILLER_27_215 vpwr vgnd scs8hd_fill_2
XFILLER_27_204 vpwr vgnd scs8hd_fill_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_104 vgnd vpwr scs8hd_decap_8
XFILLER_12_66 vpwr vgnd scs8hd_fill_2
XANTENNA__214__B _211_/B vgnd vpwr scs8hd_diode_2
XANTENNA__230__A _114_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_226 vpwr vgnd scs8hd_fill_2
X_276_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__140__A _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_270 vgnd vpwr scs8hd_decap_6
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_6_.latch data_in mem_top_track_8.LATCH_6_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_6_.latch data_in mem_right_track_0.LATCH_6_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_207 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _251_/HI mem_top_track_8.LATCH_7_.latch/Q
+ mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _107_/A _130_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__225__A _224_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_199 vgnd vpwr scs8hd_decap_4
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_259_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_97 vgnd vpwr scs8hd_fill_1
XFILLER_7_203 vgnd vpwr scs8hd_fill_1
XFILLER_11_254 vgnd vpwr scs8hd_decap_4
XFILLER_11_265 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A _114_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _196_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_7 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__222__B _220_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_20_11 vgnd vpwr scs8hd_fill_1
XFILLER_4_206 vgnd vpwr scs8hd_decap_6
XFILLER_4_228 vgnd vpwr scs8hd_decap_4
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_6_46 vpwr vgnd scs8hd_fill_2
XFILLER_6_79 vgnd vpwr scs8hd_decap_12
XFILLER_34_110 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _223_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_34_198 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__233__A _232_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_87 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_132 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_135 vpwr vgnd scs8hd_fill_2
XFILLER_31_102 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _123_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_165 vgnd vpwr scs8hd_decap_8
XFILLER_16_187 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vpwr vgnd scs8hd_fill_2
XFILLER_22_102 vgnd vpwr scs8hd_decap_3
XFILLER_26_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__228__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _270_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_7_.latch data_in mem_left_track_9.LATCH_7_.latch/Q _200_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_161 vpwr vgnd scs8hd_fill_2
XFILLER_6_109 vpwr vgnd scs8hd_fill_2
XFILLER_10_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_45 vpwr vgnd scs8hd_fill_2
XFILLER_12_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__230__B _231_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_97 vpwr vgnd scs8hd_fill_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
X_275_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_5_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_219 vpwr vgnd scs8hd_fill_2
XFILLER_23_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_252 vpwr vgnd scs8hd_fill_2
XFILLER_23_241 vgnd vpwr scs8hd_decap_3
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_3
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XFILLER_2_112 vpwr vgnd scs8hd_fill_2
XFILLER_2_101 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_13 vgnd vpwr scs8hd_decap_3
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
X_258_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
X_189_ _200_/A _188_/X _189_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_211 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_34_43 vgnd vpwr scs8hd_fill_1
XFILLER_34_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__236__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_237 vgnd vpwr scs8hd_fill_1
X_112_ address[1] address[2] _106_/C _113_/A vgnd vpwr scs8hd_or3_4
XANTENNA__146__A _130_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_152 vgnd vpwr scs8hd_decap_4
XFILLER_37_141 vpwr vgnd scs8hd_fill_2
XFILLER_37_130 vpwr vgnd scs8hd_fill_2
XFILLER_1_91 vpwr vgnd scs8hd_fill_2
XFILLER_20_67 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_6_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_76 vgnd vpwr scs8hd_decap_4
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_196 vgnd vpwr scs8hd_decap_12
XFILLER_6_58 vgnd vpwr scs8hd_decap_4
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_100 vgnd vpwr scs8hd_fill_1
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_66 vgnd vpwr scs8hd_decap_4
XFILLER_31_11 vgnd vpwr scs8hd_decap_3
XFILLER_0_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _240_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_144 vgnd vpwr scs8hd_decap_6
XFILLER_31_147 vgnd vpwr scs8hd_fill_1
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_136 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
XANTENNA__228__B _231_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_206 vgnd vpwr scs8hd_decap_8
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__154__A _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_206 vgnd vpwr scs8hd_decap_6
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_76 vgnd vpwr scs8hd_decap_4
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_274_ _274_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _117_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_7_.latch data_in mem_right_track_8.LATCH_7_.latch/Q _155_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_275 vpwr vgnd scs8hd_fill_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XFILLER_2_168 vpwr vgnd scs8hd_fill_2
XFILLER_2_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _236_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_257_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_188_ _187_/X _188_/X vgnd vpwr scs8hd_buf_1
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
XANTENNA__151__B _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_201 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_45 vgnd vpwr scs8hd_decap_4
XFILLER_18_23 vgnd vpwr scs8hd_decap_6
XFILLER_34_88 vpwr vgnd scs8hd_fill_2
XFILLER_34_77 vgnd vpwr scs8hd_decap_4
XANTENNA__236__B _233_/X vgnd vpwr scs8hd_diode_2
XANTENNA__252__A _252_/A vgnd vpwr scs8hd_diode_2
X_111_ _114_/A _237_/A _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__146__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_66 vgnd vpwr scs8hd_fill_1
XFILLER_28_186 vgnd vpwr scs8hd_fill_1
XFILLER_28_164 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_131 vpwr vgnd scs8hd_fill_2
XFILLER_20_7 vgnd vpwr scs8hd_decap_4
XFILLER_34_145 vgnd vpwr scs8hd_decap_8
XFILLER_34_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _127_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XFILLER_25_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_46 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_68 vpwr vgnd scs8hd_fill_2
XFILLER_31_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_215 vgnd vpwr scs8hd_decap_4
XFILLER_39_204 vgnd vpwr scs8hd_decap_3
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _195_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_23 vgnd vpwr scs8hd_decap_8
XFILLER_26_12 vgnd vpwr scs8hd_decap_8
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_108 vgnd vpwr scs8hd_fill_1
XFILLER_13_148 vgnd vpwr scs8hd_fill_1
XANTENNA__260__A _260_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_38 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_174 vpwr vgnd scs8hd_fill_2
XFILLER_12_181 vgnd vpwr scs8hd_decap_8
XANTENNA__170__A _130_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _221_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XANTENNA__239__B _233_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_262 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_8
XFILLER_26_240 vgnd vpwr scs8hd_decap_8
XANTENNA__255__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_273_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_5_111 vpwr vgnd scs8hd_fill_2
XFILLER_5_177 vgnd vpwr scs8hd_decap_4
XFILLER_5_199 vpwr vgnd scs8hd_fill_2
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_39 vpwr vgnd scs8hd_fill_2
XFILLER_9_37 vgnd vpwr scs8hd_decap_3
XFILLER_14_243 vpwr vgnd scs8hd_fill_2
XFILLER_14_254 vgnd vpwr scs8hd_decap_8
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/X vgnd vpwr scs8hd_buf_1
X_256_ _256_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_13_90 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_246 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_4
X_110_ _132_/A _237_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_239_ _239_/A _233_/X _239_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _153_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_25 vgnd vpwr scs8hd_decap_4
XFILLER_29_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_3
XFILLER_28_110 vgnd vpwr scs8hd_decap_8
XANTENNA__263__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _206_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_25 vpwr vgnd scs8hd_fill_2
XANTENNA__258__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_113 vgnd vpwr scs8hd_decap_6
XFILLER_16_124 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_227 vgnd vpwr scs8hd_decap_4
XANTENNA__168__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_182 vpwr vgnd scs8hd_fill_2
XFILLER_30_193 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_68 vgnd vpwr scs8hd_fill_1
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_17 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_197 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_4
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_23 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_272_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XANTENNA__271__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _135_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_211 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_60 vpwr vgnd scs8hd_fill_2
XANTENNA__181__A _130_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_233 vpwr vgnd scs8hd_fill_2
XFILLER_23_222 vpwr vgnd scs8hd_fill_2
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__266__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
X_255_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_14_266 vgnd vpwr scs8hd_decap_8
X_186_ _152_/A _232_/B _152_/C _224_/D _187_/A vgnd vpwr scs8hd_or4_4
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_269 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_58 vgnd vpwr scs8hd_decap_4
XFILLER_34_46 vgnd vpwr scs8hd_fill_1
XFILLER_7_218 vpwr vgnd scs8hd_fill_2
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_258 vgnd vpwr scs8hd_fill_1
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XANTENNA__086__A _085_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_238_ _114_/B _233_/X _238_/Y vgnd vpwr scs8hd_nor2_4
X_169_ _128_/X _165_/X _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_188 vgnd vpwr scs8hd_decap_12
XFILLER_1_50 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _210_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_100 vgnd vpwr scs8hd_fill_1
XFILLER_28_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_199 vgnd vpwr scs8hd_decap_4
XFILLER_19_177 vgnd vpwr scs8hd_decap_4
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_169 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_6_.latch data_in mem_top_track_0.LATCH_6_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__173__B _164_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _181_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_40_106 vgnd vpwr scs8hd_decap_8
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_33_191 vgnd vpwr scs8hd_decap_4
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_139 vpwr vgnd scs8hd_fill_2
XFILLER_31_106 vgnd vpwr scs8hd_decap_3
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__274__A _274_/A vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_239 vgnd vpwr scs8hd_decap_4
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_82 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _205_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_47 vgnd vpwr scs8hd_decap_4
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_117 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_161 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_8_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__269__A _269_/A vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XFILLER_12_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _227_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_37_35 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _212_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
X_271_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__181__B _180_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
XFILLER_4_83 vgnd vpwr scs8hd_decap_3
XFILLER_23_201 vgnd vpwr scs8hd_decap_8
XFILLER_2_127 vpwr vgnd scs8hd_fill_2
XFILLER_2_116 vpwr vgnd scs8hd_fill_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
XANTENNA__282__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_254_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
X_185_ address[5] _150_/Y _224_/D vgnd vpwr scs8hd_or2_4
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_7 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vpwr vgnd scs8hd_fill_2
XANTENNA__192__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_7_.latch data_in mem_left_track_1.LATCH_7_.latch/Q _189_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__277__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_8_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_237_ _237_/A _233_/X _237_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_track_9.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_168_ _127_/A _165_/X _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_099_ _114_/A _099_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_112 vpwr vgnd scs8hd_fill_2
XFILLER_37_101 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_fill_1
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_6_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_36 vgnd vpwr scs8hd_decap_6
XANTENNA__097__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_266 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_156 vgnd vpwr scs8hd_decap_3
XFILLER_19_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_38 vpwr vgnd scs8hd_fill_2
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _228_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_107 vgnd vpwr scs8hd_decap_3
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__184__B _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_94 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _191_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__285__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_80 vgnd vpwr scs8hd_fill_1
XFILLER_8_133 vgnd vpwr scs8hd_decap_3
XFILLER_16_81 vgnd vpwr scs8hd_decap_8
XANTENNA__179__B _180_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_243 vgnd vpwr scs8hd_fill_1
XANTENNA__195__A _135_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_37_47 vgnd vpwr scs8hd_decap_3
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
X_270_ _270_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_5_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _218_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
XFILLER_4_40 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_202 vpwr vgnd scs8hd_fill_2
X_253_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_184_ _149_/A _176_/A _184_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_161 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_6_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_20_205 vgnd vpwr scs8hd_decap_6
XANTENNA__192__B _188_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_205 vpwr vgnd scs8hd_fill_2
XFILLER_11_216 vpwr vgnd scs8hd_fill_2
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_236_ _220_/A _233_/X _236_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_242 vgnd vpwr scs8hd_decap_3
X_167_ _125_/A _165_/X _167_/Y vgnd vpwr scs8hd_nor2_4
X_098_ _097_/X _099_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_179 vgnd vpwr scs8hd_decap_4
XFILLER_1_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__097__B _103_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _236_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_223 vgnd vpwr scs8hd_fill_1
XFILLER_3_212 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_7_.latch data_in mem_right_track_0.LATCH_7_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_72 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_7_.latch data_in mem_top_track_8.LATCH_7_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_168 vgnd vpwr scs8hd_decap_3
X_219_ _211_/A _220_/B _219_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_127 vgnd vpwr scs8hd_fill_1
XFILLER_25_116 vgnd vpwr scs8hd_decap_4
XFILLER_18_190 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _250_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _245_/HI mem_left_track_9.LATCH_7_.latch/Q
+ mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_119 vgnd vpwr scs8hd_decap_8
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_decap_4
XFILLER_15_193 vgnd vpwr scs8hd_decap_4
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _244_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_123 vgnd vpwr scs8hd_fill_1
XFILLER_8_145 vgnd vpwr scs8hd_decap_8
XFILLER_8_178 vpwr vgnd scs8hd_fill_2
XFILLER_12_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__195__B _187_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _260_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_252_ _252_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _135_/A _176_/A _183_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_72 vgnd vpwr scs8hd_decap_3
XFILLER_13_94 vpwr vgnd scs8hd_fill_2
XFILLER_29_8 vpwr vgnd scs8hd_fill_2
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_273 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_235_ _211_/A _233_/X _235_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XFILLER_6_210 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_232 vgnd vpwr scs8hd_fill_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_10_272 vgnd vpwr scs8hd_decap_3
X_166_ _123_/A _165_/X _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _106_/A _103_/B address[0] _097_/X vgnd vpwr scs8hd_or3_4
XFILLER_1_20 vpwr vgnd scs8hd_fill_2
XFILLER_37_169 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__097__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_235 vgnd vpwr scs8hd_decap_3
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_4
XFILLER_35_92 vpwr vgnd scs8hd_fill_2
XFILLER_34_128 vgnd vpwr scs8hd_decap_4
X_218_ _234_/A _220_/B _218_/Y vgnd vpwr scs8hd_nor2_4
X_149_ _149_/A _149_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_106 vgnd vpwr scs8hd_decap_4
XFILLER_33_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_128 vpwr vgnd scs8hd_fill_2
XFILLER_24_183 vpwr vgnd scs8hd_fill_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_30_142 vgnd vpwr scs8hd_decap_8
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_186 vgnd vpwr scs8hd_decap_4
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_197 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XFILLER_8_113 vpwr vgnd scs8hd_fill_2
XFILLER_8_157 vpwr vgnd scs8hd_fill_2
XFILLER_12_164 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_160 vpwr vgnd scs8hd_fill_2
XFILLER_4_171 vpwr vgnd scs8hd_fill_2
XFILLER_4_64 vpwr vgnd scs8hd_fill_2
XFILLER_4_75 vpwr vgnd scs8hd_fill_2
XFILLER_23_259 vpwr vgnd scs8hd_fill_2
XFILLER_23_248 vpwr vgnd scs8hd_fill_2
XFILLER_23_237 vpwr vgnd scs8hd_fill_2
XFILLER_23_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_251_ _251_/HI _251_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_182_ _133_/A _180_/B _182_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_237 vgnd vpwr scs8hd_decap_4
XFILLER_13_62 vgnd vpwr scs8hd_fill_1
XFILLER_38_70 vpwr vgnd scs8hd_fill_2
XFILLER_1_174 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_229 vgnd vpwr scs8hd_decap_8
XFILLER_9_241 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_39 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _240_/HI mem_bottom_track_1.LATCH_7_.latch/Q
+ mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_165_ _164_/X _165_/X vgnd vpwr scs8hd_buf_1
X_234_ _234_/A _233_/X _234_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _213_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_8
X_096_ _117_/A _114_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_148 vpwr vgnd scs8hd_fill_2
XFILLER_37_137 vpwr vgnd scs8hd_fill_2
XFILLER_37_126 vpwr vgnd scs8hd_fill_2
XFILLER_1_54 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _114_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_170 vgnd vpwr scs8hd_decap_12
XFILLER_28_148 vgnd vpwr scs8hd_decap_4
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
XFILLER_34_118 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_217_ _217_/A _220_/B vgnd vpwr scs8hd_buf_1
X_148_ _135_/A _149_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_162 vgnd vpwr scs8hd_fill_1
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _235_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_228 vpwr vgnd scs8hd_fill_2
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XFILLER_24_140 vgnd vpwr scs8hd_decap_8
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_21_95 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_165 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_140 vgnd vpwr scs8hd_fill_1
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_165 vgnd vpwr scs8hd_decap_4
XFILLER_12_154 vgnd vpwr scs8hd_fill_1
XFILLER_16_62 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _230_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__103__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_235 vpwr vgnd scs8hd_fill_2
XFILLER_17_224 vpwr vgnd scs8hd_fill_2
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_54 vgnd vpwr scs8hd_decap_4
XFILLER_4_183 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB _201_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_19 vpwr vgnd scs8hd_fill_2
X_250_ _250_/HI _250_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
X_181_ _130_/X _180_/B _181_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_142 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _194_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__100__B _103_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_219 vgnd vpwr scs8hd_fill_1
XFILLER_9_220 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _099_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _220_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_51 vgnd vpwr scs8hd_decap_6
XFILLER_24_40 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_233_ _232_/X _233_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_164_ _163_/X _164_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_84 vgnd vpwr scs8hd_decap_6
X_095_ _123_/A _117_/A _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XFILLER_37_116 vgnd vpwr scs8hd_decap_6
XANTENNA__111__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_33 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_182 vgnd vpwr scs8hd_decap_12
XFILLER_36_160 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_20 vpwr vgnd scs8hd_fill_2
XFILLER_10_53 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_127 vpwr vgnd scs8hd_fill_2
XFILLER_19_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_73 vpwr vgnd scs8hd_fill_2
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ _133_/A _142_/B _147_/Y vgnd vpwr scs8hd_nor2_4
X_216_ _152_/A _232_/B _232_/C _152_/D _217_/A vgnd vpwr scs8hd_or4_4
XFILLER_31_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_fill_1
XFILLER_24_163 vgnd vpwr scs8hd_decap_3
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_85 vpwr vgnd scs8hd_fill_2
XFILLER_21_74 vpwr vgnd scs8hd_fill_2
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _194_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_122 vgnd vpwr scs8hd_fill_1
XFILLER_30_111 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_32 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_8_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_87 vpwr vgnd scs8hd_fill_2
XFILLER_7_98 vpwr vgnd scs8hd_fill_2
XFILLER_38_200 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_96 vgnd vpwr scs8hd_decap_8
XFILLER_32_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _221_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__204__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XFILLER_27_51 vpwr vgnd scs8hd_fill_2
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XFILLER_4_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_180_ _128_/X _180_/B _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_31 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__100__C _106_/C vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _243_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_209 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_180 vgnd vpwr scs8hd_fill_1
XANTENNA__201__B _205_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_74 vpwr vgnd scs8hd_fill_2
X_232_ _232_/A _232_/B _232_/C _224_/D _232_/X vgnd vpwr scs8hd_or4_4
X_094_ _094_/A _117_/A vgnd vpwr scs8hd_buf_1
X_163_ _232_/C _152_/D _232_/A _152_/B _163_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_202 vpwr vgnd scs8hd_fill_2
XFILLER_6_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_253 vgnd vpwr scs8hd_decap_8
XFILLER_10_264 vgnd vpwr scs8hd_decap_8
XANTENNA__111__B _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _239_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _133_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _147_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_19 vpwr vgnd scs8hd_fill_2
XFILLER_36_194 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_216 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__212__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_40 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_62 vpwr vgnd scs8hd_fill_2
X_215_ _239_/A _211_/B _215_/Y vgnd vpwr scs8hd_nor2_4
X_146_ _130_/X _142_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__106__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_6 vgnd vpwr scs8hd_decap_12
XFILLER_18_194 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _239_/A vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vgnd vpwr scs8hd_fill_1
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_66 vgnd vpwr scs8hd_fill_1
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
X_129_ _128_/X _123_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_74 vgnd vpwr scs8hd_decap_6
XFILLER_8_138 vpwr vgnd scs8hd_fill_2
XFILLER_12_134 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_189 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__103__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_215 vgnd vpwr scs8hd_decap_12
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_7_.latch data_in mem_top_track_0.LATCH_7_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _180_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__204__B _205_/B vgnd vpwr scs8hd_diode_2
XANTENNA__220__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_30 vpwr vgnd scs8hd_fill_2
XFILLER_17_204 vgnd vpwr scs8hd_decap_3
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _114_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _107_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_218 vgnd vpwr scs8hd_decap_6
XANTENNA__215__A _239_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _204_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_188 vgnd vpwr scs8hd_decap_3
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
XFILLER_9_233 vpwr vgnd scs8hd_fill_2
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XFILLER_13_273 vgnd vpwr scs8hd_decap_4
XANTENNA__109__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vgnd vpwr scs8hd_decap_12
XFILLER_39_170 vpwr vgnd scs8hd_fill_2
X_231_ _239_/A _231_/B _231_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_162_ _149_/A _153_/X _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_221 vpwr vgnd scs8hd_fill_2
X_093_ _152_/A _152_/B _232_/C _208_/D _094_/A vgnd vpwr scs8hd_or4_4
XFILLER_6_247 vgnd vpwr scs8hd_decap_3
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _211_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__212__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vgnd vpwr scs8hd_decap_3
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_10_88 vgnd vpwr scs8hd_fill_1
XFILLER_27_140 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XFILLER_35_96 vpwr vgnd scs8hd_fill_2
X_214_ _114_/B _211_/B _214_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _128_/X _142_/B _145_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XFILLER_33_198 vpwr vgnd scs8hd_fill_2
XFILLER_33_187 vpwr vgnd scs8hd_fill_2
XFILLER_33_176 vgnd vpwr scs8hd_fill_1
XFILLER_33_154 vpwr vgnd scs8hd_fill_2
XFILLER_33_143 vpwr vgnd scs8hd_fill_2
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_121 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_187 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__B _198_/X vgnd vpwr scs8hd_diode_2
XANTENNA__223__A _239_/A vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_154 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _239_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _128_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_78 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XANTENNA__218__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_32_53 vgnd vpwr scs8hd_decap_4
XFILLER_8_106 vgnd vpwr scs8hd_decap_4
XFILLER_8_117 vgnd vpwr scs8hd_decap_6
XFILLER_12_168 vgnd vpwr scs8hd_decap_4
XFILLER_35_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_150 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__220__B _220_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_131 vgnd vpwr scs8hd_fill_1
XFILLER_4_175 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_79 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _227_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_241 vgnd vpwr scs8hd_decap_3
XFILLER_22_241 vgnd vpwr scs8hd_decap_4
XANTENNA__215__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_55 vpwr vgnd scs8hd_fill_2
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XANTENNA__231__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_178 vgnd vpwr scs8hd_decap_3
XFILLER_1_112 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vpwr vgnd scs8hd_fill_2
XFILLER_38_74 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA__109__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _248_/HI mem_right_track_8.LATCH_7_.latch/Q
+ mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_160 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
X_230_ _114_/B _231_/B _230_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_200 vgnd vpwr scs8hd_decap_12
X_161_ _135_/A _153_/X _161_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__226__A _234_/A vgnd vpwr scs8hd_diode_2
X_092_ address[5] address[6] _208_/D vgnd vpwr scs8hd_or2_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_259 vpwr vgnd scs8hd_fill_2
XFILLER_37_108 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_45 vpwr vgnd scs8hd_fill_2
XFILLER_10_67 vgnd vpwr scs8hd_decap_3
XFILLER_19_21 vpwr vgnd scs8hd_fill_2
XFILLER_19_10 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_174 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _237_/A _211_/B _213_/Y vgnd vpwr scs8hd_nor2_4
X_144_ _127_/A _142_/B _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_111 vgnd vpwr scs8hd_decap_8
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_55 vpwr vgnd scs8hd_fill_2
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XANTENNA__223__B _220_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_100 vpwr vgnd scs8hd_fill_2
XFILLER_30_169 vgnd vpwr scs8hd_decap_4
XFILLER_30_125 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_127_ _127_/A _123_/B _127_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _278_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_169 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_6_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA__218__B _220_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_8
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_180 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_239 vgnd vpwr scs8hd_decap_4
XANTENNA__144__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _204_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__229__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_239 vgnd vpwr scs8hd_decap_3
XFILLER_17_228 vpwr vgnd scs8hd_fill_2
XFILLER_4_36 vpwr vgnd scs8hd_fill_2
XFILLER_4_143 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _249_/HI mem_top_track_0.LATCH_7_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_250 vpwr vgnd scs8hd_fill_2
XFILLER_31_275 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_64 vgnd vpwr scs8hd_decap_3
XANTENNA__231__B _231_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XFILLER_13_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _249_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_11 vgnd vpwr scs8hd_decap_4
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_091_ _091_/A _232_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_212 vpwr vgnd scs8hd_fill_2
X_160_ _133_/A _154_/X _160_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__226__B _231_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_219 vgnd vpwr scs8hd_decap_4
XFILLER_10_24 vpwr vgnd scs8hd_fill_2
XFILLER_27_120 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_212_ _220_/A _211_/B _212_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_197 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
X_143_ _125_/A _142_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_186 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _133_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.INVTX1_8_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_89 vgnd vpwr scs8hd_decap_4
XFILLER_21_78 vgnd vpwr scs8hd_decap_4
XFILLER_21_34 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_178 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _101_/A _127_/A vgnd vpwr scs8hd_buf_1
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_148 vpwr vgnd scs8hd_fill_2
XFILLER_29_226 vgnd vpwr scs8hd_decap_12
XFILLER_29_215 vgnd vpwr scs8hd_decap_8
XFILLER_29_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _246_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_16_45 vgnd vpwr scs8hd_decap_8
XFILLER_16_89 vgnd vpwr scs8hd_decap_3
XFILLER_32_88 vgnd vpwr scs8hd_decap_4
XANTENNA__234__B _233_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_163 vpwr vgnd scs8hd_fill_2
XFILLER_7_174 vpwr vgnd scs8hd_fill_2
XFILLER_11_192 vpwr vgnd scs8hd_fill_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_4
XANTENNA__160__A _133_/A vgnd vpwr scs8hd_diode_2
X_109_ _106_/A address[2] address[0] _132_/A vgnd vpwr scs8hd_or3_4
XFILLER_26_229 vgnd vpwr scs8hd_decap_8
XFILLER_26_218 vgnd vpwr scs8hd_decap_8
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vpwr vgnd scs8hd_fill_2
XFILLER_27_55 vgnd vpwr scs8hd_decap_4
XANTENNA__229__B _231_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_199 vgnd vpwr scs8hd_decap_4
XFILLER_31_221 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _232_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_240 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_22_210 vgnd vpwr scs8hd_fill_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_203 vpwr vgnd scs8hd_fill_2
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_9_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_4
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_24_78 vgnd vpwr scs8hd_decap_3
X_090_ enable _091_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
XFILLER_6_228 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_16 vpwr vgnd scs8hd_fill_2
XFILLER_1_38 vgnd vpwr scs8hd_decap_3
XANTENNA__152__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_11 vgnd vpwr scs8hd_decap_12
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_44 vgnd vpwr scs8hd_decap_4
X_211_ _211_/A _211_/B _211_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__237__B _233_/X vgnd vpwr scs8hd_diode_2
X_142_ _123_/A _142_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__253__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_2_253 vpwr vgnd scs8hd_fill_2
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
XFILLER_18_143 vgnd vpwr scs8hd_decap_8
XANTENNA__147__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _232_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_168 vgnd vpwr scs8hd_decap_6
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_138 vpwr vgnd scs8hd_fill_2
X_125_ _125_/A _123_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_15 vpwr vgnd scs8hd_fill_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XFILLER_21_116 vgnd vpwr scs8hd_decap_4
XFILLER_21_105 vgnd vpwr scs8hd_decap_4
XANTENNA__158__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_238 vgnd vpwr scs8hd_decap_6
XFILLER_32_23 vgnd vpwr scs8hd_decap_8
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_138 vgnd vpwr scs8hd_decap_4
X_108_ _114_/A _220_/A _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_171 vgnd vpwr scs8hd_fill_1
XFILLER_21_3 vgnd vpwr scs8hd_decap_3
XANTENNA__160__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _283_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_34 vpwr vgnd scs8hd_fill_2
XFILLER_27_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_200 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _234_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_123 vgnd vpwr scs8hd_decap_8
XANTENNA__261__A _261_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XANTENNA__139__C _152_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_233 vgnd vpwr scs8hd_decap_8
XANTENNA__155__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_14 vpwr vgnd scs8hd_fill_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA__256__A _256_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_237 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB _189_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_174 vgnd vpwr scs8hd_decap_6
XFILLER_39_152 vgnd vpwr scs8hd_decap_8
XFILLER_39_130 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_236 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
X_287_ _287_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__152__C _152_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_46 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_23 vgnd vpwr scs8hd_decap_12
XFILLER_27_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
X_210_ _234_/A _211_/B _210_/Y vgnd vpwr scs8hd_nor2_4
X_141_ _149_/B _142_/B vgnd vpwr scs8hd_buf_1
XFILLER_2_232 vpwr vgnd scs8hd_fill_2
XFILLER_2_210 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_111 vgnd vpwr scs8hd_decap_8
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_158 vpwr vgnd scs8hd_fill_2
XFILLER_33_147 vgnd vpwr scs8hd_decap_4
XANTENNA__163__B _152_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _193_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_125 vpwr vgnd scs8hd_fill_2
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_47 vpwr vgnd scs8hd_fill_2
XFILLER_15_136 vgnd vpwr scs8hd_decap_4
XFILLER_15_158 vpwr vgnd scs8hd_fill_2
XANTENNA__264__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_7_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_124_ _099_/B _125_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__158__B _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _219_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vgnd vpwr scs8hd_decap_12
XFILLER_32_68 vgnd vpwr scs8hd_decap_4
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__259__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _234_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
X_107_ _107_/A _220_/A vgnd vpwr scs8hd_buf_1
XANTENNA__169__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_209 vpwr vgnd scs8hd_fill_2
XFILLER_40_212 vpwr vgnd scs8hd_fill_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XFILLER_4_179 vgnd vpwr scs8hd_decap_4
XANTENNA__139__D _208_/D vgnd vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_116 vgnd vpwr scs8hd_decap_4
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__272__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__182__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_36 vpwr vgnd scs8hd_fill_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_4
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__267__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
X_286_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XFILLER_5_241 vgnd vpwr scs8hd_fill_1
XANTENNA__152__D _152_/D vgnd vpwr scs8hd_diode_2
XFILLER_36_145 vgnd vpwr scs8hd_decap_8
XANTENNA__177__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_49 vpwr vgnd scs8hd_fill_2
XFILLER_19_58 vgnd vpwr scs8hd_decap_3
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XFILLER_19_14 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_79 vpwr vgnd scs8hd_fill_2
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_35_35 vpwr vgnd scs8hd_fill_2
XFILLER_27_178 vgnd vpwr scs8hd_decap_3
XFILLER_27_123 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _200_/A vgnd vpwr scs8hd_diode_2
X_140_ _139_/X _149_/B vgnd vpwr scs8hd_buf_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_266 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_167 vgnd vpwr scs8hd_decap_8
XFILLER_18_101 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_269_ _269_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__163__C _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_148 vgnd vpwr scs8hd_fill_1
XFILLER_24_104 vgnd vpwr scs8hd_decap_8
XFILLER_21_15 vpwr vgnd scs8hd_fill_2
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_118 vgnd vpwr scs8hd_decap_4
XFILLER_30_107 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_104 vpwr vgnd scs8hd_fill_2
XFILLER_15_115 vgnd vpwr scs8hd_decap_4
XANTENNA__280__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
X_123_ _123_/A _123_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_8 vpwr vgnd scs8hd_fill_2
XFILLER_11_81 vpwr vgnd scs8hd_fill_2
XANTENNA__174__B _232_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _131_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _146_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_118 vgnd vpwr scs8hd_fill_1
XFILLER_20_184 vpwr vgnd scs8hd_fill_2
XFILLER_20_140 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__275__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _207_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_133 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
X_106_ _106_/A address[2] _106_/C _107_/A vgnd vpwr scs8hd_or3_4
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XANTENNA__169__B _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_210 vgnd vpwr scs8hd_decap_4
XANTENNA__185__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_82 vpwr vgnd scs8hd_fill_2
XFILLER_27_47 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_4
XFILLER_25_221 vpwr vgnd scs8hd_fill_2
XFILLER_25_210 vpwr vgnd scs8hd_fill_2
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_147 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_202 vpwr vgnd scs8hd_fill_2
XFILLER_16_254 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_90 vpwr vgnd scs8hd_fill_2
XFILLER_22_224 vpwr vgnd scs8hd_fill_2
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vgnd vpwr scs8hd_decap_4
XFILLER_13_224 vgnd vpwr scs8hd_fill_1
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__182__B _180_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_250 vpwr vgnd scs8hd_fill_2
XFILLER_5_94 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_fill_1
XANTENNA__092__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__283__A _283_/A vgnd vpwr scs8hd_diode_2
X_285_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _179_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_80 vgnd vpwr scs8hd_fill_1
XFILLER_36_124 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__177__B _180_/B vgnd vpwr scs8hd_diode_2
XANTENNA__193__A _130_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_10_28 vgnd vpwr scs8hd_decap_3
XFILLER_27_113 vgnd vpwr scs8hd_fill_1
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_127 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_135 vpwr vgnd scs8hd_fill_2
XANTENNA__278__A _278_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_91 vpwr vgnd scs8hd_fill_2
XFILLER_25_80 vgnd vpwr scs8hd_decap_4
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_268_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_199_ _198_/X _205_/B vgnd vpwr scs8hd_buf_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _203_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__163__D _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__188__A _187_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_62 vgnd vpwr scs8hd_fill_1
XFILLER_2_51 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_171 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A _097_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_122_ _135_/B _123_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _211_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_90 vpwr vgnd scs8hd_fill_2
XANTENNA__174__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _242_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_171 vgnd vpwr scs8hd_decap_3
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _210_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__190__B _188_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vpwr vgnd scs8hd_fill_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_105_ _114_/A _211_/A _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_152 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
XFILLER_7_167 vpwr vgnd scs8hd_fill_2
XFILLER_7_178 vgnd vpwr scs8hd_decap_3
XFILLER_19_263 vpwr vgnd scs8hd_fill_2
XFILLER_19_252 vpwr vgnd scs8hd_fill_2
XANTENNA__185__B _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_61 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _117_/A vgnd vpwr scs8hd_diode_2
XANTENNA__286__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_233 vgnd vpwr scs8hd_fill_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__196__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_247 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _228_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_73 vpwr vgnd scs8hd_fill_2
XFILLER_39_166 vpwr vgnd scs8hd_fill_2
XFILLER_39_111 vgnd vpwr scs8hd_decap_3
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
X_284_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_6_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_210 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XFILLER_5_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_6
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__193__B _188_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _226_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_191 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
X_267_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_198_ _198_/A _198_/X vgnd vpwr scs8hd_buf_1
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
XFILLER_7_19 vpwr vgnd scs8hd_fill_2
X_121_ _120_/X _135_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_21_109 vgnd vpwr scs8hd_fill_1
XANTENNA__174__D _152_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__199__A _198_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_49 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _239_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_60 vgnd vpwr scs8hd_decap_4
XFILLER_7_146 vpwr vgnd scs8hd_fill_2
X_104_ _128_/A _211_/A vgnd vpwr scs8hd_buf_1
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_3
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_267 vgnd vpwr scs8hd_decap_8
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_212 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_259 vpwr vgnd scs8hd_fill_2
XFILLER_16_267 vgnd vpwr scs8hd_decap_8
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_3_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _192_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__196__B _187_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
XFILLER_13_18 vpwr vgnd scs8hd_fill_2
XFILLER_1_108 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_163 vpwr vgnd scs8hd_fill_2
XFILLER_0_152 vgnd vpwr scs8hd_fill_1
XFILLER_0_141 vgnd vpwr scs8hd_decap_4
XFILLER_28_81 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _219_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
X_283_ _283_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_30_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_233 vpwr vgnd scs8hd_fill_2
XFILLER_5_266 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_27_159 vpwr vgnd scs8hd_fill_2
XFILLER_2_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_107 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_192 vgnd vpwr scs8hd_decap_4
XFILLER_26_170 vgnd vpwr scs8hd_decap_6
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
X_266_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _232_/A _152_/B _152_/C _224_/D _198_/A vgnd vpwr scs8hd_or4_4
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _279_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_97 vpwr vgnd scs8hd_fill_2
XFILLER_2_75 vpwr vgnd scs8hd_fill_2
XFILLER_32_151 vpwr vgnd scs8hd_fill_2
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _243_/HI mem_left_track_1.LATCH_7_.latch/Q
+ mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_120_ _152_/A _232_/B _152_/C _208_/D _120_/X vgnd vpwr scs8hd_or4_4
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_249_ _249_/HI _249_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _237_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_243 vgnd vpwr scs8hd_decap_12
XFILLER_28_232 vgnd vpwr scs8hd_decap_8
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_22_83 vpwr vgnd scs8hd_fill_2
XFILLER_22_50 vgnd vpwr scs8hd_fill_1
X_103_ address[1] _103_/B address[0] _128_/A vgnd vpwr scs8hd_or3_4
XFILLER_19_210 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_106 vpwr vgnd scs8hd_fill_2
XFILLER_16_224 vgnd vpwr scs8hd_decap_3
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_271 vgnd vpwr scs8hd_decap_4
XFILLER_13_205 vpwr vgnd scs8hd_fill_2
XFILLER_13_216 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_4
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_29 vpwr vgnd scs8hd_fill_2
XFILLER_24_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_282_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _265_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_72 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_92 vgnd vpwr scs8hd_decap_4
XFILLER_36_116 vgnd vpwr scs8hd_decap_6
XFILLER_36_105 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_265_ _265_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_196_ _149_/A _187_/X _196_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
XFILLER_2_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_270 vpwr vgnd scs8hd_fill_2
XFILLER_2_65 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_163 vpwr vgnd scs8hd_fill_2
XFILLER_23_130 vpwr vgnd scs8hd_fill_2
XFILLER_15_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vpwr vgnd scs8hd_fill_2
XFILLER_14_185 vpwr vgnd scs8hd_fill_2
X_248_ _248_/HI _248_/LO vgnd vpwr scs8hd_conb_1
X_179_ _127_/A _180_/B _179_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_200 vgnd vpwr scs8hd_decap_12
XFILLER_32_18 vpwr vgnd scs8hd_fill_2
XFILLER_28_255 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_144 vgnd vpwr scs8hd_fill_1
X_102_ _114_/A _234_/A _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_115 vgnd vpwr scs8hd_decap_4
XFILLER_11_188 vpwr vgnd scs8hd_fill_2
XFILLER_8_42 vpwr vgnd scs8hd_fill_2
XFILLER_8_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_214 vpwr vgnd scs8hd_fill_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_236 vgnd vpwr scs8hd_fill_1
XFILLER_25_225 vpwr vgnd scs8hd_fill_2
XFILLER_16_236 vgnd vpwr scs8hd_decap_4
XFILLER_17_51 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_94 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__104__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_228 vpwr vgnd scs8hd_fill_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_198 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_254 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _184_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_32 vgnd vpwr scs8hd_decap_3
XFILLER_5_98 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
X_281_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_14_74 vgnd vpwr scs8hd_fill_1
XFILLER_30_84 vgnd vpwr scs8hd_decap_6
XFILLER_39_82 vgnd vpwr scs8hd_decap_3
XFILLER_36_139 vgnd vpwr scs8hd_decap_4
XFILLER_36_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__202__A _234_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_249 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_139 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_264_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_84 vgnd vpwr scs8hd_fill_1
XFILLER_25_62 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ _135_/A _187_/X _195_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _214_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _215_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_247_ _247_/HI _247_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_142 vgnd vpwr scs8hd_fill_1
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _125_/A _180_/B _178_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_37_212 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_41 vgnd vpwr scs8hd_decap_3
X_101_ _101_/A _234_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_11_167 vgnd vpwr scs8hd_decap_4
XFILLER_11_178 vgnd vpwr scs8hd_decap_3
XFILLER_19_256 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_4
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_19_267 vgnd vpwr scs8hd_decap_8
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vgnd vpwr scs8hd_fill_1
XFILLER_8_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_182 vpwr vgnd scs8hd_fill_2
XFILLER_27_19 vpwr vgnd scs8hd_fill_2
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_119 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _192_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__210__A _234_/A vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_73 vpwr vgnd scs8hd_fill_2
XFILLER_33_40 vpwr vgnd scs8hd_fill_2
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
XFILLER_3_130 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _231_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _218_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_251 vpwr vgnd scs8hd_fill_2
XFILLER_12_262 vgnd vpwr scs8hd_decap_12
XFILLER_8_233 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_148 vpwr vgnd scs8hd_fill_2
XFILLER_39_126 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_77 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_181 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _231_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
X_280_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _202_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_203 vgnd vpwr scs8hd_decap_3
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vgnd vpwr scs8hd_decap_4
XFILLER_29_170 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_173 vpwr vgnd scs8hd_fill_2
XANTENNA__202__B _205_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
X_263_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _133_/A _188_/X _194_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XANTENNA__112__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_6
XFILLER_32_143 vgnd vpwr scs8hd_decap_8
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_17_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__213__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_98 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
X_246_ _246_/HI _246_/LO vgnd vpwr scs8hd_conb_1
X_177_ _123_/A _180_/B _177_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_37_224 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_64 vgnd vpwr scs8hd_fill_1
XANTENNA__208__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_102 vpwr vgnd scs8hd_fill_2
X_100_ address[1] _103_/B _106_/C _101_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A address[3] vgnd vpwr scs8hd_diode_2
X_229_ _237_/A _231_/B _229_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _195_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__210__B _211_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_20 vpwr vgnd scs8hd_fill_2
XFILLER_17_31 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_164 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _232_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_260 vpwr vgnd scs8hd_fill_2
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XANTENNA__205__B _205_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _222_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__221__A _237_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _145_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _129_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XFILLER_8_267 vgnd vpwr scs8hd_decap_8
XANTENNA__115__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_39_116 vgnd vpwr scs8hd_decap_6
XFILLER_39_105 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _130_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_30_97 vgnd vpwr scs8hd_fill_1
XFILLER_30_42 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__216__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_237 vgnd vpwr scs8hd_decap_4
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
X_262_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _130_/X _188_/X _193_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XANTENNA__112__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_79 vgnd vpwr scs8hd_decap_3
XFILLER_32_199 vgnd vpwr scs8hd_decap_12
XFILLER_32_188 vgnd vpwr scs8hd_decap_8
XFILLER_17_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__213__B _211_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_11_55 vpwr vgnd scs8hd_fill_2
XFILLER_11_66 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_85 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_8_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_245_ _245_/HI _245_/LO vgnd vpwr scs8hd_conb_1
X_176_ _176_/A _180_/B vgnd vpwr scs8hd_buf_1
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_236 vgnd vpwr scs8hd_decap_8
XFILLER_20_136 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_6_.latch data_in mem_bottom_track_9.LATCH_6_.latch/Q _178_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__208__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_87 vgnd vpwr scs8hd_decap_3
XANTENNA__224__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_19_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_78 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _113_/A vgnd vpwr scs8hd_diode_2
X_228_ _220_/A _231_/B _228_/Y vgnd vpwr scs8hd_nor2_4
X_159_ _130_/X _154_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_3 vgnd vpwr scs8hd_decap_3
XFILLER_25_239 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _202_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _244_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_4
XFILLER_17_65 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_209 vgnd vpwr scs8hd_decap_12
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__219__A _211_/A vgnd vpwr scs8hd_diode_2
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__120__C _152_/C vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_242 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_209 vgnd vpwr scs8hd_decap_4
XANTENNA__221__B _220_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_102 vpwr vgnd scs8hd_fill_2
XFILLER_28_97 vgnd vpwr scs8hd_fill_1
XFILLER_28_64 vgnd vpwr scs8hd_decap_3
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _123_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__216__B _232_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_66 vgnd vpwr scs8hd_decap_6
XFILLER_14_88 vgnd vpwr scs8hd_fill_1
XFILLER_30_76 vgnd vpwr scs8hd_decap_4
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_8
XFILLER_36_109 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_109 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_6_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_219 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_142 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_87 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A _211_/A vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_261_ _261_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
X_192_ _128_/X _188_/X _192_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_58 vgnd vpwr scs8hd_decap_4
XFILLER_2_47 vpwr vgnd scs8hd_fill_2
XFILLER_32_123 vgnd vpwr scs8hd_fill_1
XANTENNA__137__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_134 vgnd vpwr scs8hd_decap_3
XFILLER_23_101 vpwr vgnd scs8hd_fill_2
XFILLER_23_167 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_244_ _244_/HI _244_/LO vgnd vpwr scs8hd_conb_1
XFILLER_36_75 vgnd vpwr scs8hd_decap_8
XFILLER_14_112 vgnd vpwr scs8hd_decap_6
XFILLER_14_145 vgnd vpwr scs8hd_decap_6
XFILLER_14_167 vpwr vgnd scs8hd_fill_2
XFILLER_14_189 vgnd vpwr scs8hd_decap_4
X_175_ _174_/X _176_/A vgnd vpwr scs8hd_buf_1
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_20_148 vgnd vpwr scs8hd_decap_3
XFILLER_20_115 vgnd vpwr scs8hd_decap_8
XFILLER_20_104 vgnd vpwr scs8hd_decap_8
XFILLER_28_226 vgnd vpwr scs8hd_decap_3
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__208__C _232_/C vgnd vpwr scs8hd_diode_2
XANTENNA__224__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_119 vgnd vpwr scs8hd_fill_1
XFILLER_11_148 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_46 vpwr vgnd scs8hd_fill_2
X_227_ _211_/A _231_/B _227_/Y vgnd vpwr scs8hd_nor2_4
X_089_ address[3] _152_/B vgnd vpwr scs8hd_buf_1
X_158_ _128_/X _154_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__150__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__219__B _220_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_229 vgnd vpwr scs8hd_decap_4
XFILLER_17_44 vgnd vpwr scs8hd_decap_4
XFILLER_17_55 vgnd vpwr scs8hd_decap_6
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_32 vpwr vgnd scs8hd_fill_2
XFILLER_33_21 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _211_/A vgnd vpwr scs8hd_diode_2
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_199 vpwr vgnd scs8hd_fill_2
XANTENNA__120__D _208_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_15_273 vgnd vpwr scs8hd_decap_4
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_30_254 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_80 vpwr vgnd scs8hd_fill_2
XFILLER_21_265 vpwr vgnd scs8hd_fill_2
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_87 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _246_/HI mem_right_track_0.LATCH_7_.latch/Q
+ mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _238_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_173 vgnd vpwr scs8hd_decap_8
XANTENNA__216__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_30_55 vgnd vpwr scs8hd_decap_8
XANTENNA__232__B _232_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _247_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_187 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_176 vgnd vpwr scs8hd_fill_1
XFILLER_26_154 vgnd vpwr scs8hd_decap_3
XFILLER_25_44 vpwr vgnd scs8hd_fill_2
XFILLER_25_11 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
X_260_ _260_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XANTENNA__227__B _231_/B vgnd vpwr scs8hd_diode_2
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _127_/A _188_/X _191_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_23_146 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _114_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _173_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_243_ _243_/HI _243_/LO vgnd vpwr scs8hd_conb_1
X_174_ _232_/A _232_/B _152_/C _152_/D _174_/X vgnd vpwr scs8hd_or4_4
XANTENNA__148__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_4
XANTENNA__208__D _208_/D vgnd vpwr scs8hd_diode_2
XFILLER_11_138 vgnd vpwr scs8hd_decap_4
XFILLER_22_67 vgnd vpwr scs8hd_decap_3
XANTENNA__224__C _232_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _127_/A _154_/X _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_160 vpwr vgnd scs8hd_fill_2
X_226_ _234_/A _231_/B _226_/Y vgnd vpwr scs8hd_nor2_4
X_088_ address[4] _152_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_186 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_230 vgnd vpwr scs8hd_decap_4
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_77 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _223_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__235__B _233_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
X_209_ _208_/X _211_/B vgnd vpwr scs8hd_buf_1
XANTENNA__145__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_159 vpwr vgnd scs8hd_fill_2
XFILLER_0_148 vgnd vpwr scs8hd_decap_4
XFILLER_0_137 vpwr vgnd scs8hd_fill_2
XFILLER_5_15 vpwr vgnd scs8hd_fill_2
XFILLER_5_37 vgnd vpwr scs8hd_decap_3
XFILLER_8_204 vgnd vpwr scs8hd_decap_3
XFILLER_8_215 vgnd vpwr scs8hd_decap_4
XFILLER_8_237 vpwr vgnd scs8hd_fill_2
XFILLER_12_255 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _205_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vpwr vgnd scs8hd_fill_2
XANTENNA__156__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_270 vgnd vpwr scs8hd_decap_6
XFILLER_30_23 vgnd vpwr scs8hd_decap_4
XFILLER_30_12 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _245_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_229 vpwr vgnd scs8hd_fill_2
XANTENNA__216__D _152_/D vgnd vpwr scs8hd_diode_2
XANTENNA__232__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_262 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_177 vgnd vpwr scs8hd_decap_6
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_188 vpwr vgnd scs8hd_fill_2
XFILLER_26_166 vpwr vgnd scs8hd_fill_2
XFILLER_25_67 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_190_ _125_/A _188_/X _190_/Y vgnd vpwr scs8hd_nor2_4
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_254 vpwr vgnd scs8hd_fill_2
XFILLER_17_177 vpwr vgnd scs8hd_fill_2
XFILLER_17_133 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_31_191 vgnd vpwr scs8hd_decap_4
XFILLER_11_14 vpwr vgnd scs8hd_fill_2
XANTENNA__238__B _233_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
XANTENNA__254__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
X_242_ _242_/HI _242_/LO vgnd vpwr scs8hd_conb_1
X_173_ _149_/A _164_/X _173_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_3
XFILLER_13_191 vpwr vgnd scs8hd_fill_2
XFILLER_22_46 vpwr vgnd scs8hd_fill_2
XFILLER_11_106 vgnd vpwr scs8hd_decap_3
XFILLER_22_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XANTENNA__224__D _224_/D vgnd vpwr scs8hd_diode_2
XFILLER_19_206 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_087_ _200_/A _123_/A vgnd vpwr scs8hd_buf_1
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_132 vpwr vgnd scs8hd_fill_2
XFILLER_6_165 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_225_ _224_/X _231_/B vgnd vpwr scs8hd_buf_1
X_156_ _125_/A _154_/X _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_272 vgnd vpwr scs8hd_decap_3
XANTENNA__159__A _130_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_30_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_139_ _232_/A _232_/B _152_/C _208_/D _139_/X vgnd vpwr scs8hd_or4_4
X_208_ _232_/A _152_/B _232_/C _208_/D _208_/X vgnd vpwr scs8hd_or4_4
XANTENNA__161__B _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_212 vgnd vpwr scs8hd_decap_3
XFILLER_21_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_45 vpwr vgnd scs8hd_fill_2
XFILLER_28_23 vgnd vpwr scs8hd_decap_4
XFILLER_28_12 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_201 vpwr vgnd scs8hd_fill_2
XFILLER_12_234 vpwr vgnd scs8hd_fill_2
XANTENNA__262__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_5_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_260 vpwr vgnd scs8hd_fill_2
XANTENNA__156__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_36 vpwr vgnd scs8hd_fill_2
XFILLER_30_35 vgnd vpwr scs8hd_decap_4
XANTENNA__082__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_99 vgnd vpwr scs8hd_decap_4
XFILLER_39_88 vpwr vgnd scs8hd_fill_2
XFILLER_39_11 vgnd vpwr scs8hd_decap_12
XANTENNA__232__D _224_/D vgnd vpwr scs8hd_diode_2
XANTENNA__257__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_197 vpwr vgnd scs8hd_fill_2
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_252 vgnd vpwr scs8hd_fill_1
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_35_156 vpwr vgnd scs8hd_fill_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _125_/A vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_200 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_266 vpwr vgnd scs8hd_fill_2
XFILLER_32_126 vpwr vgnd scs8hd_fill_2
XFILLER_32_115 vgnd vpwr scs8hd_decap_8
XFILLER_32_104 vgnd vpwr scs8hd_decap_8
XFILLER_17_189 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_fill_1
XFILLER_17_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _226_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_181 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
XFILLER_11_37 vgnd vpwr scs8hd_decap_3
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _183_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_241_ _241_/HI _241_/LO vgnd vpwr scs8hd_conb_1
X_172_ _135_/A _164_/X _172_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__270__A _270_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_130 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_218 vgnd vpwr scs8hd_decap_8
XFILLER_3_71 vpwr vgnd scs8hd_fill_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _207_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_229 vpwr vgnd scs8hd_fill_2
XANTENNA__265__A _265_/A vgnd vpwr scs8hd_diode_2
X_224_ _152_/A _152_/B _232_/C _224_/D _224_/X vgnd vpwr scs8hd_or4_4
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
X_155_ _123_/A _154_/X _155_/Y vgnd vpwr scs8hd_nor2_4
X_086_ _085_/X _200_/A vgnd vpwr scs8hd_buf_1
XANTENNA__159__B _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _174_/X vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_13 vgnd vpwr scs8hd_decap_4
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_69 vpwr vgnd scs8hd_fill_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_103 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vgnd vpwr scs8hd_decap_3
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _214_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_90 vgnd vpwr scs8hd_decap_4
XFILLER_15_254 vgnd vpwr scs8hd_decap_4
XFILLER_15_265 vpwr vgnd scs8hd_fill_2
X_207_ _239_/A _198_/X _207_/Y vgnd vpwr scs8hd_nor2_4
X_138_ address[4] _232_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_106 vgnd vpwr scs8hd_fill_1
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_1.LATCH_6_.latch data_in mem_bottom_track_1.LATCH_6_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vpwr vgnd scs8hd_fill_2
XFILLER_38_132 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_23 vgnd vpwr scs8hd_decap_12
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__273__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _191_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_135 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__183__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB _190_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _287_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_146 vgnd vpwr scs8hd_decap_4
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XFILLER_25_25 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _152_/A vgnd vpwr scs8hd_diode_2
XANTENNA__268__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA__088__A address[4] vgnd vpwr scs8hd_diode_2
X_240_ _240_/HI _240_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_138 vgnd vpwr scs8hd_decap_4
XFILLER_22_171 vgnd vpwr scs8hd_decap_3
X_171_ _133_/A _165_/X _171_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _230_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vgnd vpwr scs8hd_decap_4
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XANTENNA__180__B _180_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_208 vgnd vpwr scs8hd_decap_6
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_230 vpwr vgnd scs8hd_fill_2
X_223_ _239_/A _220_/B _223_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__281__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
X_154_ _153_/X _154_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_196 vpwr vgnd scs8hd_fill_2
XFILLER_12_81 vpwr vgnd scs8hd_fill_2
X_085_ _106_/A _103_/B _106_/C _085_/X vgnd vpwr scs8hd_or3_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_230 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_200 vpwr vgnd scs8hd_fill_2
XFILLER_17_48 vgnd vpwr scs8hd_fill_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_36 vpwr vgnd scs8hd_fill_2
XFILLER_33_25 vgnd vpwr scs8hd_decap_4
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _103_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_148 vpwr vgnd scs8hd_fill_2
XFILLER_3_126 vpwr vgnd scs8hd_fill_2
XANTENNA__276__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _162_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_137_ _149_/A _135_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_206_ _114_/B _198_/X _206_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_21_258 vgnd vpwr scs8hd_decap_4
XANTENNA__186__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _252_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _235_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_69 vgnd vpwr scs8hd_decap_3
XANTENNA__096__A _117_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_6_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_38_188 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_14_49 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_35 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _251_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_232 vgnd vpwr scs8hd_fill_1
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_169 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _256_/A vgnd vpwr scs8hd_inv_1
XANTENNA__183__B _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_48 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_169 vpwr vgnd scs8hd_fill_2
XFILLER_17_103 vpwr vgnd scs8hd_fill_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XANTENNA__284__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_139 vpwr vgnd scs8hd_fill_2
XFILLER_15_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__178__B _180_/B vgnd vpwr scs8hd_diode_2
XANTENNA__194__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_191 vpwr vgnd scs8hd_fill_2
XFILLER_31_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_58 vgnd vpwr scs8hd_decap_8
XFILLER_36_47 vgnd vpwr scs8hd_decap_8
XFILLER_22_150 vgnd vpwr scs8hd_fill_1
X_170_ _130_/X _165_/X _170_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__279__A _279_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_80 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_51 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _114_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
XFILLER_27_242 vpwr vgnd scs8hd_fill_2
X_153_ _152_/X _153_/X vgnd vpwr scs8hd_buf_1
X_222_ _114_/B _220_/B _222_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_113 vgnd vpwr scs8hd_decap_6
XFILLER_10_131 vgnd vpwr scs8hd_decap_3
XFILLER_10_164 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _248_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_9 vpwr vgnd scs8hd_fill_2
X_084_ address[0] _106_/C vgnd vpwr scs8hd_inv_8
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__191__B _188_/X vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XFILLER_17_16 vpwr vgnd scs8hd_fill_2
XFILLER_17_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _247_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__085__C _106_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_223 vpwr vgnd scs8hd_fill_2
XFILLER_30_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_205_ _237_/A _205_/B _205_/Y vgnd vpwr scs8hd_nor2_4
X_136_ _116_/A _149_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_182 vpwr vgnd scs8hd_fill_2
XANTENNA__186__B _232_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XFILLER_5_19 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_7_.latch data_in mem_bottom_track_9.LATCH_7_.latch/Q _177_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_219 vgnd vpwr scs8hd_fill_1
XANTENNA__287__A _287_/A vgnd vpwr scs8hd_diode_2
X_119_ _091_/A _152_/C vgnd vpwr scs8hd_buf_1
XFILLER_38_167 vgnd vpwr scs8hd_decap_3
XANTENNA__197__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_47 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_156 vgnd vpwr scs8hd_decap_3
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_6_.latch data_in mem_left_track_9.LATCH_6_.latch/Q _201_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_80 vgnd vpwr scs8hd_fill_1
XFILLER_20_71 vpwr vgnd scs8hd_fill_2
XFILLER_35_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C _232_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_258 vpwr vgnd scs8hd_fill_2
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_137 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XANTENNA__194__B _188_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_18 vpwr vgnd scs8hd_fill_2
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_3
XFILLER_9_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_166 vpwr vgnd scs8hd_fill_2
XFILLER_9_199 vpwr vgnd scs8hd_fill_2
XFILLER_13_195 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__B _188_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__099__B _099_/B vgnd vpwr scs8hd_diode_2
X_221_ _237_/A _220_/B _221_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_154 vgnd vpwr scs8hd_decap_3
X_152_ _152_/A _152_/B _152_/C _152_/D _152_/X vgnd vpwr scs8hd_or4_4
X_083_ address[2] _103_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_37_80 vgnd vpwr scs8hd_fill_1
XFILLER_33_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_243 vpwr vgnd scs8hd_fill_2
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _212_/Y vgnd vpwr scs8hd_diode_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_204_ _220_/A _205_/B _204_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _135_/A _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__186__C _152_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_238 vgnd vpwr scs8hd_decap_4
XFILLER_28_49 vgnd vpwr scs8hd_decap_4
XFILLER_8_209 vgnd vpwr scs8hd_decap_4
XFILLER_12_205 vgnd vpwr scs8hd_decap_8
XFILLER_12_238 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_118_ address[3] _232_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_124 vgnd vpwr scs8hd_decap_8
XFILLER_38_113 vgnd vpwr scs8hd_decap_8
XFILLER_38_102 vgnd vpwr scs8hd_decap_6
XANTENNA__197__B _152_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _242_/HI mem_bottom_track_9.LATCH_7_.latch/Q
+ mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_39 vgnd vpwr scs8hd_fill_1
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_245 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _229_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__093__D _208_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_6_.latch data_in mem_right_track_8.LATCH_6_.latch/Q _156_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_14_108 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _237_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB _200_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_60 vpwr vgnd scs8hd_fill_2
XFILLER_9_112 vpwr vgnd scs8hd_fill_2
XFILLER_9_145 vpwr vgnd scs8hd_fill_2
XFILLER_9_189 vgnd vpwr scs8hd_fill_1
XFILLER_3_86 vpwr vgnd scs8hd_fill_2
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
X_220_ _220_/A _220_/B _220_/Y vgnd vpwr scs8hd_nor2_4
X_151_ address[5] _150_/Y _152_/D vgnd vpwr scs8hd_nand2_4
X_082_ address[1] _106_/A vgnd vpwr scs8hd_inv_8
XFILLER_12_62 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _250_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_214 vgnd vpwr scs8hd_decap_12
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_17 vgnd vpwr scs8hd_fill_1
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_107 vpwr vgnd scs8hd_fill_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_203 vgnd vpwr scs8hd_decap_4
X_203_ _211_/A _205_/B _203_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_269 vpwr vgnd scs8hd_fill_2
XFILLER_23_94 vgnd vpwr scs8hd_fill_1
X_134_ _113_/A _135_/A vgnd vpwr scs8hd_buf_1
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_195 vpwr vgnd scs8hd_fill_2
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_217 vgnd vpwr scs8hd_decap_3
XANTENNA__186__D _224_/D vgnd vpwr scs8hd_diode_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_72 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_4
X_117_ _117_/A _239_/A _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_254 vgnd vpwr scs8hd_decap_4
XFILLER_11_261 vgnd vpwr scs8hd_fill_1
XFILLER_7_276 vgnd vpwr scs8hd_fill_1
XANTENNA__197__C _152_/C vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _196_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_30_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _193_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_20_51 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_235 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_139 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _222_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_75 vpwr vgnd scs8hd_fill_2
XFILLER_6_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_106 vpwr vgnd scs8hd_fill_2
XFILLER_25_29 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_205 vgnd vpwr scs8hd_decap_3
XFILLER_9_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _220_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_83 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_150 vgnd vpwr scs8hd_fill_1
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_120 vpwr vgnd scs8hd_fill_2
XFILLER_13_142 vgnd vpwr scs8hd_decap_6
XFILLER_13_175 vgnd vpwr scs8hd_fill_1
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_21 vpwr vgnd scs8hd_fill_2
XFILLER_22_19 vgnd vpwr scs8hd_fill_1
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
XFILLER_27_234 vgnd vpwr scs8hd_decap_6
XFILLER_10_123 vpwr vgnd scs8hd_fill_2
X_150_ address[6] _150_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_149 vgnd vpwr scs8hd_decap_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_41 vpwr vgnd scs8hd_fill_2
XFILLER_12_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_226 vgnd vpwr scs8hd_decap_12
X_279_ _279_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_248 vgnd vpwr scs8hd_decap_8
XFILLER_24_237 vgnd vpwr scs8hd_decap_8
XFILLER_24_226 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _238_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_218 vgnd vpwr scs8hd_decap_12
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
X_202_ _234_/A _205_/B _202_/Y vgnd vpwr scs8hd_nor2_4
X_133_ _133_/A _123_/B _133_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_163 vgnd vpwr scs8hd_decap_3
XANTENNA__110__A _132_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_229 vgnd vpwr scs8hd_decap_3
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_3
XFILLER_28_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_50 vgnd vpwr scs8hd_decap_6
XFILLER_18_84 vgnd vpwr scs8hd_decap_8
XANTENNA__105__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_200 vgnd vpwr scs8hd_fill_1
XFILLER_7_233 vgnd vpwr scs8hd_decap_4
XFILLER_7_266 vpwr vgnd scs8hd_fill_2
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
X_116_ _116_/A _239_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_159 vgnd vpwr scs8hd_decap_8
XANTENNA__197__D _224_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_83 vgnd vpwr scs8hd_decap_3
XFILLER_6_10 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_3
XFILLER_6_54 vpwr vgnd scs8hd_fill_2
XFILLER_34_173 vgnd vpwr scs8hd_decap_4
XFILLER_26_129 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _137_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_107 vpwr vgnd scs8hd_fill_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_176 vgnd vpwr scs8hd_decap_8
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_85 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vpwr vgnd scs8hd_fill_2
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
XANTENNA__102__B _234_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_173 vgnd vpwr scs8hd_decap_3
XFILLER_31_198 vpwr vgnd scs8hd_fill_2
XFILLER_31_187 vpwr vgnd scs8hd_fill_2
XFILLER_31_176 vgnd vpwr scs8hd_decap_3
XFILLER_31_165 vpwr vgnd scs8hd_fill_2
XFILLER_31_143 vgnd vpwr scs8hd_decap_4
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_195 vpwr vgnd scs8hd_fill_2
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_176 vpwr vgnd scs8hd_fill_2
XFILLER_22_187 vgnd vpwr scs8hd_decap_8
XANTENNA__203__A _211_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_154 vpwr vgnd scs8hd_fill_2
XFILLER_13_187 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_55 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _269_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_3
XFILLER_6_128 vpwr vgnd scs8hd_fill_2
XFILLER_10_179 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_83 vgnd vpwr scs8hd_decap_3
XFILLER_33_238 vgnd vpwr scs8hd_decap_6
XANTENNA__108__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
X_278_ _278_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_150 vgnd vpwr scs8hd_decap_4
XANTENNA__200__B _205_/B vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_201_ _099_/B _205_/B _201_/Y vgnd vpwr scs8hd_nor2_4
X_132_ _132_/A _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_131 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _182_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _261_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_219 vpwr vgnd scs8hd_fill_2
XANTENNA__211__A _211_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_84 vpwr vgnd scs8hd_fill_2
XFILLER_34_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__105__B _211_/A vgnd vpwr scs8hd_diode_2
X_115_ address[1] address[2] address[0] _116_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__121__A _120_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _206_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_138 vgnd vpwr scs8hd_decap_12
XFILLER_29_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vpwr vgnd scs8hd_fill_2
XANTENNA__206__A _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_119 vgnd vpwr scs8hd_fill_1
XFILLER_28_160 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _213_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_119 vgnd vpwr scs8hd_decap_8
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_1_229 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_188 vgnd vpwr scs8hd_decap_12
XFILLER_40_166 vgnd vpwr scs8hd_decap_6
XFILLER_15_42 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_1.LATCH_7_.latch data_in mem_bottom_track_1.LATCH_7_.latch/Q _166_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
.ends

