VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_right
  CLASS BLOCK ;
  FOREIGN grid_io_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 1665.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 47.600 83.000 50.000 83.600 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 1662.600 3.130 1665.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 1662.600 9.110 1665.000 ;
    END
  END address[3]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 47.600 248.920 50.000 249.520 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 1662.600 15.550 1665.000 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 47.600 415.520 50.000 416.120 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 2.400 356.280 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 47.600 582.120 50.000 582.720 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 47.600 748.720 50.000 749.320 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 1662.600 21.530 1665.000 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 47.600 1415.120 50.000 1415.720 ;
    END
  END left_width_0_height_0__pin_10_
  PIN left_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END left_width_0_height_0__pin_11_
  PIN left_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.680 2.400 1070.280 ;
    END
  END left_width_0_height_0__pin_12_
  PIN left_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 47.600 1581.720 50.000 1582.320 ;
    END
  END left_width_0_height_0__pin_13_
  PIN left_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.680 2.400 1308.280 ;
    END
  END left_width_0_height_0__pin_14_
  PIN left_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1545.680 2.400 1546.280 ;
    END
  END left_width_0_height_0__pin_15_
  PIN left_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 47.600 915.320 50.000 915.920 ;
    END
  END left_width_0_height_0__pin_1_
  PIN left_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 2.400 594.280 ;
    END
  END left_width_0_height_0__pin_2_
  PIN left_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 47.600 1081.920 50.000 1082.520 ;
    END
  END left_width_0_height_0__pin_3_
  PIN left_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 1662.600 27.970 1665.000 ;
    END
  END left_width_0_height_0__pin_4_
  PIN left_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 47.600 1248.520 50.000 1249.120 ;
    END
  END left_width_0_height_0__pin_5_
  PIN left_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 1662.600 34.410 1665.000 ;
    END
  END left_width_0_height_0__pin_6_
  PIN left_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.110 1662.600 40.390 1665.000 ;
    END
  END left_width_0_height_0__pin_7_
  PIN left_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 1662.600 46.830 1665.000 ;
    END
  END left_width_0_height_0__pin_8_
  PIN left_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.680 2.400 832.280 ;
    END
  END left_width_0_height_0__pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 13.055 10.640 14.655 1654.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 21.385 10.640 22.985 1654.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 44.160 1653.845 ;
      LAYER met1 ;
        RECT 0.070 0.380 46.850 1662.900 ;
      LAYER met2 ;
        RECT 0.090 1662.320 2.570 1663.010 ;
        RECT 3.410 1662.320 8.550 1663.010 ;
        RECT 9.390 1662.320 14.990 1663.010 ;
        RECT 15.830 1662.320 20.970 1663.010 ;
        RECT 21.810 1662.320 27.410 1663.010 ;
        RECT 28.250 1662.320 33.850 1663.010 ;
        RECT 34.690 1662.320 39.830 1663.010 ;
        RECT 40.670 1662.320 46.270 1663.010 ;
        RECT 0.090 2.680 46.760 1662.320 ;
        RECT 0.090 0.270 4.410 2.680 ;
        RECT 5.250 0.270 14.070 2.680 ;
        RECT 14.910 0.270 24.190 2.680 ;
        RECT 25.030 0.270 34.310 2.680 ;
        RECT 35.150 0.270 44.430 2.680 ;
        RECT 45.270 0.270 46.760 2.680 ;
      LAYER met3 ;
        RECT 0.310 1582.720 48.450 1653.925 ;
        RECT 0.310 1581.320 47.200 1582.720 ;
        RECT 0.310 1546.680 48.450 1581.320 ;
        RECT 2.800 1545.280 48.450 1546.680 ;
        RECT 0.310 1416.120 48.450 1545.280 ;
        RECT 0.310 1414.720 47.200 1416.120 ;
        RECT 0.310 1308.680 48.450 1414.720 ;
        RECT 2.800 1307.280 48.450 1308.680 ;
        RECT 0.310 1249.520 48.450 1307.280 ;
        RECT 0.310 1248.120 47.200 1249.520 ;
        RECT 0.310 1082.920 48.450 1248.120 ;
        RECT 0.310 1081.520 47.200 1082.920 ;
        RECT 0.310 1070.680 48.450 1081.520 ;
        RECT 2.800 1069.280 48.450 1070.680 ;
        RECT 0.310 916.320 48.450 1069.280 ;
        RECT 0.310 914.920 47.200 916.320 ;
        RECT 0.310 832.680 48.450 914.920 ;
        RECT 2.800 831.280 48.450 832.680 ;
        RECT 0.310 749.720 48.450 831.280 ;
        RECT 0.310 748.320 47.200 749.720 ;
        RECT 0.310 594.680 48.450 748.320 ;
        RECT 2.800 593.280 48.450 594.680 ;
        RECT 0.310 583.120 48.450 593.280 ;
        RECT 0.310 581.720 47.200 583.120 ;
        RECT 0.310 416.520 48.450 581.720 ;
        RECT 0.310 415.120 47.200 416.520 ;
        RECT 0.310 356.680 48.450 415.120 ;
        RECT 2.800 355.280 48.450 356.680 ;
        RECT 0.310 249.920 48.450 355.280 ;
        RECT 0.310 248.520 47.200 249.920 ;
        RECT 0.310 119.360 48.450 248.520 ;
        RECT 2.800 117.960 48.450 119.360 ;
        RECT 0.310 84.000 48.450 117.960 ;
        RECT 0.310 82.600 47.200 84.000 ;
        RECT 0.310 10.715 48.450 82.600 ;
      LAYER met4 ;
        RECT 15.055 10.640 20.985 1654.000 ;
        RECT 23.385 10.640 39.650 1654.000 ;
  END
END grid_io_right
END LIBRARY

