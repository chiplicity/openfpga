* NGSPICE file created from sb_0__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_0__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_11_
+ top_left_grid_pin_13_ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_
+ top_left_grid_pin_5_ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_
+ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_211 vgnd vpwr scs8hd_decap_4
XFILLER_39_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_188 vpwr vgnd scs8hd_fill_2
XFILLER_36_247 vpwr vgnd scs8hd_fill_2
XFILLER_36_258 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_192 vgnd vpwr scs8hd_decap_4
XFILLER_27_258 vgnd vpwr scs8hd_decap_4
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_158 vgnd vpwr scs8hd_fill_1
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _202_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_84 vgnd vpwr scs8hd_fill_1
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XFILLER_33_228 vgnd vpwr scs8hd_decap_3
XANTENNA__124__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_239 vpwr vgnd scs8hd_fill_2
XFILLER_15_217 vpwr vgnd scs8hd_fill_2
X_131_ _129_/X _130_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__110__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_97 vgnd vpwr scs8hd_fill_1
X_114_ _163_/B _114_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_235 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _206_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _172_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_6
XFILLER_35_109 vpwr vgnd scs8hd_fill_2
XFILLER_28_150 vgnd vpwr scs8hd_decap_3
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_120 vgnd vpwr scs8hd_decap_6
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_40_101 vgnd vpwr scs8hd_fill_1
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_156 vpwr vgnd scs8hd_fill_2
XFILLER_31_167 vgnd vpwr scs8hd_decap_4
XFILLER_31_123 vpwr vgnd scs8hd_fill_2
XFILLER_16_120 vgnd vpwr scs8hd_decap_3
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_22_101 vgnd vpwr scs8hd_decap_6
Xmem_top_track_4.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_8
XFILLER_36_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_171 vgnd vpwr scs8hd_decap_6
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_4
XFILLER_37_96 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_41_262 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_32_240 vgnd vpwr scs8hd_fill_1
XFILLER_24_229 vgnd vpwr scs8hd_decap_3
XFILLER_24_207 vgnd vpwr scs8hd_decap_6
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_130_ _126_/A _114_/X _134_/C _169_/A _130_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
XANTENNA__110__D _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_240 vgnd vpwr scs8hd_decap_8
XANTENNA__135__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_243 vpwr vgnd scs8hd_fill_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
X_113_ address[2] _163_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_221 vpwr vgnd scs8hd_fill_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_28_184 vpwr vgnd scs8hd_fill_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_124 vgnd vpwr scs8hd_decap_3
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_135 vgnd vpwr scs8hd_fill_1
XFILLER_16_143 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vgnd vpwr scs8hd_decap_3
XFILLER_22_168 vgnd vpwr scs8hd_decap_4
XFILLER_22_146 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_146 vpwr vgnd scs8hd_fill_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_161 vgnd vpwr scs8hd_fill_1
XFILLER_27_227 vgnd vpwr scs8hd_fill_1
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_41_274 vgnd vpwr scs8hd_decap_3
XFILLER_41_241 vgnd vpwr scs8hd_decap_3
XANTENNA__140__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__135__B _134_/X vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
X_112_ _125_/A _112_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_29_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_130 vpwr vgnd scs8hd_fill_2
XFILLER_37_152 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _192_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_163 vpwr vgnd scs8hd_fill_2
XFILLER_19_163 vgnd vpwr scs8hd_fill_1
XFILLER_25_133 vpwr vgnd scs8hd_fill_2
XFILLER_31_99 vgnd vpwr scs8hd_decap_4
XFILLER_16_133 vgnd vpwr scs8hd_fill_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_147 vgnd vpwr scs8hd_decap_3
XFILLER_31_114 vgnd vpwr scs8hd_decap_8
XFILLER_16_199 vgnd vpwr scs8hd_decap_4
XANTENNA__143__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _196_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_206 vpwr vgnd scs8hd_fill_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_206 vpwr vgnd scs8hd_fill_2
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_261 vgnd vpwr scs8hd_decap_12
XFILLER_26_250 vpwr vgnd scs8hd_fill_2
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_253 vpwr vgnd scs8hd_fill_2
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__C _153_/C vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_264 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _200_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__151__B _151_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ _119_/A _112_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B _114_/X vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
XFILLER_37_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_142 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _204_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_123 vgnd vpwr scs8hd_fill_1
XFILLER_25_156 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_259 vgnd vpwr scs8hd_decap_3
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_159 vpwr vgnd scs8hd_fill_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_270 vgnd vpwr scs8hd_decap_6
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _156_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_196 vgnd vpwr scs8hd_fill_1
XFILLER_8_141 vgnd vpwr scs8hd_decap_8
XANTENNA__170__A _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_26_273 vpwr vgnd scs8hd_fill_2
XANTENNA__140__D _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_188 vgnd vpwr scs8hd_decap_12
XANTENNA__149__B _114_/X vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_243 vgnd vpwr scs8hd_decap_3
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_221 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _123_/B _123_/C _170_/A _112_/B vgnd vpwr scs8hd_or4_4
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
X_239_ _239_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _153_/C vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_121 vgnd vpwr scs8hd_decap_4
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_40_116 vgnd vpwr scs8hd_decap_8
XFILLER_40_105 vgnd vpwr scs8hd_decap_8
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_127 vpwr vgnd scs8hd_fill_2
XFILLER_24_190 vpwr vgnd scs8hd_fill_2
XFILLER_16_168 vgnd vpwr scs8hd_decap_4
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_21_90 vpwr vgnd scs8hd_fill_2
XANTENNA__168__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_227 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_230 vgnd vpwr scs8hd_decap_3
XFILLER_18_219 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_266 vgnd vpwr scs8hd_decap_8
Xmem_top_track_8.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_32_222 vgnd vpwr scs8hd_decap_3
XFILLER_17_263 vpwr vgnd scs8hd_fill_2
XFILLER_17_252 vpwr vgnd scs8hd_fill_2
XFILLER_17_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _164_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_255 vgnd vpwr scs8hd_decap_3
XFILLER_32_266 vgnd vpwr scs8hd_decap_8
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_200 vpwr vgnd scs8hd_fill_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_4
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vpwr vgnd scs8hd_fill_2
XFILLER_11_258 vpwr vgnd scs8hd_fill_2
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_225 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_169_ _169_/A _170_/B _165_/A _169_/Y vgnd vpwr scs8hd_nor3_4
X_238_ _238_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__D _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_188 vgnd vpwr scs8hd_decap_4
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_19_155 vpwr vgnd scs8hd_fill_2
XFILLER_19_111 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__157__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_169 vgnd vpwr scs8hd_decap_4
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_25_114 vgnd vpwr scs8hd_decap_6
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_180 vgnd vpwr scs8hd_decap_4
XFILLER_16_147 vgnd vpwr scs8hd_decap_4
XFILLER_16_125 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _190_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_217 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_117 vgnd vpwr scs8hd_decap_8
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_14.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_194 vgnd vpwr scs8hd_decap_3
XFILLER_12_161 vgnd vpwr scs8hd_decap_12
XFILLER_8_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__170__C _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_8
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XANTENNA__149__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _194_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_4
XFILLER_23_201 vgnd vpwr scs8hd_fill_1
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_14_223 vgnd vpwr scs8hd_decap_3
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_226 vgnd vpwr scs8hd_decap_8
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
X_168_ _169_/A _170_/B _164_/A _168_/Y vgnd vpwr scs8hd_nor3_4
X_237_ _237_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
XFILLER_10_270 vgnd vpwr scs8hd_decap_4
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XFILLER_6_252 vgnd vpwr scs8hd_decap_3
X_099_ address[4] address[5] _134_/C vgnd vpwr scs8hd_or2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_134 vgnd vpwr scs8hd_decap_3
XFILLER_37_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_145 vgnd vpwr scs8hd_decap_3
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_167 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_104 vpwr vgnd scs8hd_fill_2
XFILLER_34_137 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_4
XANTENNA__157__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_181 vpwr vgnd scs8hd_fill_2
XFILLER_25_137 vpwr vgnd scs8hd_fill_2
XFILLER_25_104 vgnd vpwr scs8hd_decap_8
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_129 vpwr vgnd scs8hd_fill_2
XFILLER_22_107 vgnd vpwr scs8hd_fill_1
XFILLER_30_184 vpwr vgnd scs8hd_fill_2
XFILLER_30_140 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XFILLER_38_273 vpwr vgnd scs8hd_fill_2
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_162 vpwr vgnd scs8hd_fill_2
XFILLER_21_151 vpwr vgnd scs8hd_fill_2
XFILLER_13_129 vpwr vgnd scs8hd_fill_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _202_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_173 vpwr vgnd scs8hd_fill_2
XFILLER_12_140 vgnd vpwr scs8hd_decap_8
XFILLER_8_188 vpwr vgnd scs8hd_fill_2
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_254 vpwr vgnd scs8hd_fill_2
XFILLER_35_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_254 vgnd vpwr scs8hd_decap_4
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_27_91 vpwr vgnd scs8hd_fill_2
XFILLER_23_213 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XFILLER_14_257 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_205 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_098_ address[2] _123_/B vgnd vpwr scs8hd_buf_1
X_167_ _166_/X _170_/B vgnd vpwr scs8hd_buf_1
X_236_ _236_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_37_113 vpwr vgnd scs8hd_fill_2
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_163 vpwr vgnd scs8hd_fill_2
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_130 vpwr vgnd scs8hd_fill_2
XFILLER_29_230 vgnd vpwr scs8hd_decap_3
XFILLER_16_93 vgnd vpwr scs8hd_decap_6
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
Xmem_top_track_10.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_236 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_8
XFILLER_9_273 vgnd vpwr scs8hd_decap_4
XFILLER_9_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_235_ _235_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
X_097_ address[3] _110_/A vgnd vpwr scs8hd_buf_1
X_166_ address[3] address[2] address[4] _137_/Y _166_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_125 vgnd vpwr scs8hd_fill_1
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
X_149_ address[3] _114_/X _153_/C _163_/D _151_/B vgnd vpwr scs8hd_or4_4
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_161 vpwr vgnd scs8hd_fill_2
XFILLER_24_150 vgnd vpwr scs8hd_fill_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_186 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_267 vgnd vpwr scs8hd_decap_8
XFILLER_17_223 vgnd vpwr scs8hd_fill_1
XFILLER_32_215 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_204 vgnd vpwr scs8hd_decap_4
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_215 vgnd vpwr scs8hd_decap_4
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_38_81 vgnd vpwr scs8hd_decap_8
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_241 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _192_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
X_165_ _165_/A _164_/B _165_/Y vgnd vpwr scs8hd_nor2_4
X_234_ _234_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
X_096_ _096_/A _119_/A vgnd vpwr scs8hd_buf_1
XFILLER_40_93 vgnd vpwr scs8hd_decap_8
XFILLER_40_60 vgnd vpwr scs8hd_decap_12
XFILLER_37_126 vpwr vgnd scs8hd_fill_2
XFILLER_37_148 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_104 vgnd vpwr scs8hd_decap_8
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_4
XFILLER_19_115 vgnd vpwr scs8hd_fill_1
XFILLER_19_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_60 vgnd vpwr scs8hd_fill_1
X_148_ _151_/A _147_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_192 vgnd vpwr scs8hd_decap_3
XFILLER_33_173 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_6
XFILLER_33_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XFILLER_15_162 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_38_254 vgnd vpwr scs8hd_decap_8
XFILLER_38_265 vgnd vpwr scs8hd_decap_8
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_21_143 vpwr vgnd scs8hd_fill_2
XFILLER_29_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
XFILLER_29_221 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_158 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_235 vgnd vpwr scs8hd_decap_6
XFILLER_26_224 vgnd vpwr scs8hd_decap_4
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XFILLER_41_205 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _200_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_260 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
Xmem_right_track_14.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_220 vpwr vgnd scs8hd_fill_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_095_ address[0] _096_/A vgnd vpwr scs8hd_inv_8
X_164_ _164_/A _164_/B _164_/Y vgnd vpwr scs8hd_nor2_4
X_233_ _233_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_40_72 vgnd vpwr scs8hd_decap_12
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
XANTENNA__111__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_108 vgnd vpwr scs8hd_decap_12
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_35_94 vpwr vgnd scs8hd_fill_2
X_147_ _129_/X _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XFILLER_18_171 vpwr vgnd scs8hd_fill_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_16_108 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _188_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_188 vgnd vpwr scs8hd_decap_4
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_266 vpwr vgnd scs8hd_fill_2
XFILLER_35_214 vgnd vpwr scs8hd_decap_8
XFILLER_35_258 vgnd vpwr scs8hd_decap_4
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_217 vgnd vpwr scs8hd_decap_12
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_203 vgnd vpwr scs8hd_fill_1
XFILLER_32_206 vgnd vpwr scs8hd_decap_8
XFILLER_27_95 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_236 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_31_272 vgnd vpwr scs8hd_decap_4
XFILLER_23_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_228 vgnd vpwr scs8hd_decap_3
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_13_250 vgnd vpwr scs8hd_decap_4
XFILLER_9_210 vgnd vpwr scs8hd_decap_8
X_232_ _232_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_163_ _163_/A _163_/B _163_/C _163_/D _164_/B vgnd vpwr scs8hd_or4_4
XFILLER_40_84 vgnd vpwr scs8hd_decap_8
XFILLER_24_96 vpwr vgnd scs8hd_fill_2
XFILLER_6_246 vgnd vpwr scs8hd_decap_4
XANTENNA__111__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_128 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_150 vgnd vpwr scs8hd_decap_3
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_146_ address[3] _114_/X _153_/C _153_/D _147_/B vgnd vpwr scs8hd_or4_4
XANTENNA__122__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_186 vpwr vgnd scs8hd_fill_2
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
XFILLER_21_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_167 vgnd vpwr scs8hd_decap_12
XFILLER_15_197 vgnd vpwr scs8hd_decap_4
X_129_ _096_/A _129_/X vgnd vpwr scs8hd_buf_1
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vgnd vpwr scs8hd_decap_4
XFILLER_29_201 vpwr vgnd scs8hd_fill_2
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_41_229 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_226 vpwr vgnd scs8hd_fill_2
XFILLER_17_215 vgnd vpwr scs8hd_decap_8
XFILLER_27_74 vgnd vpwr scs8hd_decap_6
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XFILLER_17_248 vpwr vgnd scs8hd_fill_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
Xmem_top_track_14.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
X_162_ _165_/A _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
X_231_ _231_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_10_210 vgnd vpwr scs8hd_decap_4
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_4
XFILLER_27_195 vpwr vgnd scs8hd_fill_2
XFILLER_19_86 vgnd vpwr scs8hd_decap_8
X_145_ _151_/A _143_/X _145_/Y vgnd vpwr scs8hd_nor2_4
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _190_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_154 vpwr vgnd scs8hd_fill_2
XFILLER_18_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_176 vpwr vgnd scs8hd_fill_2
XFILLER_24_165 vpwr vgnd scs8hd_fill_2
XFILLER_24_154 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_30_135 vgnd vpwr scs8hd_decap_3
XFILLER_30_102 vgnd vpwr scs8hd_decap_6
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
XFILLER_15_121 vgnd vpwr scs8hd_fill_1
X_128_ _125_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_179 vpwr vgnd scs8hd_fill_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_190 vpwr vgnd scs8hd_fill_2
XFILLER_12_157 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_219 vgnd vpwr scs8hd_fill_1
XANTENNA__130__B _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_219 vgnd vpwr scs8hd_fill_1
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_96 vgnd vpwr scs8hd_decap_6
Xmem_right_track_6.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_230 vgnd vpwr scs8hd_fill_1
XFILLER_9_245 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _129_/X vgnd vpwr scs8hd_diode_2
X_161_ _164_/A _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
X_230_ _230_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XANTENNA__136__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_185 vpwr vgnd scs8hd_fill_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_42 vgnd vpwr scs8hd_decap_12
XFILLER_27_141 vpwr vgnd scs8hd_fill_2
X_144_ _129_/X _143_/X _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_4
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_33_177 vpwr vgnd scs8hd_fill_2
XFILLER_33_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_144 vgnd vpwr scs8hd_decap_6
XFILLER_24_100 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ _119_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__B _130_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_158 vpwr vgnd scs8hd_fill_2
XFILLER_21_147 vpwr vgnd scs8hd_fill_2
XFILLER_21_114 vgnd vpwr scs8hd_decap_6
XFILLER_29_258 vgnd vpwr scs8hd_decap_4
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_239 vgnd vpwr scs8hd_decap_3
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_fill_1
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _186_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_34_250 vgnd vpwr scs8hd_decap_8
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_231 vgnd vpwr scs8hd_decap_12
XFILLER_25_272 vgnd vpwr scs8hd_decap_4
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XANTENNA__130__C _134_/C vgnd vpwr scs8hd_diode_2
XANTENNA__139__A _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_253 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_275 vpwr vgnd scs8hd_fill_2
XFILLER_9_235 vgnd vpwr scs8hd_decap_6
XANTENNA__141__B _140_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_194 vpwr vgnd scs8hd_fill_2
X_160_ _163_/A _163_/B _163_/C _153_/D _162_/B vgnd vpwr scs8hd_or4_4
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_223 vgnd vpwr scs8hd_fill_1
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _134_/X vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _096_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_131 vpwr vgnd scs8hd_fill_2
XFILLER_36_142 vgnd vpwr scs8hd_decap_8
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_54 vgnd vpwr scs8hd_decap_6
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_143_ _110_/A _123_/B _153_/C _163_/D _143_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vgnd vpwr scs8hd_decap_3
XANTENNA__147__A _129_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_123 vgnd vpwr scs8hd_fill_1
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vgnd vpwr scs8hd_decap_12
X_126_ _126_/A _123_/B _123_/C _170_/A _127_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_226 vpwr vgnd scs8hd_fill_2
XFILLER_38_237 vgnd vpwr scs8hd_decap_8
XFILLER_29_226 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_148 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _143_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_181 vpwr vgnd scs8hd_fill_2
X_109_ _163_/D _170_/A vgnd vpwr scs8hd_buf_1
XANTENNA__160__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_196 vgnd vpwr scs8hd_fill_1
XFILLER_26_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_240 vgnd vpwr scs8hd_fill_1
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_243 vpwr vgnd scs8hd_fill_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_38_76 vpwr vgnd scs8hd_fill_2
XFILLER_13_254 vgnd vpwr scs8hd_fill_1
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_9_269 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_39_162 vgnd vpwr scs8hd_decap_6
XFILLER_39_184 vgnd vpwr scs8hd_fill_1
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_235 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_154 vgnd vpwr scs8hd_decap_3
XFILLER_27_154 vpwr vgnd scs8hd_fill_2
X_142_ _151_/A _140_/X _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vpwr vgnd scs8hd_fill_2
XFILLER_18_110 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_15_113 vgnd vpwr scs8hd_decap_8
X_125_ _125_/A _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__158__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_127 vgnd vpwr scs8hd_fill_1
XFILLER_21_105 vgnd vpwr scs8hd_decap_3
XFILLER_14_190 vgnd vpwr scs8hd_fill_1
XFILLER_29_205 vgnd vpwr scs8hd_decap_4
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_20_182 vpwr vgnd scs8hd_fill_2
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
X_108_ address[1] enable _163_/D vgnd vpwr scs8hd_nand2_4
XFILLER_11_193 vgnd vpwr scs8hd_decap_4
XFILLER_7_164 vgnd vpwr scs8hd_decap_8
XANTENNA__160__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_40_200 vpwr vgnd scs8hd_fill_2
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_233 vgnd vpwr scs8hd_decap_4
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _170_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_233 vpwr vgnd scs8hd_fill_2
XFILLER_13_211 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_141 vpwr vgnd scs8hd_fill_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_fill_1
XFILLER_10_258 vgnd vpwr scs8hd_decap_12
XFILLER_10_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_111 vgnd vpwr scs8hd_decap_12
XFILLER_36_166 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_199 vpwr vgnd scs8hd_fill_2
X_141_ _129_/X _140_/X _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_78 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _180_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_100 vgnd vpwr scs8hd_fill_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_158 vgnd vpwr scs8hd_decap_4
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_169 vpwr vgnd scs8hd_fill_2
XFILLER_15_158 vpwr vgnd scs8hd_fill_2
X_124_ _119_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_206 vgnd vpwr scs8hd_decap_8
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_20_194 vgnd vpwr scs8hd_decap_3
XFILLER_20_161 vgnd vpwr scs8hd_decap_4
XFILLER_11_150 vgnd vpwr scs8hd_fill_1
X_107_ _125_/A _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XANTENNA__160__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_212 vpwr vgnd scs8hd_fill_2
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_212 vgnd vpwr scs8hd_decap_6
XFILLER_31_245 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__171__B _170_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_245 vgnd vpwr scs8hd_decap_6
XFILLER_22_234 vpwr vgnd scs8hd_fill_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _184_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_38_89 vgnd vpwr scs8hd_decap_3
XFILLER_13_245 vgnd vpwr scs8hd_decap_3
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_123 vgnd vpwr scs8hd_decap_8
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_189 vgnd vpwr scs8hd_decap_8
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_3
X_140_ _110_/A _123_/B _153_/C _153_/D _140_/X vgnd vpwr scs8hd_or4_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _188_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_167 vpwr vgnd scs8hd_fill_2
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XFILLER_18_134 vpwr vgnd scs8hd_fill_2
XFILLER_18_123 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_126 vgnd vpwr scs8hd_decap_3
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
Xmem_top_track_6.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_118 vgnd vpwr scs8hd_decap_6
X_123_ _126_/A _123_/B _123_/C _169_/A _125_/B vgnd vpwr scs8hd_or4_4
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_38_218 vgnd vpwr scs8hd_decap_8
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_129 vpwr vgnd scs8hd_fill_2
XFILLER_11_162 vgnd vpwr scs8hd_decap_12
X_106_ address[0] _125_/A vgnd vpwr scs8hd_buf_1
XANTENNA__160__D _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_80 vpwr vgnd scs8hd_fill_2
XFILLER_7_199 vgnd vpwr scs8hd_decap_12
XFILLER_7_188 vgnd vpwr scs8hd_decap_8
XFILLER_7_177 vpwr vgnd scs8hd_fill_2
XANTENNA__169__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_221 vgnd vpwr scs8hd_fill_1
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_25_276 vgnd vpwr scs8hd_fill_1
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_8
XFILLER_31_268 vpwr vgnd scs8hd_fill_2
XANTENNA__171__C _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_38_68 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_39_198 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_193 vgnd vpwr scs8hd_decap_12
XFILLER_25_91 vpwr vgnd scs8hd_fill_2
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__163__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_41_90 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_108 vgnd vpwr scs8hd_fill_1
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
XFILLER_23_171 vpwr vgnd scs8hd_fill_2
XFILLER_23_160 vpwr vgnd scs8hd_fill_2
X_122_ _163_/A _126_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_182 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_10.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_130 vpwr vgnd scs8hd_fill_2
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
X_105_ _119_/A _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_174 vgnd vpwr scs8hd_fill_1
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XANTENNA__169__C _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_233 vgnd vpwr scs8hd_decap_8
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_91 vpwr vgnd scs8hd_fill_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XFILLER_28_80 vgnd vpwr scs8hd_decap_3
XANTENNA__166__D _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_39_133 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vgnd vpwr scs8hd_decap_8
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_33_139 vpwr vgnd scs8hd_fill_2
XFILLER_26_180 vgnd vpwr scs8hd_decap_4
XFILLER_18_114 vgnd vpwr scs8hd_decap_6
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_117 vgnd vpwr scs8hd_decap_6
XFILLER_17_191 vpwr vgnd scs8hd_fill_2
Xmem_right_track_6.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_194 vgnd vpwr scs8hd_decap_3
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_139 vpwr vgnd scs8hd_fill_2
X_121_ address[3] _163_/A vgnd vpwr scs8hd_inv_8
XFILLER_36_80 vgnd vpwr scs8hd_decap_6
XFILLER_14_172 vgnd vpwr scs8hd_fill_1
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _178_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_209 vgnd vpwr scs8hd_fill_1
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_186 vpwr vgnd scs8hd_fill_2
XFILLER_28_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
X_104_ _110_/A _123_/B _123_/C _169_/A _105_/B vgnd vpwr scs8hd_or4_4
Xmem_top_track_2.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vgnd vpwr scs8hd_decap_6
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_267 vgnd vpwr scs8hd_decap_8
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_204 vgnd vpwr scs8hd_decap_8
XFILLER_25_256 vgnd vpwr scs8hd_decap_8
XFILLER_25_245 vpwr vgnd scs8hd_fill_2
XFILLER_25_201 vpwr vgnd scs8hd_fill_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_237 vgnd vpwr scs8hd_fill_1
XFILLER_16_234 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_22_215 vgnd vpwr scs8hd_decap_4
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
XFILLER_13_237 vgnd vpwr scs8hd_decap_6
XFILLER_13_226 vgnd vpwr scs8hd_decap_4
XFILLER_21_270 vgnd vpwr scs8hd_decap_6
XFILLER_8_230 vgnd vpwr scs8hd_decap_3
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vpwr vgnd scs8hd_fill_2
XFILLER_39_145 vpwr vgnd scs8hd_fill_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _182_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_6
XFILLER_5_200 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_8
XFILLER_35_38 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_27_137 vpwr vgnd scs8hd_fill_2
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_192 vgnd vpwr scs8hd_fill_1
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XFILLER_41_140 vgnd vpwr scs8hd_decap_8
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_151 vpwr vgnd scs8hd_fill_2
XFILLER_25_82 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_120_ _125_/A _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _186_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_210 vgnd vpwr scs8hd_decap_4
XFILLER_37_254 vgnd vpwr scs8hd_decap_8
XFILLER_37_265 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vgnd vpwr scs8hd_fill_1
XFILLER_20_143 vgnd vpwr scs8hd_decap_3
XFILLER_28_210 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
X_103_ _153_/D _169_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_19_265 vgnd vpwr scs8hd_decap_12
XFILLER_19_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_249 vgnd vpwr scs8hd_decap_8
XFILLER_25_268 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_16_246 vgnd vpwr scs8hd_decap_8
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_82 vgnd vpwr scs8hd_decap_3
XFILLER_17_94 vpwr vgnd scs8hd_fill_2
XFILLER_30_271 vgnd vpwr scs8hd_decap_4
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XFILLER_8_242 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_168 vgnd vpwr scs8hd_fill_1
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_212 vgnd vpwr scs8hd_decap_12
XFILLER_5_245 vgnd vpwr scs8hd_decap_8
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XFILLER_18_138 vpwr vgnd scs8hd_fill_2
XFILLER_18_127 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_108 vgnd vpwr scs8hd_decap_8
XFILLER_41_174 vpwr vgnd scs8hd_fill_2
XFILLER_41_163 vpwr vgnd scs8hd_fill_2
XFILLER_41_130 vgnd vpwr scs8hd_decap_6
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_160 vgnd vpwr scs8hd_decap_4
XFILLER_32_163 vpwr vgnd scs8hd_fill_2
XFILLER_23_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_4
XFILLER_14_163 vgnd vpwr scs8hd_decap_3
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_133 vgnd vpwr scs8hd_decap_6
X_102_ address[1] _102_/B _153_/D vgnd vpwr scs8hd_or2_4
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
XFILLER_11_199 vgnd vpwr scs8hd_decap_6
XFILLER_11_177 vpwr vgnd scs8hd_fill_2
XFILLER_7_159 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_203 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_214 vpwr vgnd scs8hd_fill_2
XFILLER_25_236 vgnd vpwr scs8hd_decap_4
XFILLER_25_225 vpwr vgnd scs8hd_fill_2
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_22_228 vgnd vpwr scs8hd_decap_4
XFILLER_22_206 vgnd vpwr scs8hd_decap_8
XFILLER_30_250 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_110 vgnd vpwr scs8hd_fill_1
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XFILLER_5_224 vgnd vpwr scs8hd_decap_12
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_39_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_161 vgnd vpwr scs8hd_fill_1
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_94 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_186 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_197 vgnd vpwr scs8hd_decap_4
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_23_164 vpwr vgnd scs8hd_fill_2
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA__107__A _125_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_223 vpwr vgnd scs8hd_fill_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_267 vgnd vpwr scs8hd_decap_8
XFILLER_28_256 vgnd vpwr scs8hd_decap_8
X_101_ enable _102_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_123 vgnd vpwr scs8hd_decap_8
XFILLER_19_212 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_6
XFILLER_42_270 vgnd vpwr scs8hd_decap_6
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _176_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_229 vpwr vgnd scs8hd_fill_2
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__120__A _125_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_207 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_12_251 vgnd vpwr scs8hd_decap_4
XFILLER_8_200 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_115 vgnd vpwr scs8hd_decap_6
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_181 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _180_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_236 vgnd vpwr scs8hd_decap_8
XFILLER_39_83 vpwr vgnd scs8hd_fill_2
XFILLER_36_107 vpwr vgnd scs8hd_fill_2
XFILLER_39_94 vpwr vgnd scs8hd_fill_2
XFILLER_29_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_8
XFILLER_35_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XFILLER_25_74 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_121 vgnd vpwr scs8hd_decap_3
XFILLER_17_195 vpwr vgnd scs8hd_fill_2
XFILLER_23_143 vpwr vgnd scs8hd_fill_2
XFILLER_23_110 vpwr vgnd scs8hd_fill_2
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_14_143 vgnd vpwr scs8hd_decap_4
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__123__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_157 vpwr vgnd scs8hd_fill_2
XFILLER_20_168 vgnd vpwr scs8hd_decap_3
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
XFILLER_28_202 vgnd vpwr scs8hd_decap_8
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
X_100_ _134_/C _123_/C vgnd vpwr scs8hd_buf_1
XFILLER_11_146 vgnd vpwr scs8hd_decap_4
XANTENNA__118__A _110_/A vgnd vpwr scs8hd_diode_2
X_229_ _229_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_260 vpwr vgnd scs8hd_fill_2
XFILLER_40_219 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _184_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_260 vgnd vpwr scs8hd_decap_12
XFILLER_17_86 vgnd vpwr scs8hd_decap_6
XFILLER_33_74 vgnd vpwr scs8hd_decap_8
Xmem_top_track_6.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__104__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_230 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_85 vgnd vpwr scs8hd_decap_6
XFILLER_8_223 vgnd vpwr scs8hd_fill_1
XANTENNA__115__B _114_/X vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _129_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_62 vgnd vpwr scs8hd_decap_6
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_270 vgnd vpwr scs8hd_decap_4
XFILLER_35_130 vpwr vgnd scs8hd_fill_2
XFILLER_27_108 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_155 vgnd vpwr scs8hd_decap_4
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_133 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_214 vgnd vpwr scs8hd_fill_1
XFILLER_37_236 vpwr vgnd scs8hd_fill_2
XFILLER_37_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
Xmem_top_track_12.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_258 vpwr vgnd scs8hd_fill_2
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
X_159_ _165_/A _159_/B _159_/Y vgnd vpwr scs8hd_nor2_4
X_228_ _228_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA__134__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_228 vgnd vpwr scs8hd_decap_6
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_272 vgnd vpwr scs8hd_decap_3
XFILLER_17_98 vpwr vgnd scs8hd_fill_2
XANTENNA__104__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__129__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_250 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_220 vgnd vpwr scs8hd_decap_4
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _130_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_194 vpwr vgnd scs8hd_fill_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_30 vgnd vpwr scs8hd_decap_12
XFILLER_29_161 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_153 vpwr vgnd scs8hd_fill_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_197 vgnd vpwr scs8hd_decap_8
XFILLER_26_186 vpwr vgnd scs8hd_fill_2
XFILLER_26_164 vgnd vpwr scs8hd_decap_3
XFILLER_25_87 vpwr vgnd scs8hd_fill_2
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_178 vgnd vpwr scs8hd_decap_3
XFILLER_41_167 vgnd vpwr scs8hd_decap_4
XFILLER_41_86 vgnd vpwr scs8hd_decap_4
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_153 vgnd vpwr scs8hd_fill_1
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_145 vgnd vpwr scs8hd_decap_6
XFILLER_32_167 vgnd vpwr scs8hd_decap_8
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_86 vgnd vpwr scs8hd_fill_1
XFILLER_36_97 vgnd vpwr scs8hd_fill_1
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_148 vpwr vgnd scs8hd_fill_2
XFILLER_20_126 vpwr vgnd scs8hd_fill_2
XFILLER_20_115 vgnd vpwr scs8hd_decap_8
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_28_215 vpwr vgnd scs8hd_fill_2
XFILLER_36_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_204 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_207 vgnd vpwr scs8hd_decap_6
XFILLER_27_270 vgnd vpwr scs8hd_decap_6
X_227_ _227_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__118__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_170 vpwr vgnd scs8hd_fill_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
X_158_ _164_/A _159_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__B _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_240 vpwr vgnd scs8hd_fill_2
XFILLER_25_229 vpwr vgnd scs8hd_fill_2
XFILLER_25_218 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_87 vpwr vgnd scs8hd_fill_2
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_30_254 vgnd vpwr scs8hd_fill_1
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_0_114 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _174_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_129 vpwr vgnd scs8hd_fill_2
Xmem_top_track_2.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_151 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_39_42 vgnd vpwr scs8hd_decap_4
XFILLER_30_99 vgnd vpwr scs8hd_fill_1
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_53 vgnd vpwr scs8hd_decap_4
XFILLER_39_75 vgnd vpwr scs8hd_decap_4
XFILLER_29_184 vpwr vgnd scs8hd_fill_2
XFILLER_29_173 vgnd vpwr scs8hd_decap_8
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _140_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_121 vgnd vpwr scs8hd_fill_1
XFILLER_26_121 vgnd vpwr scs8hd_decap_4
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_143 vpwr vgnd scs8hd_fill_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_102 vgnd vpwr scs8hd_decap_8
XFILLER_32_113 vgnd vpwr scs8hd_decap_8
XFILLER_17_187 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_fill_1
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _178_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
X_243_ _243_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_14_168 vgnd vpwr scs8hd_decap_4
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_227 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_157_ _126_/A address[2] _153_/C _163_/D _159_/B vgnd vpwr scs8hd_or4_4
X_226_ _226_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__134__C _134_/C vgnd vpwr scs8hd_diode_2
XANTENNA__118__D _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_193 vgnd vpwr scs8hd_decap_4
XANTENNA__150__B _151_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_263 vpwr vgnd scs8hd_fill_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__145__B _143_/X vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_12_244 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _182_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_259 vgnd vpwr scs8hd_decap_12
XFILLER_8_226 vpwr vgnd scs8hd_fill_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_8
XFILLER_8_204 vpwr vgnd scs8hd_fill_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vpwr vgnd scs8hd_fill_2
XFILLER_38_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_39_87 vgnd vpwr scs8hd_decap_4
XFILLER_39_98 vpwr vgnd scs8hd_fill_2
XANTENNA__126__D _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_199 vgnd vpwr scs8hd_decap_4
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_136 vgnd vpwr scs8hd_fill_1
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_17_199 vgnd vpwr scs8hd_decap_4
XFILLER_17_111 vgnd vpwr scs8hd_decap_8
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_147 vpwr vgnd scs8hd_fill_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vgnd vpwr scs8hd_decap_3
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
X_242_ _242_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_22_191 vpwr vgnd scs8hd_fill_2
XFILLER_37_217 vgnd vpwr scs8hd_decap_4
XANTENNA__148__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_6
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_156_ _165_/A _156_/B _156_/Y vgnd vpwr scs8hd_nor2_4
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__134__D _170_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_187 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_220 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_30_201 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
X_139_ _163_/C _153_/C vgnd vpwr scs8hd_buf_1
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA__156__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_22 vgnd vpwr scs8hd_fill_1
XFILLER_29_197 vpwr vgnd scs8hd_fill_2
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XANTENNA__167__A _166_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_4
XFILLER_35_145 vgnd vpwr scs8hd_decap_8
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_fill_1
XFILLER_41_126 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_137 vgnd vpwr scs8hd_decap_6
XFILLER_17_156 vpwr vgnd scs8hd_fill_2
XFILLER_17_134 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _153_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _198_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_36_89 vgnd vpwr scs8hd_decap_3
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
X_241_ _241_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__164__B _164_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_192 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_4
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ address[0] _165_/A vgnd vpwr scs8hd_buf_1
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_199 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_254 vgnd vpwr scs8hd_decap_4
XFILLER_33_265 vpwr vgnd scs8hd_fill_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_243 vgnd vpwr scs8hd_decap_4
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
XFILLER_15_221 vpwr vgnd scs8hd_fill_2
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_224 vgnd vpwr scs8hd_fill_1
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
X_138_ address[4] _137_/Y _163_/C vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_213 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vgnd vpwr scs8hd_decap_4
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_198 vgnd vpwr scs8hd_decap_4
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _206_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_113 vgnd vpwr scs8hd_decap_8
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vgnd vpwr scs8hd_decap_4
XFILLER_34_190 vpwr vgnd scs8hd_fill_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA__153__D _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_182 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
X_171_ _170_/A _170_/B _165_/A _171_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_171 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vgnd vpwr scs8hd_decap_3
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XFILLER_36_230 vpwr vgnd scs8hd_fill_2
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _176_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_230 vgnd vpwr scs8hd_decap_3
XFILLER_19_208 vpwr vgnd scs8hd_fill_2
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
X_154_ _164_/A _156_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_174 vgnd vpwr scs8hd_decap_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_6
XFILLER_18_274 vgnd vpwr scs8hd_fill_1
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_137_ address[5] _137_/Y vgnd vpwr scs8hd_inv_8
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_247 vgnd vpwr scs8hd_fill_1
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr scs8hd_diode_2
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_177 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_79 vgnd vpwr scs8hd_fill_1
XFILLER_29_144 vpwr vgnd scs8hd_fill_2
XFILLER_29_111 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_158 vpwr vgnd scs8hd_fill_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_147 vgnd vpwr scs8hd_decap_4
XFILLER_26_125 vgnd vpwr scs8hd_fill_1
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_40_150 vgnd vpwr scs8hd_decap_3
XFILLER_31_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
X_170_ _170_/A _170_/B _164_/A _170_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_22_183 vpwr vgnd scs8hd_fill_2
XFILLER_22_150 vgnd vpwr scs8hd_fill_1
XFILLER_14_139 vpwr vgnd scs8hd_fill_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_8
XFILLER_26_80 vpwr vgnd scs8hd_fill_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
X_153_ _126_/A address[2] _153_/C _153_/D _156_/B vgnd vpwr scs8hd_or4_4
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_212 vgnd vpwr scs8hd_decap_8
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vpwr vgnd scs8hd_fill_2
XFILLER_15_267 vgnd vpwr scs8hd_decap_8
XFILLER_15_245 vgnd vpwr scs8hd_decap_3
XFILLER_15_201 vgnd vpwr scs8hd_fill_1
X_136_ _151_/A _134_/X _136_/Y vgnd vpwr scs8hd_nor2_4
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_21_204 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_215 vgnd vpwr scs8hd_decap_3
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XFILLER_12_248 vgnd vpwr scs8hd_fill_1
XFILLER_8_208 vgnd vpwr scs8hd_decap_6
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _119_/A _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_12.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_241 vgnd vpwr scs8hd_fill_1
XFILLER_38_145 vgnd vpwr scs8hd_decap_4
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_80 vgnd vpwr scs8hd_fill_1
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_31_92 vgnd vpwr scs8hd_fill_1
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_173 vpwr vgnd scs8hd_fill_2
XFILLER_31_195 vpwr vgnd scs8hd_fill_2
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_240 vpwr vgnd scs8hd_fill_2
XFILLER_22_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_210 vgnd vpwr scs8hd_decap_4
XFILLER_36_243 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_210 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_254 vpwr vgnd scs8hd_fill_2
X_152_ _096_/A _164_/A vgnd vpwr scs8hd_buf_1
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _196_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_80 vgnd vpwr scs8hd_decap_4
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_254 vgnd vpwr scs8hd_decap_8
XFILLER_18_243 vpwr vgnd scs8hd_fill_2
XFILLER_33_224 vpwr vgnd scs8hd_fill_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_224 vgnd vpwr scs8hd_decap_3
XFILLER_24_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_227 vgnd vpwr scs8hd_fill_1
XFILLER_30_205 vgnd vpwr scs8hd_decap_8
XFILLER_15_235 vpwr vgnd scs8hd_fill_2
X_135_ _129_/X _134_/X _135_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_21_238 vgnd vpwr scs8hd_decap_4
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vgnd vpwr scs8hd_decap_8
XFILLER_20_260 vgnd vpwr scs8hd_decap_12
XFILLER_18_93 vgnd vpwr scs8hd_decap_4
XFILLER_7_231 vpwr vgnd scs8hd_fill_2
X_118_ _110_/A _114_/X _123_/C _170_/A _119_/B vgnd vpwr scs8hd_or4_4
Xmem_right_track_4.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_113 vgnd vpwr scs8hd_decap_8
XFILLER_38_124 vgnd vpwr scs8hd_decap_8
XFILLER_38_168 vgnd vpwr scs8hd_decap_6
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_26 vpwr vgnd scs8hd_fill_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_168 vgnd vpwr scs8hd_decap_3
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XFILLER_29_92 vgnd vpwr scs8hd_decap_6
XFILLER_35_127 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_138 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_34_182 vgnd vpwr scs8hd_decap_8
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_17_149 vgnd vpwr scs8hd_decap_4
XFILLER_40_174 vgnd vpwr scs8hd_decap_8
XFILLER_40_163 vgnd vpwr scs8hd_decap_8
XFILLER_31_152 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _204_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_13_163 vgnd vpwr scs8hd_decap_8
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_258 vgnd vpwr scs8hd_decap_12
XFILLER_27_266 vpwr vgnd scs8hd_fill_2
X_151_ _151_/A _151_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_236 vpwr vgnd scs8hd_fill_2
XFILLER_18_266 vgnd vpwr scs8hd_decap_8
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_203 vpwr vgnd scs8hd_fill_2
XFILLER_15_225 vgnd vpwr scs8hd_fill_1
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _174_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_8
X_134_ _126_/A _114_/X _134_/C _170_/A _134_/X vgnd vpwr scs8hd_or4_4
XFILLER_21_217 vpwr vgnd scs8hd_fill_2
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
XFILLER_20_272 vgnd vpwr scs8hd_decap_3
X_117_ _125_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_265 vpwr vgnd scs8hd_fill_2
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_39_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_128 vgnd vpwr scs8hd_fill_1
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_142 vgnd vpwr scs8hd_decap_8
XFILLER_40_131 vgnd vpwr scs8hd_decap_6
XFILLER_25_150 vgnd vpwr scs8hd_decap_4
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_40_186 vgnd vpwr scs8hd_decap_4
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_131 vgnd vpwr scs8hd_decap_4
XFILLER_16_194 vgnd vpwr scs8hd_decap_3
XFILLER_16_183 vgnd vpwr scs8hd_decap_6
XFILLER_22_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_175 vgnd vpwr scs8hd_decap_8
XFILLER_13_142 vpwr vgnd scs8hd_fill_2
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_36_223 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_223 vgnd vpwr scs8hd_decap_4
X_150_ _129_/X _151_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_189 vpwr vgnd scs8hd_fill_2
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_223 vgnd vpwr scs8hd_fill_1
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
X_133_ _151_/A _130_/X _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
X_116_ _119_/A _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_273 vgnd vpwr scs8hd_decap_4
XFILLER_11_262 vgnd vpwr scs8hd_decap_4
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_7_211 vgnd vpwr scs8hd_decap_12
XFILLER_29_115 vpwr vgnd scs8hd_fill_2
XFILLER_4_258 vgnd vpwr scs8hd_decap_12
XFILLER_28_192 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_84 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_254 vgnd vpwr scs8hd_decap_3
XFILLER_39_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_187 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_8
XFILLER_9_158 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_6
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_235 vgnd vpwr scs8hd_decap_8
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_260 vgnd vpwr scs8hd_decap_3
XFILLER_24_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_132_ address[0] _151_/A vgnd vpwr scs8hd_buf_1
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_260 vpwr vgnd scs8hd_fill_2
XFILLER_23_74 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA__110__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_208 vgnd vpwr scs8hd_decap_3
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _194_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
X_115_ _110_/A _114_/X _123_/C _169_/A _116_/B vgnd vpwr scs8hd_or4_4
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_223 vgnd vpwr scs8hd_decap_8
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_160 vgnd vpwr scs8hd_decap_4
XFILLER_29_127 vpwr vgnd scs8hd_fill_2
XFILLER_37_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XANTENNA__116__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_26_108 vgnd vpwr scs8hd_decap_4
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_193 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _198_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_119 vgnd vpwr scs8hd_fill_1
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vgnd vpwr scs8hd_decap_3
XFILLER_0_262 vgnd vpwr scs8hd_decap_12
XFILLER_16_163 vgnd vpwr scs8hd_decap_3
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_177 vgnd vpwr scs8hd_decap_4
XFILLER_31_199 vpwr vgnd scs8hd_fill_2
.ends

