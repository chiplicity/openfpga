VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 197.160 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 2.400 ;
    END
  END Test_en
  PIN bottom_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END bottom_width_0_height_0__pin_16_
  PIN bottom_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END bottom_width_0_height_0__pin_17_
  PIN bottom_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END bottom_width_0_height_0__pin_18_
  PIN bottom_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.400 ;
    END
  END bottom_width_0_height_0__pin_19_
  PIN bottom_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END bottom_width_0_height_0__pin_20_
  PIN bottom_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 2.400 ;
    END
  END bottom_width_0_height_0__pin_21_
  PIN bottom_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END bottom_width_0_height_0__pin_22_
  PIN bottom_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 2.400 ;
    END
  END bottom_width_0_height_0__pin_23_
  PIN bottom_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 2.400 ;
    END
  END bottom_width_0_height_0__pin_24_
  PIN bottom_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END bottom_width_0_height_0__pin_25_
  PIN bottom_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 2.400 ;
    END
  END bottom_width_0_height_0__pin_26_
  PIN bottom_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END bottom_width_0_height_0__pin_27_
  PIN bottom_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END bottom_width_0_height_0__pin_28_
  PIN bottom_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 2.400 ;
    END
  END bottom_width_0_height_0__pin_29_
  PIN bottom_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END bottom_width_0_height_0__pin_30_
  PIN bottom_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 2.400 ;
    END
  END bottom_width_0_height_0__pin_31_
  PIN bottom_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 2.400 ;
    END
  END bottom_width_0_height_0__pin_42_lower
  PIN bottom_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END bottom_width_0_height_0__pin_42_upper
  PIN bottom_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 2.400 ;
    END
  END bottom_width_0_height_0__pin_43_lower
  PIN bottom_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 2.400 ;
    END
  END bottom_width_0_height_0__pin_43_upper
  PIN bottom_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 2.400 ;
    END
  END bottom_width_0_height_0__pin_44_lower
  PIN bottom_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.400 ;
    END
  END bottom_width_0_height_0__pin_44_upper
  PIN bottom_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 2.400 ;
    END
  END bottom_width_0_height_0__pin_45_lower
  PIN bottom_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END bottom_width_0_height_0__pin_45_upper
  PIN bottom_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.400 ;
    END
  END bottom_width_0_height_0__pin_46_lower
  PIN bottom_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END bottom_width_0_height_0__pin_46_upper
  PIN bottom_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 2.400 ;
    END
  END bottom_width_0_height_0__pin_47_lower
  PIN bottom_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.400 ;
    END
  END bottom_width_0_height_0__pin_47_upper
  PIN bottom_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 2.400 ;
    END
  END bottom_width_0_height_0__pin_48_lower
  PIN bottom_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END bottom_width_0_height_0__pin_48_upper
  PIN bottom_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 2.400 ;
    END
  END bottom_width_0_height_0__pin_49_lower
  PIN bottom_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.400 ;
    END
  END bottom_width_0_height_0__pin_49_upper
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 2.400 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 2.400 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 59.880 200.000 60.480 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 2.400 ;
    END
  END clk
  PIN left_width_0_height_0__pin_52_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_width_0_height_0__pin_52_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 65.320 200.000 65.920 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 122.440 200.000 123.040 ;
    END
  END right_width_0_height_0__pin_10_
  PIN right_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 127.880 200.000 128.480 ;
    END
  END right_width_0_height_0__pin_11_
  PIN right_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 134.000 200.000 134.600 ;
    END
  END right_width_0_height_0__pin_12_
  PIN right_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 139.440 200.000 140.040 ;
    END
  END right_width_0_height_0__pin_13_
  PIN right_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 145.560 200.000 146.160 ;
    END
  END right_width_0_height_0__pin_14_
  PIN right_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 151.000 200.000 151.600 ;
    END
  END right_width_0_height_0__pin_15_
  PIN right_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 70.760 200.000 71.360 ;
    END
  END right_width_0_height_0__pin_1_
  PIN right_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 76.880 200.000 77.480 ;
    END
  END right_width_0_height_0__pin_2_
  PIN right_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 25.200 200.000 25.800 ;
    END
  END right_width_0_height_0__pin_34_lower
  PIN right_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 156.440 200.000 157.040 ;
    END
  END right_width_0_height_0__pin_34_upper
  PIN right_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 31.320 200.000 31.920 ;
    END
  END right_width_0_height_0__pin_35_lower
  PIN right_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 162.560 200.000 163.160 ;
    END
  END right_width_0_height_0__pin_35_upper
  PIN right_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 36.760 200.000 37.360 ;
    END
  END right_width_0_height_0__pin_36_lower
  PIN right_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 168.000 200.000 168.600 ;
    END
  END right_width_0_height_0__pin_36_upper
  PIN right_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 42.200 200.000 42.800 ;
    END
  END right_width_0_height_0__pin_37_lower
  PIN right_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 174.120 200.000 174.720 ;
    END
  END right_width_0_height_0__pin_37_upper
  PIN right_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 48.320 200.000 48.920 ;
    END
  END right_width_0_height_0__pin_38_lower
  PIN right_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 179.560 200.000 180.160 ;
    END
  END right_width_0_height_0__pin_38_upper
  PIN right_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 53.760 200.000 54.360 ;
    END
  END right_width_0_height_0__pin_39_lower
  PIN right_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 185.000 200.000 185.600 ;
    END
  END right_width_0_height_0__pin_39_upper
  PIN right_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 82.320 200.000 82.920 ;
    END
  END right_width_0_height_0__pin_3_
  PIN right_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 13.640 200.000 14.240 ;
    END
  END right_width_0_height_0__pin_40_lower
  PIN right_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 191.120 200.000 191.720 ;
    END
  END right_width_0_height_0__pin_40_upper
  PIN right_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 19.760 200.000 20.360 ;
    END
  END right_width_0_height_0__pin_41_lower
  PIN right_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 196.560 200.000 197.160 ;
    END
  END right_width_0_height_0__pin_41_upper
  PIN right_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 88.440 200.000 89.040 ;
    END
  END right_width_0_height_0__pin_4_
  PIN right_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 93.880 200.000 94.480 ;
    END
  END right_width_0_height_0__pin_5_
  PIN right_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 99.320 200.000 99.920 ;
    END
  END right_width_0_height_0__pin_6_
  PIN right_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 105.440 200.000 106.040 ;
    END
  END right_width_0_height_0__pin_7_
  PIN right_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 110.880 200.000 111.480 ;
    END
  END right_width_0_height_0__pin_8_
  PIN right_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 117.000 200.000 117.600 ;
    END
  END right_width_0_height_0__pin_9_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.760 200.000 3.360 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 8.200 200.000 8.800 ;
    END
  END top_width_0_height_0__pin_33_
  PIN vpwr
    USE POWER ; 
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 2.850 2.680 197.250 197.045 ;
        RECT 3.410 2.400 8.090 2.680 ;
        RECT 8.930 2.400 13.610 2.680 ;
        RECT 14.450 2.400 19.130 2.680 ;
        RECT 19.970 2.400 24.650 2.680 ;
        RECT 25.490 2.400 30.170 2.680 ;
        RECT 31.010 2.400 35.690 2.680 ;
        RECT 36.530 2.400 41.210 2.680 ;
        RECT 42.050 2.400 46.730 2.680 ;
        RECT 47.570 2.400 52.250 2.680 ;
        RECT 53.090 2.400 57.770 2.680 ;
        RECT 58.610 2.400 63.290 2.680 ;
        RECT 64.130 2.400 69.270 2.680 ;
        RECT 70.110 2.400 74.790 2.680 ;
        RECT 75.630 2.400 80.310 2.680 ;
        RECT 81.150 2.400 85.830 2.680 ;
        RECT 86.670 2.400 91.350 2.680 ;
        RECT 92.190 2.400 96.870 2.680 ;
        RECT 97.710 2.400 102.390 2.680 ;
        RECT 103.230 2.400 107.910 2.680 ;
        RECT 108.750 2.400 113.430 2.680 ;
        RECT 114.270 2.400 118.950 2.680 ;
        RECT 119.790 2.400 124.470 2.680 ;
        RECT 125.310 2.400 129.990 2.680 ;
        RECT 130.830 2.400 135.970 2.680 ;
        RECT 136.810 2.400 141.490 2.680 ;
        RECT 142.330 2.400 147.010 2.680 ;
        RECT 147.850 2.400 152.530 2.680 ;
        RECT 153.370 2.400 158.050 2.680 ;
        RECT 158.890 2.400 163.570 2.680 ;
        RECT 164.410 2.400 169.090 2.680 ;
        RECT 169.930 2.400 174.610 2.680 ;
        RECT 175.450 2.400 180.130 2.680 ;
        RECT 180.970 2.400 185.650 2.680 ;
        RECT 186.490 2.400 191.170 2.680 ;
        RECT 192.010 2.400 196.690 2.680 ;
      LAYER met3 ;
        RECT 2.400 196.160 197.200 197.025 ;
        RECT 2.400 192.120 197.600 196.160 ;
        RECT 2.400 190.720 197.200 192.120 ;
        RECT 2.400 186.000 197.600 190.720 ;
        RECT 2.400 184.600 197.200 186.000 ;
        RECT 2.400 180.560 197.600 184.600 ;
        RECT 2.400 179.160 197.200 180.560 ;
        RECT 2.400 175.120 197.600 179.160 ;
        RECT 2.400 173.720 197.200 175.120 ;
        RECT 2.400 169.000 197.600 173.720 ;
        RECT 2.400 167.640 197.200 169.000 ;
        RECT 2.800 167.600 197.200 167.640 ;
        RECT 2.800 166.240 197.600 167.600 ;
        RECT 2.400 163.560 197.600 166.240 ;
        RECT 2.400 162.160 197.200 163.560 ;
        RECT 2.400 157.440 197.600 162.160 ;
        RECT 2.400 156.040 197.200 157.440 ;
        RECT 2.400 152.000 197.600 156.040 ;
        RECT 2.400 150.600 197.200 152.000 ;
        RECT 2.400 146.560 197.600 150.600 ;
        RECT 2.400 145.160 197.200 146.560 ;
        RECT 2.400 140.440 197.600 145.160 ;
        RECT 2.400 139.040 197.200 140.440 ;
        RECT 2.400 135.000 197.600 139.040 ;
        RECT 2.400 133.600 197.200 135.000 ;
        RECT 2.400 128.880 197.600 133.600 ;
        RECT 2.400 127.480 197.200 128.880 ;
        RECT 2.400 123.440 197.600 127.480 ;
        RECT 2.400 122.040 197.200 123.440 ;
        RECT 2.400 118.000 197.600 122.040 ;
        RECT 2.400 116.600 197.200 118.000 ;
        RECT 2.400 111.880 197.600 116.600 ;
        RECT 2.400 110.480 197.200 111.880 ;
        RECT 2.400 106.440 197.600 110.480 ;
        RECT 2.400 105.040 197.200 106.440 ;
        RECT 2.400 101.000 197.600 105.040 ;
        RECT 2.800 100.320 197.600 101.000 ;
        RECT 2.800 99.600 197.200 100.320 ;
        RECT 2.400 98.920 197.200 99.600 ;
        RECT 2.400 94.880 197.600 98.920 ;
        RECT 2.400 93.480 197.200 94.880 ;
        RECT 2.400 89.440 197.600 93.480 ;
        RECT 2.400 88.040 197.200 89.440 ;
        RECT 2.400 83.320 197.600 88.040 ;
        RECT 2.400 81.920 197.200 83.320 ;
        RECT 2.400 77.880 197.600 81.920 ;
        RECT 2.400 76.480 197.200 77.880 ;
        RECT 2.400 71.760 197.600 76.480 ;
        RECT 2.400 70.360 197.200 71.760 ;
        RECT 2.400 66.320 197.600 70.360 ;
        RECT 2.400 64.920 197.200 66.320 ;
        RECT 2.400 60.880 197.600 64.920 ;
        RECT 2.400 59.480 197.200 60.880 ;
        RECT 2.400 54.760 197.600 59.480 ;
        RECT 2.400 53.360 197.200 54.760 ;
        RECT 2.400 49.320 197.600 53.360 ;
        RECT 2.400 47.920 197.200 49.320 ;
        RECT 2.400 43.200 197.600 47.920 ;
        RECT 2.400 41.800 197.200 43.200 ;
        RECT 2.400 37.760 197.600 41.800 ;
        RECT 2.400 36.360 197.200 37.760 ;
        RECT 2.400 34.360 197.600 36.360 ;
        RECT 2.800 32.960 197.600 34.360 ;
        RECT 2.400 32.320 197.600 32.960 ;
        RECT 2.400 30.920 197.200 32.320 ;
        RECT 2.400 26.200 197.600 30.920 ;
        RECT 2.400 24.800 197.200 26.200 ;
        RECT 2.400 20.760 197.600 24.800 ;
        RECT 2.400 19.360 197.200 20.760 ;
        RECT 2.400 14.640 197.600 19.360 ;
        RECT 2.400 13.240 197.200 14.640 ;
        RECT 2.400 9.200 197.600 13.240 ;
        RECT 2.400 7.800 197.200 9.200 ;
        RECT 2.400 3.760 197.600 7.800 ;
        RECT 2.400 2.895 197.200 3.760 ;
      LAYER met4 ;
        RECT 174.640 10.640 179.105 187.920 ;
  END
END grid_clb
END LIBRARY

