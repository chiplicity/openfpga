* NGSPICE file created from sb_3__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_3__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_
+ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ left_top_grid_pin_10_ top_left_grid_pin_13_
+ top_right_grid_pin_11_ top_right_grid_pin_13_ top_right_grid_pin_15_ top_right_grid_pin_1_
+ top_right_grid_pin_3_ top_right_grid_pin_5_ top_right_grid_pin_7_ top_right_grid_pin_9_
+ vpwr vgnd
XFILLER_39_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_74 vpwr vgnd scs8hd_fill_2
XFILLER_26_96 vgnd vpwr scs8hd_decap_4
XFILLER_42_84 vgnd vpwr scs8hd_decap_8
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_115 vgnd vpwr scs8hd_decap_6
XFILLER_36_203 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_7_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_21 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vpwr vgnd scs8hd_fill_2
XFILLER_37_95 vpwr vgnd scs8hd_fill_2
XFILLER_33_239 vgnd vpwr scs8hd_decap_4
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_206 vgnd vpwr scs8hd_decap_8
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _190_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_209 vgnd vpwr scs8hd_decap_4
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
X_131_ _129_/X _133_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__110__C _118_/C vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_86 vgnd vpwr scs8hd_decap_4
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd vpwr
+ scs8hd_diode_2
X_114_ _114_/A _118_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_106 vpwr vgnd scs8hd_fill_2
XFILLER_22_7 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _172_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_172 vpwr vgnd scs8hd_fill_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_10 vgnd vpwr scs8hd_decap_4
XFILLER_20_32 vgnd vpwr scs8hd_decap_8
XFILLER_20_76 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _194_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_142 vgnd vpwr scs8hd_decap_8
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_15_21 vpwr vgnd scs8hd_fill_2
XFILLER_25_175 vgnd vpwr scs8hd_decap_6
XFILLER_31_31 vgnd vpwr scs8hd_decap_3
XFILLER_25_197 vgnd vpwr scs8hd_fill_1
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_39_212 vpwr vgnd scs8hd_fill_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XFILLER_22_123 vpwr vgnd scs8hd_fill_2
Xmem_top_track_4.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_26_86 vgnd vpwr scs8hd_decap_3
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_204 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_11 vgnd vpwr scs8hd_fill_1
XFILLER_12_55 vgnd vpwr scs8hd_fill_1
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA__140__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_5_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_130_ _134_/A _118_/B _100_/A _104_/D _133_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_76 vpwr vgnd scs8hd_fill_2
XANTENNA__110__D _109_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XANTENNA__135__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_4
XFILLER_18_98 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
X_113_ address[2] _114_/A vgnd vpwr scs8hd_inv_8
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_6
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_55 vgnd vpwr scs8hd_decap_8
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_20 vpwr vgnd scs8hd_fill_2
XFILLER_6_79 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_151 vgnd vpwr scs8hd_decap_12
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_165 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_102 vgnd vpwr scs8hd_decap_8
XFILLER_15_55 vgnd vpwr scs8hd_decap_4
XFILLER_25_110 vpwr vgnd scs8hd_fill_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_97 vgnd vpwr scs8hd_decap_8
XFILLER_42_75 vgnd vpwr scs8hd_decap_6
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_216 vgnd vpwr scs8hd_decap_12
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_6 vgnd vpwr scs8hd_decap_8
XANTENNA__140__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_9_24 vpwr vgnd scs8hd_fill_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_79 vgnd vpwr scs8hd_decap_12
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_6
XANTENNA__151__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_54 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_4
X_112_ _125_/A _112_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_65 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_3_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_119 vgnd vpwr scs8hd_decap_4
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_152 vgnd vpwr scs8hd_decap_4
XFILLER_20_23 vgnd vpwr scs8hd_decap_8
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XFILLER_34_111 vpwr vgnd scs8hd_fill_2
XFILLER_19_163 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_147 vgnd vpwr scs8hd_decap_6
XFILLER_40_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_125 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XFILLER_15_89 vgnd vpwr scs8hd_decap_6
XFILLER_25_133 vpwr vgnd scs8hd_fill_2
XFILLER_31_99 vpwr vgnd scs8hd_fill_2
XFILLER_31_77 vgnd vpwr scs8hd_fill_1
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_136 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XFILLER_22_136 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_228 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_37_32 vgnd vpwr scs8hd_decap_12
XFILLER_37_21 vpwr vgnd scs8hd_fill_2
XFILLER_37_10 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_76 vpwr vgnd scs8hd_fill_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_15.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__C _143_/C vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_47 vgnd vpwr scs8hd_decap_8
XFILLER_9_36 vgnd vpwr scs8hd_decap_4
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_6
XFILLER_18_56 vpwr vgnd scs8hd_fill_2
X_111_ _127_/A _112_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XANTENNA__146__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_33 vgnd vpwr scs8hd_decap_3
XFILLER_29_99 vpwr vgnd scs8hd_fill_2
XFILLER_28_186 vgnd vpwr scs8hd_decap_4
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_29_66 vgnd vpwr scs8hd_fill_1
XANTENNA__157__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vgnd vpwr scs8hd_decap_8
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_1_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_123 vgnd vpwr scs8hd_fill_1
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_112 vgnd vpwr scs8hd_decap_4
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_159 vpwr vgnd scs8hd_fill_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_204 vgnd vpwr scs8hd_decap_4
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _192_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_1.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_26_78 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _109_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_25 vpwr vgnd scs8hd_fill_2
XFILLER_12_47 vgnd vpwr scs8hd_decap_8
XFILLER_12_69 vpwr vgnd scs8hd_fill_2
XFILLER_37_66 vgnd vpwr scs8hd_decap_3
XFILLER_37_44 vgnd vpwr scs8hd_decap_12
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_99 vgnd vpwr scs8hd_decap_4
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_111 vgnd vpwr scs8hd_decap_8
XANTENNA__140__D _140_/D vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_13 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
X_110_ _118_/A _104_/B _118_/C _109_/X _112_/B vgnd vpwr scs8hd_or4_4
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
X_239_ _239_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _160_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_132 vgnd vpwr scs8hd_decap_4
XFILLER_37_187 vpwr vgnd scs8hd_fill_2
XFILLER_37_176 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_78 vpwr vgnd scs8hd_fill_2
XFILLER_28_110 vgnd vpwr scs8hd_fill_1
XFILLER_28_132 vpwr vgnd scs8hd_fill_2
XFILLER_28_165 vgnd vpwr scs8hd_decap_8
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vgnd vpwr scs8hd_decap_3
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_143 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_47 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__143__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_216 vgnd vpwr scs8hd_decap_4
XFILLER_39_227 vgnd vpwr scs8hd_decap_12
XANTENNA__168__A _104_/D vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_81 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_127 vgnd vpwr scs8hd_decap_12
XFILLER_26_57 vgnd vpwr scs8hd_decap_8
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_160 vpwr vgnd scs8hd_fill_2
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_89 vgnd vpwr scs8hd_decap_4
XFILLER_37_56 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XFILLER_32_200 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C _143_/C vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_36 vgnd vpwr scs8hd_fill_1
XFILLER_18_69 vpwr vgnd scs8hd_fill_2
XFILLER_34_46 vgnd vpwr scs8hd_decap_8
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
X_238_ _238_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__D _140_/D vgnd vpwr scs8hd_diode_2
X_169_ _104_/D _168_/B _155_/X _169_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_1_50 vgnd vpwr scs8hd_decap_8
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_17 vgnd vpwr scs8hd_decap_12
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_169 vgnd vpwr scs8hd_decap_8
XFILLER_34_125 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_33_191 vgnd vpwr scs8hd_decap_12
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_239 vgnd vpwr scs8hd_decap_4
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_106 vpwr vgnd scs8hd_fill_2
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_139 vgnd vpwr scs8hd_decap_12
XFILLER_26_36 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_212 vpwr vgnd scs8hd_fill_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XANTENNA__149__D _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_36 vgnd vpwr scs8hd_fill_1
XFILLER_18_48 vgnd vpwr scs8hd_decap_8
XFILLER_34_69 vpwr vgnd scs8hd_fill_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
X_237_ _237_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_168_ _104_/D _168_/B _152_/X _168_/Y vgnd vpwr scs8hd_nor3_4
X_099_ address[4] address[5] _100_/A vgnd vpwr scs8hd_or2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_3
XFILLER_37_156 vgnd vpwr scs8hd_fill_1
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_145 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_115 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__157__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_137 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _152_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_173 vpwr vgnd scs8hd_fill_2
XFILLER_30_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_50 vgnd vpwr scs8hd_decap_8
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vgnd vpwr scs8hd_decap_4
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _190_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_38 vpwr vgnd scs8hd_fill_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_60 vgnd vpwr scs8hd_fill_1
Xmem_top_track_4.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_81 vgnd vpwr scs8hd_decap_3
XFILLER_40_91 vgnd vpwr scs8hd_fill_1
X_236_ _236_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_167_ _166_/X _168_/B vgnd vpwr scs8hd_buf_1
X_098_ address[2] _104_/B vgnd vpwr scs8hd_buf_1
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XFILLER_28_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_119 vgnd vpwr scs8hd_decap_4
XFILLER_15_17 vpwr vgnd scs8hd_fill_2
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_182 vgnd vpwr scs8hd_decap_12
XFILLER_39_208 vgnd vpwr scs8hd_fill_1
XFILLER_11_7 vgnd vpwr scs8hd_decap_3
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_22_119 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_8
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_241 vgnd vpwr scs8hd_decap_3
XFILLER_16_60 vpwr vgnd scs8hd_fill_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_32_81 vpwr vgnd scs8hd_fill_2
XFILLER_32_70 vgnd vpwr scs8hd_decap_4
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_200 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
Xmem_top_track_10.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_81 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_17 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vpwr vgnd scs8hd_fill_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_60 vgnd vpwr scs8hd_decap_3
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
X_235_ _235_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_40_81 vpwr vgnd scs8hd_fill_2
XFILLER_40_70 vpwr vgnd scs8hd_fill_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_166_ address[3] address[2] address[4] _138_/B _166_/X vgnd vpwr scs8hd_or4_4
X_097_ address[3] _118_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_6 vgnd vpwr scs8hd_decap_8
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_29_38 vgnd vpwr scs8hd_decap_3
XFILLER_36_191 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_73 vgnd vpwr scs8hd_decap_4
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_19_147 vpwr vgnd scs8hd_fill_2
XFILLER_35_70 vpwr vgnd scs8hd_fill_2
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ address[3] _118_/B _143_/C _109_/A _149_/X vgnd vpwr scs8hd_or4_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_29 vgnd vpwr scs8hd_decap_3
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_194 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_197 vgnd vpwr scs8hd_decap_12
XFILLER_30_186 vgnd vpwr scs8hd_decap_8
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_153 vgnd vpwr scs8hd_fill_1
XFILLER_21_164 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_35_212 vgnd vpwr scs8hd_decap_12
XFILLER_26_201 vgnd vpwr scs8hd_decap_12
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_51 vgnd vpwr scs8hd_decap_3
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XFILLER_13_84 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_207 vgnd vpwr scs8hd_decap_6
XFILLER_34_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
X_234_ _234_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_165_ _155_/X _164_/B _165_/Y vgnd vpwr scs8hd_nor2_4
X_096_ _096_/A _127_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_159 vpwr vgnd scs8hd_fill_2
XFILLER_1_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_15.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_126 vgnd vpwr scs8hd_decap_4
XFILLER_10_41 vgnd vpwr scs8hd_decap_12
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_19_50 vpwr vgnd scs8hd_fill_2
XFILLER_19_94 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vpwr vgnd scs8hd_fill_2
XFILLER_42_162 vgnd vpwr scs8hd_decap_12
XFILLER_34_107 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_170 vgnd vpwr scs8hd_decap_3
XFILLER_27_192 vgnd vpwr scs8hd_decap_12
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
X_148_ _133_/A _148_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_fill_1
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_33_173 vgnd vpwr scs8hd_decap_4
XFILLER_31_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_4
XFILLER_30_143 vgnd vpwr scs8hd_decap_8
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XANTENNA__103__A _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_224 vgnd vpwr scs8hd_decap_12
XFILLER_37_28 vpwr vgnd scs8hd_fill_2
XFILLER_37_17 vpwr vgnd scs8hd_fill_2
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_233_ _233_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_164_ _152_/X _164_/B _164_/Y vgnd vpwr scs8hd_nor2_4
X_095_ address[0] _096_/A vgnd vpwr scs8hd_inv_8
XFILLER_37_138 vgnd vpwr scs8hd_decap_3
XANTENNA__111__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_149 vgnd vpwr scs8hd_decap_4
XFILLER_10_53 vgnd vpwr scs8hd_decap_4
XFILLER_34_119 vgnd vpwr scs8hd_decap_4
XFILLER_19_62 vpwr vgnd scs8hd_fill_2
XFILLER_42_174 vgnd vpwr scs8hd_decap_12
XFILLER_42_141 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_4
XFILLER_35_83 vpwr vgnd scs8hd_fill_2
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
X_147_ _129_/X _148_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_152 vpwr vgnd scs8hd_fill_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_16_108 vpwr vgnd scs8hd_fill_2
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
XFILLER_21_74 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _188_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_122 vgnd vpwr scs8hd_decap_8
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_32_51 vgnd vpwr scs8hd_decap_4
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _206_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_35_236 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_97 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XFILLER_39_191 vpwr vgnd scs8hd_fill_2
X_232_ _232_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_40_62 vgnd vpwr scs8hd_decap_8
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_163_ _121_/Y _114_/A _138_/Y _109_/A _164_/B vgnd vpwr scs8hd_or4_4
XANTENNA__111__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
XFILLER_36_161 vpwr vgnd scs8hd_fill_2
XFILLER_27_150 vgnd vpwr scs8hd_decap_3
XFILLER_42_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_62 vgnd vpwr scs8hd_fill_1
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__122__A _121_/Y vgnd vpwr scs8hd_diode_2
X_146_ address[3] _118_/B _143_/C _140_/D _148_/B vgnd vpwr scs8hd_or4_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_11.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_7_22 vpwr vgnd scs8hd_fill_2
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _125_/A vgnd vpwr scs8hd_diode_2
X_129_ _096_/A _129_/X vgnd vpwr scs8hd_buf_1
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
XFILLER_38_201 vgnd vpwr scs8hd_decap_12
XFILLER_21_112 vgnd vpwr scs8hd_decap_4
XFILLER_21_156 vgnd vpwr scs8hd_fill_1
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_16_64 vgnd vpwr scs8hd_decap_3
XFILLER_16_86 vgnd vpwr scs8hd_decap_6
XFILLER_32_85 vgnd vpwr scs8hd_decap_4
XFILLER_32_74 vgnd vpwr scs8hd_fill_1
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_119 vgnd vpwr scs8hd_decap_3
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_3
Xmem_left_track_7.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_85 vpwr vgnd scs8hd_fill_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__130__A _134_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XFILLER_13_32 vpwr vgnd scs8hd_fill_2
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
Xmem_top_track_14.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
X_231_ _231_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_162_ _155_/X _160_/X _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_42 vpwr vgnd scs8hd_fill_2
XFILLER_24_86 vgnd vpwr scs8hd_decap_4
XFILLER_40_85 vgnd vpwr scs8hd_decap_6
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
X_145_ _133_/A _145_/B _145_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_187 vpwr vgnd scs8hd_fill_2
XFILLER_33_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_110 vgnd vpwr scs8hd_decap_3
XFILLER_24_143 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_165 vpwr vgnd scs8hd_fill_2
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_110 vgnd vpwr scs8hd_decap_6
XFILLER_15_132 vgnd vpwr scs8hd_decap_12
X_128_ _125_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_fill_1
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_168 vgnd vpwr scs8hd_fill_1
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_102 vgnd vpwr scs8hd_decap_4
XFILLER_12_113 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_4
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XFILLER_31_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_11 vpwr vgnd scs8hd_fill_2
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_63 vgnd vpwr scs8hd_decap_8
XFILLER_38_52 vgnd vpwr scs8hd_decap_8
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_171 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_230_ _230_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
X_161_ _152_/X _160_/X _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_21 vpwr vgnd scs8hd_fill_2
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_65 vgnd vpwr scs8hd_decap_3
XFILLER_1_14 vgnd vpwr scs8hd_decap_12
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_174 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_23 vgnd vpwr scs8hd_decap_8
XFILLER_19_21 vpwr vgnd scs8hd_fill_2
XFILLER_19_54 vgnd vpwr scs8hd_decap_4
XFILLER_19_98 vgnd vpwr scs8hd_decap_3
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _129_/X _145_/B _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XFILLER_33_133 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_122 vpwr vgnd scs8hd_fill_2
XFILLER_21_55 vpwr vgnd scs8hd_fill_2
XFILLER_30_169 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_144 vgnd vpwr scs8hd_decap_12
X_127_ _127_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_125 vgnd vpwr scs8hd_decap_12
XFILLER_16_22 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_4
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _186_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XANTENNA__130__C _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__A _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _204_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_56 vpwr vgnd scs8hd_fill_2
XFILLER_13_78 vgnd vpwr scs8hd_decap_4
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
Xmem_left_track_3.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__141__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_11 vgnd vpwr scs8hd_fill_1
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_160_ _121_/Y _114_/A _138_/Y _140_/D _160_/X vgnd vpwr scs8hd_or4_4
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_26 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _096_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_57 vgnd vpwr scs8hd_fill_1
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vgnd vpwr scs8hd_decap_4
XFILLER_42_156 vgnd vpwr scs8hd_decap_3
XFILLER_42_145 vgnd vpwr scs8hd_decap_8
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_98 vgnd vpwr scs8hd_fill_1
XFILLER_35_87 vpwr vgnd scs8hd_fill_2
XFILLER_35_43 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_4
XFILLER_35_21 vpwr vgnd scs8hd_fill_2
XFILLER_35_10 vpwr vgnd scs8hd_fill_2
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XFILLER_27_175 vgnd vpwr scs8hd_decap_6
X_143_ _118_/A _104_/B _143_/C _109_/A _145_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vgnd vpwr scs8hd_decap_3
XANTENNA__147__A _129_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_34 vgnd vpwr scs8hd_decap_4
XFILLER_21_78 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vgnd vpwr scs8hd_decap_12
XFILLER_7_58 vgnd vpwr scs8hd_decap_3
X_126_ _134_/A _104_/B _118_/C _109_/X _127_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_32_55 vgnd vpwr scs8hd_fill_1
XFILLER_12_137 vgnd vpwr scs8hd_decap_12
XFILLER_16_78 vpwr vgnd scs8hd_fill_2
XFILLER_32_77 vgnd vpwr scs8hd_fill_1
XANTENNA__144__B _145_/B vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _109_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XANTENNA__160__A _121_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _104_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_221 vgnd vpwr scs8hd_decap_12
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_39_195 vpwr vgnd scs8hd_fill_2
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_202 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_1_38 vgnd vpwr scs8hd_decap_12
XFILLER_36_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_69 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
XFILLER_35_66 vpwr vgnd scs8hd_fill_2
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _133_/A _141_/B _142_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XFILLER_33_179 vgnd vpwr scs8hd_decap_4
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _148_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_13 vpwr vgnd scs8hd_fill_2
XFILLER_15_168 vgnd vpwr scs8hd_decap_12
X_125_ _125_/A _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_26 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XFILLER_11_90 vgnd vpwr scs8hd_decap_3
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _152_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XFILLER_21_149 vgnd vpwr scs8hd_decap_4
XFILLER_29_205 vgnd vpwr scs8hd_decap_12
XFILLER_32_89 vgnd vpwr scs8hd_fill_1
XFILLER_12_149 vgnd vpwr scs8hd_decap_4
XFILLER_20_171 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
X_108_ address[1] enable _109_/A vgnd vpwr scs8hd_nand2_4
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
XFILLER_21_3 vgnd vpwr scs8hd_fill_1
XANTENNA__160__B _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_27_34 vpwr vgnd scs8hd_fill_2
XFILLER_40_200 vgnd vpwr scs8hd_decap_12
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_233 vgnd vpwr scs8hd_decap_8
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _109_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_47 vpwr vgnd scs8hd_fill_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XFILLER_38_44 vgnd vpwr scs8hd_decap_4
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_fill_1
XFILLER_14_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_133 vpwr vgnd scs8hd_fill_2
XFILLER_27_155 vpwr vgnd scs8hd_fill_2
XFILLER_27_188 vpwr vgnd scs8hd_fill_2
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _129_/X _141_/B _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _180_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_133 vpwr vgnd scs8hd_fill_2
XFILLER_33_169 vpwr vgnd scs8hd_fill_2
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_147 vgnd vpwr scs8hd_decap_6
XFILLER_24_169 vgnd vpwr scs8hd_decap_4
XFILLER_30_106 vgnd vpwr scs8hd_decap_3
X_124_ _127_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_139 vpwr vgnd scs8hd_fill_2
XFILLER_7_38 vgnd vpwr scs8hd_decap_12
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _157_/X vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_217 vgnd vpwr scs8hd_decap_12
XFILLER_12_106 vgnd vpwr scs8hd_fill_1
XFILLER_16_36 vgnd vpwr scs8hd_fill_1
XFILLER_20_183 vgnd vpwr scs8hd_decap_12
XFILLER_7_121 vgnd vpwr scs8hd_fill_1
X_107_ _125_/A _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__160__C _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__169__A _104_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_40_212 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA__171__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _184_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_39_175 vgnd vpwr scs8hd_decap_8
XFILLER_39_142 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _202_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_25 vgnd vpwr scs8hd_decap_4
XFILLER_24_36 vgnd vpwr scs8hd_decap_4
XFILLER_40_35 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_145 vpwr vgnd scs8hd_fill_2
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XFILLER_19_58 vgnd vpwr scs8hd_fill_1
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_fill_1
X_140_ _118_/A _104_/B _143_/C _140_/D _141_/B vgnd vpwr scs8hd_or4_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _188_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_112 vpwr vgnd scs8hd_fill_2
XFILLER_33_148 vpwr vgnd scs8hd_fill_2
XFILLER_33_115 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XANTENNA__163__C _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
XFILLER_32_170 vgnd vpwr scs8hd_decap_4
Xmem_top_track_6.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _206_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_123_ _134_/A _104_/B _118_/C _104_/D _125_/B vgnd vpwr scs8hd_or4_4
XFILLER_16_7 vpwr vgnd scs8hd_fill_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_229 vgnd vpwr scs8hd_decap_12
XFILLER_16_26 vgnd vpwr scs8hd_decap_4
XFILLER_16_48 vgnd vpwr scs8hd_decap_6
XFILLER_32_58 vgnd vpwr scs8hd_decap_3
XFILLER_32_47 vpwr vgnd scs8hd_fill_2
XFILLER_20_151 vpwr vgnd scs8hd_fill_2
XFILLER_20_195 vgnd vpwr scs8hd_decap_12
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
X_106_ address[0] _125_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XANTENNA__160__D _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_80 vpwr vgnd scs8hd_fill_2
XANTENNA__169__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_257 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_90 vpwr vgnd scs8hd_fill_2
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_5_72 vpwr vgnd scs8hd_fill_2
XFILLER_39_187 vpwr vgnd scs8hd_fill_2
XFILLER_39_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_40_47 vgnd vpwr scs8hd_decap_12
XFILLER_6_6 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_36_157 vpwr vgnd scs8hd_fill_2
XFILLER_36_102 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_7.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_102 vpwr vgnd scs8hd_fill_2
XFILLER_27_113 vpwr vgnd scs8hd_fill_2
XFILLER_42_116 vgnd vpwr scs8hd_decap_8
XFILLER_42_105 vpwr vgnd scs8hd_fill_2
XFILLER_33_105 vpwr vgnd scs8hd_fill_2
XFILLER_41_182 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_80 vpwr vgnd scs8hd_fill_2
XFILLER_26_190 vgnd vpwr scs8hd_decap_8
XFILLER_41_90 vgnd vpwr scs8hd_decap_4
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__163__D _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_3
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
X_122_ _121_/Y _134_/A vgnd vpwr scs8hd_buf_1
XFILLER_21_108 vpwr vgnd scs8hd_fill_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_32_15 vpwr vgnd scs8hd_fill_2
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
X_105_ _127_/A _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XANTENNA__169__C _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_200 vgnd vpwr scs8hd_decap_12
XFILLER_40_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_92 vgnd vpwr scs8hd_fill_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_28 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA__166__D _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_8
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_3
XFILLER_39_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_32_183 vgnd vpwr scs8hd_decap_8
XFILLER_24_139 vpwr vgnd scs8hd_fill_2
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_106 vpwr vgnd scs8hd_fill_2
X_121_ address[3] _121_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
XFILLER_23_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _178_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_109 vgnd vpwr scs8hd_fill_1
Xmem_top_track_2.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_120 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _118_/A _104_/B _118_/C _104_/D _105_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_6 vgnd vpwr scs8hd_decap_3
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_212 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_27_38 vpwr vgnd scs8hd_fill_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_48 vgnd vpwr scs8hd_fill_1
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_81 vgnd vpwr scs8hd_decap_4
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_30 vgnd vpwr scs8hd_decap_12
XFILLER_39_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _182_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_60 vgnd vpwr scs8hd_fill_1
XFILLER_36_115 vpwr vgnd scs8hd_fill_2
XFILLER_35_49 vgnd vpwr scs8hd_fill_1
XFILLER_27_137 vpwr vgnd scs8hd_fill_2
XFILLER_42_129 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_129 vpwr vgnd scs8hd_fill_2
XFILLER_33_118 vgnd vpwr scs8hd_decap_4
XPHY_60 vgnd vpwr scs8hd_decap_3
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _200_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_137 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_151 vgnd vpwr scs8hd_decap_6
XFILLER_41_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_93 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_140 vgnd vpwr scs8hd_decap_4
XFILLER_17_170 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _125_/A _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XFILLER_11_95 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _186_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XFILLER_16_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_143 vgnd vpwr scs8hd_decap_8
XFILLER_20_154 vgnd vpwr scs8hd_decap_3
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_22_61 vgnd vpwr scs8hd_decap_4
X_103_ _140_/D _104_/D vgnd vpwr scs8hd_buf_1
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _204_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_17 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_224 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_71 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_42 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_4
XFILLER_30_83 vgnd vpwr scs8hd_decap_3
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_149 vgnd vpwr scs8hd_decap_4
XFILLER_36_138 vgnd vpwr scs8hd_decap_4
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_160 vpwr vgnd scs8hd_fill_2
XFILLER_35_39 vpwr vgnd scs8hd_fill_2
XFILLER_35_28 vpwr vgnd scs8hd_fill_2
XFILLER_35_17 vpwr vgnd scs8hd_fill_2
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_116 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_174 vgnd vpwr scs8hd_decap_8
XFILLER_41_163 vpwr vgnd scs8hd_fill_2
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_15_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_23_141 vpwr vgnd scs8hd_fill_2
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vpwr vgnd scs8hd_fill_2
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_122 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
X_102_ address[1] _101_/Y _140_/D vgnd vpwr scs8hd_or2_4
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_8_86 vgnd vpwr scs8hd_decap_6
XFILLER_8_64 vgnd vpwr scs8hd_decap_8
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_236 vgnd vpwr scs8hd_decap_8
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XFILLER_38_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_5_87 vgnd vpwr scs8hd_decap_12
XFILLER_5_54 vgnd vpwr scs8hd_decap_6
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XFILLER_39_136 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_63 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_109 vgnd vpwr scs8hd_decap_6
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_120 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_42 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vgnd vpwr scs8hd_decap_4
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__107__A _125_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
XFILLER_32_19 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_13_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_105 vgnd vpwr scs8hd_decap_12
X_101_ enable _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_112 vgnd vpwr scs8hd_decap_8
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _176_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__104__B _104_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _198_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_38_29 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_99 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _180_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_63 vpwr vgnd scs8hd_fill_2
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_184 vpwr vgnd scs8hd_fill_2
XFILLER_35_173 vpwr vgnd scs8hd_fill_2
XFILLER_35_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vpwr vgnd scs8hd_fill_2
XFILLER_26_162 vpwr vgnd scs8hd_fill_2
XFILLER_26_173 vgnd vpwr scs8hd_decap_8
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_132 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_4
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_165 vpwr vgnd scs8hd_fill_2
XFILLER_23_176 vpwr vgnd scs8hd_fill_2
XFILLER_36_84 vgnd vpwr scs8hd_decap_8
XFILLER_36_73 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XFILLER_7_117 vgnd vpwr scs8hd_decap_4
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
X_100_ _100_/A _118_/C vgnd vpwr scs8hd_buf_1
XFILLER_34_205 vgnd vpwr scs8hd_decap_8
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
X_229_ _229_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _184_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_6.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__104__C _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_7 vgnd vpwr scs8hd_decap_4
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_208 vgnd vpwr scs8hd_decap_6
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _202_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_28_52 vgnd vpwr scs8hd_decap_12
XFILLER_28_85 vgnd vpwr scs8hd_fill_1
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XANTENNA__115__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_116 vgnd vpwr scs8hd_decap_4
XANTENNA__131__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_3
XFILLER_39_73 vpwr vgnd scs8hd_fill_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_4
XFILLER_36_119 vgnd vpwr scs8hd_decap_4
XFILLER_29_193 vgnd vpwr scs8hd_decap_12
XFILLER_29_171 vgnd vpwr scs8hd_decap_6
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A _134_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_111 vpwr vgnd scs8hd_fill_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_31 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_6
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
XFILLER_41_96 vgnd vpwr scs8hd_decap_4
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XFILLER_32_166 vpwr vgnd scs8hd_fill_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_6 vgnd vpwr scs8hd_decap_12
XFILLER_11_77 vpwr vgnd scs8hd_fill_2
XFILLER_36_52 vgnd vpwr scs8hd_fill_1
XFILLER_14_133 vgnd vpwr scs8hd_decap_12
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_6 vpwr vgnd scs8hd_fill_2
XANTENNA__123__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_22_21 vpwr vgnd scs8hd_fill_2
Xmem_top_track_12.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_6
XFILLER_8_23 vgnd vpwr scs8hd_decap_8
XFILLER_8_12 vgnd vpwr scs8hd_decap_8
X_159_ _155_/X _157_/X _159_/Y vgnd vpwr scs8hd_nor2_4
X_228_ _228_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vpwr vgnd scs8hd_fill_2
XFILLER_33_53 vgnd vpwr scs8hd_decap_3
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_209 vgnd vpwr scs8hd_decap_12
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__104__D _104_/D vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _118_/C vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _133_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_9_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_11 vgnd vpwr scs8hd_decap_3
XFILLER_14_99 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_150 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B _104_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_109 vpwr vgnd scs8hd_fill_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_76 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_41_167 vgnd vpwr scs8hd_decap_4
XFILLER_41_86 vpwr vgnd scs8hd_fill_2
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_145 vpwr vgnd scs8hd_fill_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_126 vgnd vpwr scs8hd_fill_1
XFILLER_20_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XANTENNA__118__C _118_/C vgnd vpwr scs8hd_diode_2
X_227_ _227_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
X_158_ _152_/X _157_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XFILLER_17_88 vgnd vpwr scs8hd_decap_4
XFILLER_17_99 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_65 vgnd vpwr scs8hd_decap_4
XFILLER_33_21 vgnd vpwr scs8hd_decap_4
XFILLER_33_10 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vgnd vpwr scs8hd_decap_4
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _174_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA__115__D _104_/D vgnd vpwr scs8hd_diode_2
XFILLER_39_107 vgnd vpwr scs8hd_decap_3
XFILLER_5_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_6 vgnd vpwr scs8hd_decap_6
Xmem_top_track_2.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _196_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_22 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_67 vpwr vgnd scs8hd_fill_2
XFILLER_39_42 vpwr vgnd scs8hd_fill_2
XFILLER_30_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _118_/C vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_143 vpwr vgnd scs8hd_fill_2
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XFILLER_26_121 vpwr vgnd scs8hd_fill_2
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_26_132 vpwr vgnd scs8hd_fill_2
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XPHY_55 vgnd vpwr scs8hd_decap_3
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_102 vpwr vgnd scs8hd_fill_2
XFILLER_32_146 vgnd vpwr scs8hd_decap_6
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _178_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vgnd vpwr scs8hd_fill_1
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
X_243_ _243_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_36_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _104_/D vgnd vpwr scs8hd_diode_2
XFILLER_37_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vpwr vgnd scs8hd_fill_2
XFILLER_28_205 vgnd vpwr scs8hd_decap_8
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_45 vpwr vgnd scs8hd_fill_2
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _134_/A address[2] _143_/C _109_/A _157_/X vgnd vpwr scs8hd_or4_4
XANTENNA__134__C _100_/A vgnd vpwr scs8hd_diode_2
X_226_ _226_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__118__D _109_/X vgnd vpwr scs8hd_diode_2
XANTENNA__150__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_17_34 vpwr vgnd scs8hd_fill_2
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_28_66 vpwr vgnd scs8hd_fill_2
XFILLER_28_88 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _182_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA__156__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_4
XFILLER_30_45 vpwr vgnd scs8hd_fill_2
XFILLER_14_46 vgnd vpwr scs8hd_decap_8
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_78 vgnd vpwr scs8hd_decap_3
XFILLER_30_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _200_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__D _109_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_188 vgnd vpwr scs8hd_decap_12
XFILLER_35_177 vgnd vpwr scs8hd_decap_6
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_26_100 vgnd vpwr scs8hd_fill_1
XFILLER_41_136 vgnd vpwr scs8hd_decap_4
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_66 vgnd vpwr scs8hd_fill_1
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_32_125 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_8
XFILLER_14_103 vgnd vpwr scs8hd_decap_4
X_242_ _242_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_239 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_139 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_12_90 vpwr vgnd scs8hd_fill_2
X_156_ _155_/X _156_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__D _109_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__B _160_/X vgnd vpwr scs8hd_diode_2
X_139_ _138_/Y _143_/C vgnd vpwr scs8hd_buf_1
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_91 vgnd vpwr scs8hd_decap_12
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_23 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_39_77 vpwr vgnd scs8hd_fill_2
XFILLER_39_66 vgnd vpwr scs8hd_fill_1
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_101 vpwr vgnd scs8hd_fill_2
XFILLER_35_156 vpwr vgnd scs8hd_fill_2
XANTENNA__167__A _166_/X vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
Xmem_left_track_13.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_13 vpwr vgnd scs8hd_fill_2
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XFILLER_41_115 vgnd vpwr scs8hd_decap_4
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_6
XFILLER_17_134 vgnd vpwr scs8hd_decap_12
XANTENNA__153__C _143_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_137 vpwr vgnd scs8hd_fill_2
XFILLER_36_12 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_67 vgnd vpwr scs8hd_decap_4
XFILLER_36_56 vgnd vpwr scs8hd_decap_8
XFILLER_36_23 vgnd vpwr scs8hd_decap_8
X_241_ _241_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
XFILLER_20_129 vgnd vpwr scs8hd_fill_1
XANTENNA__164__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_107 vgnd vpwr scs8hd_decap_3
XFILLER_22_25 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_240 vgnd vpwr scs8hd_decap_4
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
X_155_ address[0] _155_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_8
XFILLER_33_243 vgnd vpwr scs8hd_fill_1
XANTENNA__159__B _157_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
X_138_ address[4] _138_/B _138_/Y vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_34 vgnd vpwr scs8hd_decap_4
XFILLER_29_154 vpwr vgnd scs8hd_fill_2
XFILLER_29_132 vgnd vpwr scs8hd_decap_4
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_80 vpwr vgnd scs8hd_fill_2
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_36 vpwr vgnd scs8hd_fill_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
XFILLER_17_146 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _194_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_90 vgnd vpwr scs8hd_decap_3
XANTENNA__153__D _140_/D vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_116 vpwr vgnd scs8hd_fill_2
XFILLER_23_127 vgnd vpwr scs8hd_fill_1
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_149 vgnd vpwr scs8hd_decap_3
X_240_ _240_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_116 vgnd vpwr scs8hd_decap_8
X_171_ _109_/X _168_/B _155_/X _171_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _176_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
X_154_ _152_/X _156_/B _154_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _198_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XFILLER_33_36 vgnd vpwr scs8hd_fill_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
X_137_ address[5] _138_/B vgnd vpwr scs8hd_inv_8
XFILLER_23_80 vgnd vpwr scs8hd_decap_4
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vgnd vpwr scs8hd_decap_6
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_26 vgnd vpwr scs8hd_decap_4
XFILLER_39_46 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_136 vgnd vpwr scs8hd_decap_4
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_26_103 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_26_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_158 vgnd vpwr scs8hd_decap_12
XFILLER_40_183 vpwr vgnd scs8hd_fill_2
XFILLER_32_106 vpwr vgnd scs8hd_fill_2
XFILLER_25_191 vgnd vpwr scs8hd_decap_6
XFILLER_31_80 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_150 vgnd vpwr scs8hd_decap_3
XFILLER_22_161 vpwr vgnd scs8hd_fill_2
XFILLER_22_172 vgnd vpwr scs8hd_decap_12
X_170_ _109_/X _168_/B _152_/X _170_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XFILLER_9_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_109 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_49 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
X_153_ _134_/A address[2] _143_/C _140_/D _156_/B vgnd vpwr scs8hd_or4_4
XFILLER_26_8 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_17_16 vpwr vgnd scs8hd_fill_2
XFILLER_17_49 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
Xmem_left_track_5.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
X_136_ _133_/A _135_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_28_15 vpwr vgnd scs8hd_fill_2
XFILLER_28_26 vgnd vpwr scs8hd_decap_4
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_119_ _127_/A _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_12.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_145 vgnd vpwr scs8hd_decap_8
XFILLER_38_189 vgnd vpwr scs8hd_decap_12
XFILLER_38_178 vgnd vpwr scs8hd_decap_8
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_25 vpwr vgnd scs8hd_fill_2
XFILLER_30_49 vgnd vpwr scs8hd_decap_4
XFILLER_39_58 vgnd vpwr scs8hd_fill_1
XFILLER_29_167 vpwr vgnd scs8hd_fill_2
XFILLER_29_112 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_181 vgnd vpwr scs8hd_decap_12
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
XFILLER_40_140 vgnd vpwr scs8hd_decap_4
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_140 vpwr vgnd scs8hd_fill_2
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_151 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_17 vpwr vgnd scs8hd_fill_2
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
X_152_ _096_/A _152_/X vgnd vpwr scs8hd_buf_1
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_8 vpwr vgnd scs8hd_fill_2
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _129_/X _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_28_38 vgnd vpwr scs8hd_decap_3
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_82 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_3
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
X_118_ _118_/A _118_/B _118_/C _109_/X _119_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_135 vgnd vpwr scs8hd_fill_1
XFILLER_38_102 vpwr vgnd scs8hd_fill_2
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_17 vgnd vpwr scs8hd_decap_3
XFILLER_26_149 vgnd vpwr scs8hd_decap_4
XFILLER_41_119 vgnd vpwr scs8hd_fill_1
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_34_193 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_32_119 vgnd vpwr scs8hd_decap_4
XFILLER_40_163 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_163 vgnd vpwr scs8hd_decap_3
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_22_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_13_163 vgnd vpwr scs8hd_decap_12
XFILLER_26_82 vpwr vgnd scs8hd_fill_2
XFILLER_42_92 vgnd vpwr scs8hd_fill_1
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _192_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_73 vpwr vgnd scs8hd_fill_2
X_151_ _133_/A _149_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_203 vgnd vpwr scs8hd_decap_12
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_29 vgnd vpwr scs8hd_decap_3
XFILLER_33_39 vgnd vpwr scs8hd_decap_3
XFILLER_33_28 vgnd vpwr scs8hd_decap_8
XFILLER_33_17 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _174_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_72 vpwr vgnd scs8hd_fill_2
X_134_ _134_/A _118_/B _100_/A _109_/X _135_/B vgnd vpwr scs8hd_or4_4
XFILLER_0_10 vgnd vpwr scs8hd_decap_4
XFILLER_24_7 vpwr vgnd scs8hd_fill_2
XFILLER_0_21 vgnd vpwr scs8hd_decap_8
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _196_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_34_93 vgnd vpwr scs8hd_decap_3
X_117_ _125_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_125 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_3
Xmem_left_track_1.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_18 vpwr vgnd scs8hd_fill_2
XFILLER_39_38 vgnd vpwr scs8hd_fill_1
XFILLER_29_136 vgnd vpwr scs8hd_fill_1
XFILLER_37_191 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_51 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_29_82 vpwr vgnd scs8hd_fill_2
XFILLER_34_150 vgnd vpwr scs8hd_fill_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_117 vpwr vgnd scs8hd_fill_2
XFILLER_26_128 vpwr vgnd scs8hd_fill_2
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vpwr vgnd scs8hd_fill_2
XFILLER_40_175 vgnd vpwr scs8hd_decap_8
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_197 vgnd vpwr scs8hd_decap_12
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_31_153 vgnd vpwr scs8hd_decap_4
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_22_142 vgnd vpwr scs8hd_decap_8
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_175 vgnd vpwr scs8hd_decap_8
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _129_/X _149_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_60 vgnd vpwr scs8hd_fill_1
XFILLER_33_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_62 vgnd vpwr scs8hd_fill_1
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
X_133_ _133_/A _133_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_9_20 vpwr vgnd scs8hd_fill_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_116_ _127_/A _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_126 vgnd vpwr scs8hd_decap_4
XFILLER_20_63 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_50 vgnd vpwr scs8hd_decap_3
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_26_107 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_73 vgnd vpwr scs8hd_decap_4
XFILLER_31_51 vgnd vpwr scs8hd_decap_4
XANTENNA__102__B _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_132 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_165 vgnd vpwr scs8hd_decap_4
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_40 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_9_103 vgnd vpwr scs8hd_decap_12
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XFILLER_37_72 vpwr vgnd scs8hd_fill_2
XFILLER_33_227 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_30 vpwr vgnd scs8hd_fill_2
X_132_ address[0] _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA__110__B _104_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_43 vpwr vgnd scs8hd_fill_2
XFILLER_9_32 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_19 vgnd vpwr scs8hd_decap_4
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_63 vgnd vpwr scs8hd_decap_4
XFILLER_34_84 vgnd vpwr scs8hd_decap_8
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
X_115_ _118_/A _118_/B _118_/C _104_/D _116_/B vgnd vpwr scs8hd_or4_4
Xmem_left_track_9.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_29 vgnd vpwr scs8hd_decap_3
XFILLER_29_116 vgnd vpwr scs8hd_decap_4
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_4
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XFILLER_28_182 vpwr vgnd scs8hd_fill_2
XFILLER_28_193 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_188 vgnd vpwr scs8hd_decap_12
XFILLER_40_144 vgnd vpwr scs8hd_fill_1
XFILLER_15_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_152 vgnd vpwr scs8hd_decap_4
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_200 vpwr vgnd scs8hd_fill_2
.ends

