* NGSPICE file created from cbx_1__2_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

.subckt cbx_1__2_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] prog_clk
+ top_grid_pin_0_ vpwr vgnd
XFILLER_26_74 vgnd vpwr scs8hd_decap_12
XFILLER_13_166 vgnd vpwr scs8hd_decap_12
XFILLER_3_56 vgnd vpwr scs8hd_decap_12
XFILLER_35_280 vgnd vpwr scs8hd_decap_12
XFILLER_27_247 vgnd vpwr scs8hd_fill_1
XFILLER_33_239 vgnd vpwr scs8hd_decap_12
XFILLER_18_269 vgnd vpwr scs8hd_decap_12
XFILLER_12_98 vgnd vpwr scs8hd_decap_12
XFILLER_12_43 vgnd vpwr scs8hd_decap_12
XFILLER_10_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_239 vgnd vpwr scs8hd_decap_8
XFILLER_21_209 vgnd vpwr scs8hd_decap_4
XFILLER_2_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_31 vgnd vpwr scs8hd_decap_12
XFILLER_7_202 vgnd vpwr scs8hd_decap_12
XFILLER_29_117 vgnd vpwr scs8hd_decap_12
XFILLER_20_98 vgnd vpwr scs8hd_decap_12
XFILLER_20_43 vgnd vpwr scs8hd_decap_12
XFILLER_4_238 vgnd vpwr scs8hd_decap_6
XFILLER_15_87 vgnd vpwr scs8hd_decap_4
XFILLER_15_32 vgnd vpwr scs8hd_decap_12
XFILLER_31_178 vgnd vpwr scs8hd_decap_12
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_22_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_86 vgnd vpwr scs8hd_decap_12
XFILLER_13_178 vgnd vpwr scs8hd_decap_12
XFILLER_3_68 vgnd vpwr scs8hd_decap_12
XFILLER_9_105 vgnd vpwr scs8hd_decap_12
XFILLER_9_138 vgnd vpwr scs8hd_decap_12
XFILLER_27_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_182 vgnd vpwr scs8hd_fill_1
XFILLER_35_292 vgnd vpwr scs8hd_decap_6
XFILLER_12_55 vgnd vpwr scs8hd_decap_6
XFILLER_10_159 vgnd vpwr scs8hd_decap_12
XFILLER_26_281 vgnd vpwr scs8hd_decap_12
XFILLER_23_251 vgnd vpwr scs8hd_decap_12
XFILLER_23_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_86 vgnd vpwr scs8hd_decap_12
XFILLER_18_43 vgnd vpwr scs8hd_decap_12
XFILLER_11_276 vgnd vpwr scs8hd_decap_12
XFILLER_7_247 vgnd vpwr scs8hd_fill_1
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
XFILLER_29_129 vgnd vpwr scs8hd_decap_12
XFILLER_20_55 vgnd vpwr scs8hd_decap_6
XFILLER_34_110 vgnd vpwr scs8hd_decap_12
XFILLER_28_184 vgnd vpwr scs8hd_decap_12
XFILLER_25_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_66 vpwr vgnd scs8hd_fill_2
XFILLER_15_44 vgnd vpwr scs8hd_decap_12
XFILLER_15_11 vpwr vgnd scs8hd_fill_2
XFILLER_31_32 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_253 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_22_135 vgnd vpwr scs8hd_decap_12
XFILLER_26_98 vgnd vpwr scs8hd_decap_12
XFILLER_21_190 vgnd vpwr scs8hd_decap_8
XFILLER_9_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_205 vgnd vpwr scs8hd_decap_8
XFILLER_26_293 vgnd vpwr scs8hd_decap_6
XFILLER_24_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_296 vgnd vpwr scs8hd_decap_3
XFILLER_23_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_55 vgnd vpwr scs8hd_decap_6
XFILLER_11_288 vgnd vpwr scs8hd_decap_8
XFILLER_7_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S mux_bottom_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_281 vgnd vpwr scs8hd_decap_12
XFILLER_1_80 vgnd vpwr scs8hd_decap_12
XFILLER_29_87 vgnd vpwr scs8hd_decap_4
XFILLER_29_32 vgnd vpwr scs8hd_decap_12
XFILLER_28_196 vgnd vpwr scs8hd_decap_12
XFILLER_19_141 vpwr vgnd scs8hd_fill_2
XFILLER_31_44 vgnd vpwr scs8hd_decap_12
XFILLER_25_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_56 vgnd vpwr scs8hd_decap_8
XANTENNA__04__A chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_0_298 vgnd vpwr scs8hd_fill_1
XFILLER_0_265 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_147 vgnd vpwr scs8hd_decap_12
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_129 vgnd vpwr scs8hd_fill_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_261 vgnd vpwr scs8hd_decap_12
XFILLER_27_239 vgnd vpwr scs8hd_decap_8
XFILLER_5_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_56 vgnd vpwr scs8hd_decap_12
XANTENNA__12__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_2_135 vgnd vpwr scs8hd_decap_12
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_190 vgnd vpwr scs8hd_decap_12
XFILLER_20_245 vgnd vpwr scs8hd_decap_12
XANTENNA__07__A chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_11_256 vgnd vpwr scs8hd_decap_12
XFILLER_11_245 vgnd vpwr scs8hd_fill_1
XFILLER_7_227 vgnd vpwr scs8hd_decap_12
X_29_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_4_208 vpwr vgnd scs8hd_fill_2
XFILLER_6_293 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_252 vpwr vgnd scs8hd_fill_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_37 vgnd vpwr scs8hd_decap_12
XFILLER_34_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_7 vgnd vpwr scs8hd_decap_12
XFILLER_3_274 vgnd vpwr scs8hd_fill_1
XFILLER_3_296 vgnd vpwr scs8hd_decap_3
XFILLER_31_56 vgnd vpwr scs8hd_decap_12
XFILLER_25_178 vgnd vpwr scs8hd_decap_12
XANTENNA__20__A chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_0_277 vpwr vgnd scs8hd_fill_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_123 vgnd vpwr scs8hd_decap_12
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_159 vgnd vpwr scs8hd_decap_12
XFILLER_7_80 vgnd vpwr scs8hd_decap_12
XANTENNA__15__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_4
XFILLER_35_273 vgnd vpwr scs8hd_decap_6
XFILLER_8_152 vgnd vpwr scs8hd_decap_12
XFILLER_8_196 vgnd vpwr scs8hd_decap_12
XFILLER_5_133 vpwr vgnd scs8hd_fill_2
XFILLER_32_232 vgnd vpwr scs8hd_decap_12
XFILLER_5_166 vgnd vpwr scs8hd_decap_12
XFILLER_23_276 vgnd vpwr scs8hd_decap_12
XFILLER_23_68 vgnd vpwr scs8hd_decap_12
XFILLER_2_147 vgnd vpwr scs8hd_decap_12
XFILLER_14_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_257 vgnd vpwr scs8hd_decap_12
XFILLER_11_268 vgnd vpwr scs8hd_decap_6
XANTENNA__23__A chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_11_202 vgnd vpwr scs8hd_decap_12
XFILLER_7_239 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_ipin_0.mux_l3_in_1_/S ccff_tail
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_93 vgnd vpwr scs8hd_decap_12
X_28_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__18__A chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_29_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_110 vgnd vpwr scs8hd_decap_12
XFILLER_34_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_198 vpwr vgnd scs8hd_fill_2
XFILLER_19_154 vgnd vpwr scs8hd_decap_12
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_6
XFILLER_6_49 vgnd vpwr scs8hd_decap_12
XFILLER_33_190 vgnd vpwr scs8hd_decap_12
XFILLER_31_68 vgnd vpwr scs8hd_decap_12
XFILLER_31_105 vgnd vpwr scs8hd_decap_12
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_135 vgnd vpwr scs8hd_decap_12
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_182 vgnd vpwr scs8hd_fill_1
XFILLER_15_190 vgnd vpwr scs8hd_decap_12
XFILLER_13_105 vgnd vpwr scs8hd_decap_12
XANTENNA__31__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_12
XFILLER_12_171 vgnd vpwr scs8hd_decap_12
XFILLER_8_164 vgnd vpwr scs8hd_decap_12
XFILLER_18_208 vgnd vpwr scs8hd_decap_12
XANTENNA__26__A chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_17_296 vgnd vpwr scs8hd_decap_3
XFILLER_17_274 vgnd vpwr scs8hd_fill_1
XFILLER_17_252 vpwr vgnd scs8hd_fill_2
XFILLER_5_178 vgnd vpwr scs8hd_decap_12
XFILLER_23_288 vgnd vpwr scs8hd_decap_8
XFILLER_23_211 vgnd vpwr scs8hd_decap_3
XFILLER_13_80 vgnd vpwr scs8hd_decap_12
XFILLER_2_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_269 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S mux_bottom_ipin_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_ipin_0.mux_l2_in_2_/S mux_bottom_ipin_0.mux_l3_in_1_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
X_27_ chanx_right_in[9] chanx_left_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_29_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_147 vgnd vpwr scs8hd_decap_12
XFILLER_19_166 vgnd vpwr scs8hd_decap_12
XANTENNA__34__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_276 vgnd vpwr scs8hd_decap_12
XFILLER_25_136 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_117 vgnd vpwr scs8hd_decap_12
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_80 vgnd vpwr scs8hd_decap_12
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_147 vgnd vpwr scs8hd_decap_12
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_257 vgnd vpwr scs8hd_decap_4
XANTENNA__29__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D mux_bottom_ipin_0.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_110 vgnd vpwr scs8hd_decap_12
XFILLER_8_176 vgnd vpwr scs8hd_decap_6
XFILLER_35_242 vgnd vpwr scs8hd_decap_6
XFILLER_32_245 vgnd vpwr scs8hd_decap_12
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA__37__A chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_14_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_11_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_ipin_0.mux_l1_in_2_/S mux_bottom_ipin_0.mux_l2_in_2_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_24_91 vgnd vpwr scs8hd_decap_12
XFILLER_28_123 vgnd vpwr scs8hd_decap_12
X_26_ chanx_right_in[10] chanx_left_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_19_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_145 vgnd vpwr scs8hd_decap_8
XFILLER_19_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0 mux_bottom_ipin_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_288 vgnd vpwr scs8hd_decap_8
XFILLER_34_159 vgnd vpwr scs8hd_decap_12
XFILLER_25_148 vgnd vpwr scs8hd_decap_4
XFILLER_15_27 vgnd vpwr scs8hd_decap_4
X_09_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_31_129 vgnd vpwr scs8hd_decap_12
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_192 vpwr vgnd scs8hd_fill_2
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_159 vgnd vpwr scs8hd_decap_12
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_269 vgnd vpwr scs8hd_decap_8
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_184 vgnd vpwr scs8hd_decap_12
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_26_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_129 vgnd vpwr scs8hd_decap_12
XFILLER_29_262 vgnd vpwr scs8hd_decap_12
XFILLER_16_81 vgnd vpwr scs8hd_decap_12
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_12_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_298 vgnd vpwr scs8hd_fill_1
XFILLER_32_257 vgnd vpwr scs8hd_decap_12
XFILLER_27_80 vgnd vpwr scs8hd_decap_12
XFILLER_17_276 vgnd vpwr scs8hd_decap_12
XFILLER_4_51 vgnd vpwr scs8hd_decap_8
XFILLER_4_62 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_205 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_250 vgnd vpwr scs8hd_decap_12
XFILLER_34_59 vpwr vgnd scs8hd_fill_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_227 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_bottom_ipin_0.mux_l1_in_2_/S
+ mem_bottom_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_220 vgnd vpwr scs8hd_decap_12
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
X_25_ chanx_right_in[11] chanx_left_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_28_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1 mux_bottom_ipin_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_212 vpwr vgnd scs8hd_fill_2
XFILLER_3_223 vgnd vpwr scs8hd_decap_12
XFILLER_3_256 vgnd vpwr scs8hd_decap_12
XFILLER_25_105 vgnd vpwr scs8hd_decap_12
X_08_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_171 vgnd vpwr scs8hd_decap_12
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_93 vgnd vpwr scs8hd_decap_12
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_7 vgnd vpwr scs8hd_decap_12
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_196 vgnd vpwr scs8hd_decap_12
XFILLER_30_174 vgnd vpwr scs8hd_decap_8
XFILLER_26_27 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vgnd vpwr scs8hd_decap_12
XFILLER_29_296 vgnd vpwr scs8hd_decap_3
XFILLER_29_274 vgnd vpwr scs8hd_fill_1
XFILLER_29_252 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_196 vgnd vpwr scs8hd_decap_12
XFILLER_8_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XFILLER_26_200 vgnd vpwr scs8hd_decap_12
XFILLER_5_137 vgnd vpwr scs8hd_decap_12
XFILLER_32_269 vgnd vpwr scs8hd_decap_12
XFILLER_17_288 vgnd vpwr scs8hd_decap_8
XFILLER_4_74 vgnd vpwr scs8hd_decap_12
XFILLER_4_181 vpwr vgnd scs8hd_fill_2
XFILLER_23_203 vgnd vpwr scs8hd_decap_8
XFILLER_14_269 vgnd vpwr scs8hd_decap_12
X_41_ chanx_left_in[15] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_12
XFILLER_20_217 vgnd vpwr scs8hd_decap_12
XFILLER_11_239 vgnd vpwr scs8hd_decap_6
XFILLER_9_262 vgnd vpwr scs8hd_decap_12
X_24_ chanx_right_in[12] chanx_left_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_6_232 vgnd vpwr scs8hd_decap_12
XFILLER_29_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_147 vgnd vpwr scs8hd_decap_12
XFILLER_10_62 vgnd vpwr scs8hd_decap_12
XFILLER_10_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_235 vgnd vpwr scs8hd_decap_12
XFILLER_3_268 vgnd vpwr scs8hd_decap_6
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_27_180 vpwr vgnd scs8hd_fill_2
XFILLER_19_93 vgnd vpwr scs8hd_decap_12
XFILLER_25_117 vgnd vpwr scs8hd_decap_12
X_07_ chanx_left_in[9] chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_120 vpwr vgnd scs8hd_fill_2
XFILLER_26_39 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_12_19 vgnd vpwr scs8hd_decap_12
XFILLER_8_135 vgnd vpwr scs8hd_decap_12
XFILLER_26_245 vgnd vpwr scs8hd_decap_12
XFILLER_26_212 vgnd vpwr scs8hd_decap_12
XFILLER_5_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_149 vgnd vpwr scs8hd_decap_4
XFILLER_7_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_93 vgnd vpwr scs8hd_decap_12
XFILLER_17_256 vgnd vpwr scs8hd_decap_12
XFILLER_23_215 vgnd vpwr scs8hd_decap_12
XFILLER_4_86 vgnd vpwr scs8hd_decap_12
X_40_ chanx_left_in[16] chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_1_141 vgnd vpwr scs8hd_decap_12
XFILLER_20_229 vgnd vpwr scs8hd_decap_12
XFILLER_9_296 vgnd vpwr scs8hd_decap_3
XFILLER_9_274 vgnd vpwr scs8hd_fill_1
XFILLER_34_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0 _01_/HI vgnd vpwr scs8hd_diode_2
X_23_ chanx_right_in[13] chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_1_32 vgnd vpwr scs8hd_decap_12
XFILLER_28_159 vgnd vpwr scs8hd_decap_12
XFILLER_20_19 vgnd vpwr scs8hd_decap_12
XFILLER_19_137 vpwr vgnd scs8hd_fill_2
XFILLER_10_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_247 vgnd vpwr scs8hd_fill_1
XFILLER_25_129 vgnd vpwr scs8hd_fill_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_06_ chanx_left_in[10] chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_24_184 vgnd vpwr scs8hd_decap_8
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_29_276 vgnd vpwr scs8hd_decap_12
XFILLER_29_210 vpwr vgnd scs8hd_fill_2
XFILLER_21_198 vgnd vpwr scs8hd_fill_1
XFILLER_21_154 vgnd vpwr scs8hd_decap_12
XFILLER_16_62 vgnd vpwr scs8hd_decap_8
XFILLER_12_110 vgnd vpwr scs8hd_decap_12
XFILLER_8_147 vgnd vpwr scs8hd_fill_1
XFILLER_26_257 vgnd vpwr scs8hd_decap_12
XFILLER_26_224 vgnd vpwr scs8hd_decap_12
XFILLER_17_268 vgnd vpwr scs8hd_decap_6
XFILLER_17_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_117 vgnd vpwr scs8hd_decap_8
XFILLER_23_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_161 vgnd vpwr scs8hd_decap_12
XFILLER_18_19 vgnd vpwr scs8hd_decap_12
XFILLER_24_62 vgnd vpwr scs8hd_decap_3
XFILLER_24_51 vgnd vpwr scs8hd_decap_8
X_22_ chanx_right_in[14] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_10_296 vgnd vpwr scs8hd_decap_3
XFILLER_10_252 vgnd vpwr scs8hd_decap_12
XFILLER_1_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_11 vgnd vpwr scs8hd_decap_12
XFILLER_6_245 vgnd vpwr scs8hd_decap_12
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
XFILLER_27_193 vgnd vpwr scs8hd_decap_12
XFILLER_19_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_141 vgnd vpwr scs8hd_decap_12
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
X_05_ chanx_left_in[11] chanx_right_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_24_196 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_100 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_15_141 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_32 vgnd vpwr scs8hd_decap_12
XFILLER_21_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_62 vgnd vpwr scs8hd_decap_12
XFILLER_32_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_288 vgnd vpwr scs8hd_decap_8
XFILLER_26_269 vgnd vpwr scs8hd_decap_12
XFILLER_26_236 vgnd vpwr scs8hd_decap_8
XFILLER_17_247 vgnd vpwr scs8hd_fill_1
XFILLER_5_129 vpwr vgnd scs8hd_fill_2
XFILLER_23_239 vgnd vpwr scs8hd_decap_12
XFILLER_4_173 vgnd vpwr scs8hd_decap_8
XFILLER_4_184 vgnd vpwr scs8hd_decap_12
XFILLER_9_276 vgnd vpwr scs8hd_decap_12
XFILLER_1_154 vgnd vpwr scs8hd_decap_12
X_21_ chanx_right_in[15] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_10_264 vgnd vpwr scs8hd_decap_12
XFILLER_10_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_23 vgnd vpwr scs8hd_decap_8
XFILLER_6_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_117 vgnd vpwr scs8hd_decap_12
XFILLER_10_98 vgnd vpwr scs8hd_decap_12
X_04_ chanx_left_in[12] chanx_right_out[12] vgnd vpwr scs8hd_buf_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_123 vgnd vpwr scs8hd_decap_12
XFILLER_30_112 vgnd vpwr scs8hd_decap_8
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_7_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_178 vgnd vpwr scs8hd_decap_12
XFILLER_32_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_256 vgnd vpwr scs8hd_decap_4
XFILLER_29_245 vgnd vpwr scs8hd_fill_1
XFILLER_16_31 vgnd vpwr scs8hd_decap_12
XFILLER_12_123 vgnd vpwr scs8hd_decap_12
XFILLER_34_281 vgnd vpwr scs8hd_decap_12
XFILLER_17_215 vgnd vpwr scs8hd_decap_12
XFILLER_4_196 vgnd vpwr scs8hd_decap_12
XFILLER_13_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_288 vgnd vpwr scs8hd_decap_8
XFILLER_10_276 vgnd vpwr scs8hd_decap_12
XFILLER_10_232 vgnd vpwr scs8hd_decap_12
XFILLER_6_269 vgnd vpwr scs8hd_decap_12
X_20_ chanx_right_in[16] chanx_left_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_1_68 vgnd vpwr scs8hd_decap_12
XFILLER_19_129 vgnd vpwr scs8hd_decap_6
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_18_151 vgnd vpwr scs8hd_decap_12
X_03_ chanx_left_in[13] chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_33_154 vgnd vpwr scs8hd_decap_12
XFILLER_24_121 vgnd vpwr scs8hd_fill_1
XFILLER_18_184 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_135 vgnd vpwr scs8hd_decap_12
XFILLER_21_32 vgnd vpwr scs8hd_decap_12
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_154 vgnd vpwr scs8hd_decap_12
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_7_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_86 vgnd vpwr scs8hd_decap_12
XFILLER_16_43 vgnd vpwr scs8hd_decap_12
XFILLER_12_135 vgnd vpwr scs8hd_decap_12
XFILLER_35_249 vgnd vpwr scs8hd_decap_12
XFILLER_11_190 vgnd vpwr scs8hd_decap_12
XFILLER_7_150 vgnd vpwr scs8hd_decap_3
XFILLER_34_293 vgnd vpwr scs8hd_decap_6
XFILLER_32_208 vgnd vpwr scs8hd_decap_12
XFILLER_17_227 vgnd vpwr scs8hd_decap_12
XFILLER_31_296 vgnd vpwr scs8hd_decap_3
XFILLER_31_274 vgnd vpwr scs8hd_fill_1
XFILLER_31_252 vpwr vgnd scs8hd_fill_2
XFILLER_22_296 vgnd vpwr scs8hd_decap_3
XFILLER_22_252 vgnd vpwr scs8hd_decap_12
XFILLER_14_208 vgnd vpwr scs8hd_decap_12
XFILLER_13_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_11 vpwr vgnd scs8hd_fill_2
XFILLER_1_178 vgnd vpwr scs8hd_decap_12
XFILLER_13_296 vgnd vpwr scs8hd_decap_3
XFILLER_13_274 vgnd vpwr scs8hd_fill_1
XFILLER_13_252 vpwr vgnd scs8hd_fill_2
XFILLER_9_234 vpwr vgnd scs8hd_fill_2
XFILLER_10_288 vgnd vpwr scs8hd_decap_8
XFILLER_3_207 vgnd vpwr scs8hd_decap_3
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
XFILLER_27_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_32 vgnd vpwr scs8hd_decap_12
XFILLER_33_166 vgnd vpwr scs8hd_decap_12
XFILLER_18_196 vgnd vpwr scs8hd_decap_12
XFILLER_18_163 vgnd vpwr scs8hd_decap_12
X_02_ chanx_left_in[14] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_21_44 vgnd vpwr scs8hd_decap_12
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_147 vgnd vpwr scs8hd_decap_8
XFILLER_15_166 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_68 vgnd vpwr scs8hd_decap_12
XFILLER_16_55 vgnd vpwr scs8hd_decap_6
XFILLER_12_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_98 vgnd vpwr scs8hd_decap_12
XFILLER_20_180 vgnd vpwr scs8hd_decap_3
XFILLER_27_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_239 vgnd vpwr scs8hd_decap_8
XFILLER_4_110 vgnd vpwr scs8hd_decap_12
XFILLER_22_264 vgnd vpwr scs8hd_decap_12
XFILLER_22_220 vgnd vpwr scs8hd_decap_12
XFILLER_13_56 vgnd vpwr scs8hd_decap_12
XANTENNA__02__A chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_9_246 vpwr vgnd scs8hd_fill_2
XFILLER_10_245 vgnd vpwr scs8hd_decap_3
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_11 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S mux_bottom_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_219 vpwr vgnd scs8hd_fill_2
XFILLER_33_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_01_ _01_/HI _01_/LO vgnd vpwr scs8hd_conb_1
XFILLER_18_175 vgnd vpwr scs8hd_decap_8
XFILLER_18_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_252 vgnd vpwr scs8hd_decap_12
XFILLER_2_296 vgnd vpwr scs8hd_decap_3
XFILLER_24_123 vgnd vpwr scs8hd_decap_12
XFILLER_21_56 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__10__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_178 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_29_215 vgnd vpwr scs8hd_decap_12
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_159 vgnd vpwr scs8hd_decap_12
XANTENNA__05__A chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_7_141 vgnd vpwr scs8hd_decap_6
XFILLER_27_44 vgnd vpwr scs8hd_decap_12
XFILLER_31_276 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_59 vpwr vgnd scs8hd_fill_2
XFILLER_4_155 vpwr vgnd scs8hd_fill_2
XFILLER_22_276 vgnd vpwr scs8hd_decap_12
XFILLER_22_232 vgnd vpwr scs8hd_decap_12
XFILLER_13_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_276 vgnd vpwr scs8hd_decap_12
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_24_67 vgnd vpwr scs8hd_decap_12
XANTENNA__13__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
XFILLER_27_154 vgnd vpwr scs8hd_decap_12
XFILLER_19_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_23 vgnd vpwr scs8hd_decap_8
XANTENNA__08__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_2_220 vgnd vpwr scs8hd_decap_12
XFILLER_2_264 vgnd vpwr scs8hd_decap_12
XFILLER_24_135 vgnd vpwr scs8hd_decap_12
XFILLER_21_68 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_190 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_227 vgnd vpwr scs8hd_decap_12
XFILLER_21_105 vgnd vpwr scs8hd_decap_12
XANTENNA__21__A chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_27_56 vgnd vpwr scs8hd_decap_12
XFILLER_25_296 vgnd vpwr scs8hd_decap_3
XFILLER_25_274 vgnd vpwr scs8hd_fill_1
XFILLER_25_252 vpwr vgnd scs8hd_fill_2
XANTENNA__16__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_31_288 vgnd vpwr scs8hd_decap_8
XFILLER_16_296 vgnd vpwr scs8hd_decap_3
XFILLER_16_252 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_12
XFILLER_4_123 vgnd vpwr scs8hd_decap_12
XFILLER_22_288 vgnd vpwr scs8hd_decap_8
XFILLER_13_288 vgnd vpwr scs8hd_decap_8
XFILLER_9_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_79 vgnd vpwr scs8hd_decap_12
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_27_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_68 vgnd vpwr scs8hd_decap_12
XFILLER_10_59 vpwr vgnd scs8hd_fill_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XANTENNA__24__A chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_2_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XFILLER_24_147 vgnd vpwr scs8hd_decap_12
XFILLER_24_103 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__19__A chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_117 vgnd vpwr scs8hd_decap_12
XFILLER_11_80 vgnd vpwr scs8hd_decap_12
XFILLER_29_239 vgnd vpwr scs8hd_decap_6
XFILLER_7_154 vgnd vpwr scs8hd_decap_12
XFILLER_34_220 vgnd vpwr scs8hd_decap_12
XFILLER_27_68 vgnd vpwr scs8hd_decap_12
XFILLER_16_264 vgnd vpwr scs8hd_decap_12
XFILLER_16_220 vgnd vpwr scs8hd_decap_12
XANTENNA__32__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_39 vgnd vpwr scs8hd_decap_12
XFILLER_4_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_256 vgnd vpwr scs8hd_decap_12
XFILLER_22_245 vgnd vpwr scs8hd_decap_3
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_256 vgnd vpwr scs8hd_decap_12
XFILLER_9_238 vgnd vpwr scs8hd_decap_8
XFILLER_9_227 vgnd vpwr scs8hd_decap_3
XFILLER_1_105 vgnd vpwr scs8hd_decap_12
XANTENNA__27__A chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_decap_12
XFILLER_5_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_208 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_252 vpwr vgnd scs8hd_fill_2
XFILLER_5_274 vgnd vpwr scs8hd_fill_1
XFILLER_5_296 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S mux_bottom_ipin_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_123 vgnd vpwr scs8hd_decap_6
XANTENNA__40__A chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_2_288 vgnd vpwr scs8hd_decap_8
XFILLER_24_159 vgnd vpwr scs8hd_decap_12
XFILLER_24_115 vgnd vpwr scs8hd_decap_6
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XANTENNA__35__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_21_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_7 vgnd vpwr scs8hd_decap_12
XFILLER_20_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_166 vgnd vpwr scs8hd_decap_12
XFILLER_34_232 vgnd vpwr scs8hd_decap_12
XFILLER_25_276 vgnd vpwr scs8hd_decap_12
XFILLER_4_147 vgnd vpwr scs8hd_decap_8
XFILLER_31_268 vgnd vpwr scs8hd_decap_6
XFILLER_31_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D mux_bottom_ipin_0.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_80 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_decap_12
XFILLER_16_232 vgnd vpwr scs8hd_decap_12
XFILLER_13_202 vgnd vpwr scs8hd_decap_12
XFILLER_13_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_268 vgnd vpwr scs8hd_decap_6
XFILLER_24_59 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_72 vgnd vpwr scs8hd_decap_12
XANTENNA__38__A chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_14_92 vgnd vpwr scs8hd_decap_12
XFILLER_30_80 vgnd vpwr scs8hd_fill_1
XFILLER_10_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_245 vgnd vpwr scs8hd_decap_3
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_105 vgnd vpwr scs8hd_decap_12
XFILLER_2_51 vgnd vpwr scs8hd_decap_8
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_62 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_171 vgnd vpwr scs8hd_decap_12
XFILLER_21_27 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l2_in_3_ _01_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_2_/S
+ mux_bottom_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_190 vgnd vpwr scs8hd_decap_12
XFILLER_15_105 vgnd vpwr scs8hd_decap_12
XFILLER_11_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_171 vgnd vpwr scs8hd_decap_12
XFILLER_32_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_296 vgnd vpwr scs8hd_decap_3
XFILLER_28_252 vgnd vpwr scs8hd_decap_12
XFILLER_11_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_296 vgnd vpwr scs8hd_decap_3
XFILLER_19_274 vgnd vpwr scs8hd_fill_1
XFILLER_19_230 vgnd vpwr scs8hd_decap_12
XFILLER_7_178 vgnd vpwr scs8hd_decap_12
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_288 vgnd vpwr scs8hd_decap_8
XFILLER_33_80 vgnd vpwr scs8hd_decap_12
XFILLER_31_247 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ ccff_tail mux_bottom_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_288 vgnd vpwr scs8hd_decap_8
XFILLER_1_129 vgnd vpwr scs8hd_decap_12
XFILLER_13_247 vgnd vpwr scs8hd_fill_1
XFILLER_24_27 vgnd vpwr scs8hd_decap_12
XFILLER_5_84 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_276 vgnd vpwr scs8hd_decap_12
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_33_117 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_2_/S
+ mux_bottom_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_74 vgnd vpwr scs8hd_decap_12
XFILLER_15_117 vgnd vpwr scs8hd_decap_12
X_39_ chanx_left_in[17] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_264 vgnd vpwr scs8hd_decap_12
XFILLER_28_220 vgnd vpwr scs8hd_decap_12
XFILLER_34_245 vgnd vpwr scs8hd_decap_12
XFILLER_19_242 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S mux_bottom_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_256 vgnd vpwr scs8hd_decap_12
XFILLER_8_62 vgnd vpwr scs8hd_decap_12
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_93 vgnd vpwr scs8hd_decap_12
XFILLER_16_245 vgnd vpwr scs8hd_decap_3
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_13_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_6
XFILLER_8_252 vgnd vpwr scs8hd_decap_12
XFILLER_8_296 vgnd vpwr scs8hd_decap_3
XFILLER_24_39 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_5_288 vgnd vpwr scs8hd_decap_8
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_129 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_181 vpwr vgnd scs8hd_fill_2
XFILLER_25_93 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_184 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_2_/S mux_bottom_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0 mux_bottom_ipin_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_129 vgnd vpwr scs8hd_decap_12
XFILLER_14_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_39 vgnd vpwr scs8hd_decap_12
X_38_ chanx_left_in[18] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_28_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_110 vgnd vpwr scs8hd_decap_12
XFILLER_34_257 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_decap_12
XFILLER_19_276 vgnd vpwr scs8hd_decap_12
XFILLER_19_254 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_7 vgnd vpwr scs8hd_decap_12
XFILLER_11_154 vgnd vpwr scs8hd_decap_12
XFILLER_7_147 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0 mux_bottom_ipin_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_268 vgnd vpwr scs8hd_decap_6
XFILLER_25_202 vgnd vpwr scs8hd_decap_12
XFILLER_6_180 vgnd vpwr scs8hd_decap_3
XFILLER_8_74 vgnd vpwr scs8hd_decap_12
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_93 vgnd vpwr scs8hd_decap_12
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_227 vgnd vpwr scs8hd_decap_12
XFILLER_3_183 vgnd vpwr scs8hd_decap_12
XFILLER_13_227 vgnd vpwr scs8hd_decap_12
XFILLER_8_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_264 vgnd vpwr scs8hd_decap_12
XFILLER_10_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_14_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_256 vgnd vpwr scs8hd_decap_12
XFILLER_27_105 vgnd vpwr scs8hd_decap_12
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_2_/S mux_bottom_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_98 vgnd vpwr scs8hd_decap_12
XFILLER_23_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1 mux_bottom_ipin_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
X_37_ chanx_left_in[19] chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_20_144 vgnd vpwr scs8hd_decap_12
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
XFILLER_28_288 vgnd vpwr scs8hd_decap_8
XFILLER_22_62 vgnd vpwr scs8hd_decap_12
XFILLER_22_51 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_166 vgnd vpwr scs8hd_decap_12
XFILLER_34_269 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1 mux_bottom_ipin_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_288 vgnd vpwr scs8hd_decap_8
XFILLER_19_266 vgnd vpwr scs8hd_decap_8
XFILLER_8_86 vgnd vpwr scs8hd_decap_12
XFILLER_25_247 vgnd vpwr scs8hd_fill_1
XFILLER_17_84 vgnd vpwr scs8hd_decap_8
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_239 vgnd vpwr scs8hd_decap_8
XFILLER_3_195 vgnd vpwr scs8hd_decap_12
XFILLER_21_250 vgnd vpwr scs8hd_decap_12
XFILLER_13_239 vgnd vpwr scs8hd_decap_8
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_decap_12
XFILLER_5_32 vpwr vgnd scs8hd_fill_2
XFILLER_30_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_268 vgnd vpwr scs8hd_decap_6
XFILLER_27_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_139 vgnd vpwr scs8hd_decap_12
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_161 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_84 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_fill_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_156 vgnd vpwr scs8hd_decap_12
XFILLER_20_123 vgnd vpwr scs8hd_decap_12
X_36_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_28_245 vgnd vpwr scs8hd_decap_3
XFILLER_22_74 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_2_/S
+ mux_bottom_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_105 vgnd vpwr scs8hd_decap_12
XFILLER_8_98 vgnd vpwr scs8hd_decap_12
XFILLER_25_215 vgnd vpwr scs8hd_decap_12
X_19_ chanx_right_in[17] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_281 vgnd vpwr scs8hd_decap_12
XFILLER_3_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_262 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_288 vgnd vpwr scs8hd_decap_8
XFILLER_30_74 vgnd vpwr scs8hd_decap_6
XFILLER_14_31 vgnd vpwr scs8hd_decap_12
XFILLER_5_247 vgnd vpwr scs8hd_fill_1
XFILLER_27_129 vgnd vpwr scs8hd_decap_12
XPHY_63 vgnd vpwr scs8hd_decap_3
XFILLER_26_184 vpwr vgnd scs8hd_fill_2
XFILLER_26_173 vgnd vpwr scs8hd_decap_8
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_fill_1
XFILLER_18_107 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_110 vgnd vpwr scs8hd_decap_12
XFILLER_23_154 vgnd vpwr scs8hd_decap_12
XFILLER_11_32 vgnd vpwr scs8hd_decap_12
X_35_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_20_168 vgnd vpwr scs8hd_decap_12
XFILLER_7_117 vgnd vpwr scs8hd_decap_12
XFILLER_22_86 vgnd vpwr scs8hd_decap_12
XFILLER_19_202 vpwr vgnd scs8hd_fill_2
X_18_ chanx_right_in[18] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_25_227 vgnd vpwr scs8hd_decap_12
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_293 vgnd vpwr scs8hd_decap_6
XFILLER_30_296 vgnd vpwr scs8hd_decap_3
XFILLER_30_252 vgnd vpwr scs8hd_decap_8
XFILLER_22_208 vgnd vpwr scs8hd_decap_12
XFILLER_12_7 vgnd vpwr scs8hd_decap_12
XFILLER_28_74 vgnd vpwr scs8hd_decap_12
XFILLER_21_296 vgnd vpwr scs8hd_decap_3
XFILLER_21_274 vgnd vpwr scs8hd_fill_1
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_12_296 vgnd vpwr scs8hd_decap_3
XFILLER_12_252 vgnd vpwr scs8hd_decap_12
XFILLER_8_245 vgnd vpwr scs8hd_decap_3
XFILLER_14_76 vpwr vgnd scs8hd_fill_2
XFILLER_14_43 vgnd vpwr scs8hd_decap_12
XFILLER_5_215 vgnd vpwr scs8hd_decap_12
XFILLER_4_281 vgnd vpwr scs8hd_decap_12
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_fill_1
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_141 vgnd vpwr scs8hd_decap_12
XFILLER_23_166 vgnd vpwr scs8hd_decap_12
XFILLER_11_44 vgnd vpwr scs8hd_decap_12
X_34_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_9_192 vpwr vgnd scs8hd_fill_2
XFILLER_22_98 vgnd vpwr scs8hd_decap_12
XFILLER_7_129 vgnd vpwr scs8hd_decap_12
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
X_17_ chanx_right_in[19] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_25_239 vgnd vpwr scs8hd_decap_8
XFILLER_6_184 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_76 vpwr vgnd scs8hd_fill_2
XFILLER_17_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_154 vgnd vpwr scs8hd_decap_3
XFILLER_30_264 vgnd vpwr scs8hd_decap_12
XFILLER_15_250 vgnd vpwr scs8hd_decap_12
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.scs8hd_buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X top_grid_pin_0_
+ vgnd vpwr scs8hd_buf_1
XFILLER_28_86 vgnd vpwr scs8hd_decap_12
XFILLER_12_264 vgnd vpwr scs8hd_decap_12
XFILLER_12_220 vgnd vpwr scs8hd_decap_12
XFILLER_14_55 vgnd vpwr scs8hd_decap_6
XFILLER_5_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_293 vgnd vpwr scs8hd_decap_6
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_32 vgnd vpwr scs8hd_decap_12
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_208 vgnd vpwr scs8hd_decap_12
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XFILLER_32_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_296 vgnd vpwr scs8hd_decap_3
XFILLER_1_274 vgnd vpwr scs8hd_fill_1
XFILLER_1_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_178 vgnd vpwr scs8hd_decap_12
XFILLER_11_56 vgnd vpwr scs8hd_decap_12
X_33_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_123 vgnd vpwr scs8hd_decap_12
XFILLER_33_251 vgnd vpwr scs8hd_decap_12
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_281 vgnd vpwr scs8hd_decap_12
X_16_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_196 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_32 vgnd vpwr scs8hd_decap_12
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_11 vgnd vpwr scs8hd_decap_12
XFILLER_30_276 vgnd vpwr scs8hd_decap_12
XFILLER_30_243 vgnd vpwr scs8hd_fill_1
XFILLER_15_262 vgnd vpwr scs8hd_decap_12
XFILLER_21_276 vgnd vpwr scs8hd_decap_12
XFILLER_28_98 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_decap_12
XFILLER_12_232 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_5_36 vgnd vpwr scs8hd_decap_12
XFILLER_29_162 vgnd vpwr scs8hd_decap_12
XANTENNA__03__A chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_5_239 vgnd vpwr scs8hd_decap_8
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_110 vgnd vpwr scs8hd_decap_12
XFILLER_25_44 vgnd vpwr scs8hd_decap_12
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XFILLER_32_135 vgnd vpwr scs8hd_decap_12
XFILLER_17_154 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S mux_bottom_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_68 vgnd vpwr scs8hd_decap_12
X_32_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_13_190 vgnd vpwr scs8hd_decap_12
XFILLER_9_150 vgnd vpwr scs8hd_decap_3
XANTENNA__11__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_11_105 vgnd vpwr scs8hd_decap_12
XFILLER_3_80 vgnd vpwr scs8hd_decap_12
XFILLER_34_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_171 vgnd vpwr scs8hd_decap_12
X_15_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_33_296 vgnd vpwr scs8hd_decap_3
XFILLER_33_263 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_293 vgnd vpwr scs8hd_decap_6
XFILLER_17_56 vgnd vpwr scs8hd_decap_12
XFILLER_17_23 vgnd vpwr scs8hd_decap_8
XFILLER_16_208 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_44 vgnd vpwr scs8hd_decap_12
XFILLER_15_296 vgnd vpwr scs8hd_decap_3
XFILLER_15_274 vgnd vpwr scs8hd_fill_1
XANTENNA__06__A chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_30_288 vgnd vpwr scs8hd_decap_8
XFILLER_21_288 vgnd vpwr scs8hd_decap_8
XFILLER_12_288 vgnd vpwr scs8hd_decap_8
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_48 vgnd vpwr scs8hd_decap_12
XFILLER_29_174 vgnd vpwr scs8hd_decap_12
XFILLER_29_141 vgnd vpwr scs8hd_decap_12
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XFILLER_32_147 vgnd vpwr scs8hd_decap_12
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_188 vgnd vpwr scs8hd_decap_12
XFILLER_25_56 vgnd vpwr scs8hd_decap_6
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_17_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_133 vpwr vgnd scs8hd_fill_2
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_12
XFILLER_1_276 vgnd vpwr scs8hd_decap_12
XANTENNA__14__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A mux_bottom_ipin_0.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_147 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_31_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_11_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_250 vgnd vpwr scs8hd_decap_12
XFILLER_19_206 vgnd vpwr scs8hd_decap_8
XFILLER_6_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_132 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_59 vpwr vgnd scs8hd_fill_2
X_14_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_56 vgnd vpwr scs8hd_decap_12
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_220 vgnd vpwr scs8hd_decap_12
XANTENNA__22__A chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_17_68 vgnd vpwr scs8hd_decap_6
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_245 vgnd vpwr scs8hd_decap_3
XFILLER_21_201 vpwr vgnd scs8hd_fill_2
XANTENNA__17__A chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_12_245 vgnd vpwr scs8hd_decap_3
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_9_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_186 vgnd vpwr scs8hd_decap_12
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_26_123 vgnd vpwr scs8hd_decap_6
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_2_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_288 vgnd vpwr scs8hd_decap_8
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__30__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_159 vgnd vpwr scs8hd_decap_12
XFILLER_17_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_159 vgnd vpwr scs8hd_decap_12
XFILLER_14_104 vgnd vpwr scs8hd_decap_12
XANTENNA__25__A chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_22_192 vpwr vgnd scs8hd_fill_2
X_30_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_11_129 vgnd vpwr scs8hd_decap_12
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_93 vgnd vpwr scs8hd_decap_12
XFILLER_27_262 vgnd vpwr scs8hd_decap_12
XFILLER_19_218 vgnd vpwr scs8hd_decap_12
XFILLER_10_184 vgnd vpwr scs8hd_decap_12
XFILLER_0_7 vpwr vgnd scs8hd_fill_2
XFILLER_6_144 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_12
XFILLER_33_276 vgnd vpwr scs8hd_decap_12
X_13_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_68 vgnd vpwr scs8hd_decap_12
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_232 vgnd vpwr scs8hd_decap_12
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S mux_bottom_ipin_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_276 vgnd vpwr scs8hd_decap_12
XFILLER_21_213 vgnd vpwr scs8hd_fill_1
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XANTENNA__33__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_7_250 vgnd vpwr scs8hd_decap_12
XFILLER_29_198 vgnd vpwr scs8hd_decap_12
XFILLER_29_154 vpwr vgnd scs8hd_fill_2
XANTENNA__28__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XFILLER_1_256 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_fill_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_25_190 vgnd vpwr scs8hd_decap_12
XFILLER_15_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D mux_bottom_ipin_0.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_105 vgnd vpwr scs8hd_decap_12
XFILLER_22_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S mux_bottom_ipin_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__41__A chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_14_116 vgnd vpwr scs8hd_decap_6
XFILLER_28_208 vgnd vpwr scs8hd_decap_12
XFILLER_9_186 vpwr vgnd scs8hd_fill_2
XFILLER_27_296 vgnd vpwr scs8hd_decap_3
XFILLER_27_274 vgnd vpwr scs8hd_fill_1
XFILLER_22_59 vpwr vgnd scs8hd_fill_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__36__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_288 vgnd vpwr scs8hd_decap_8
XFILLER_10_196 vgnd vpwr scs8hd_decap_12
X_12_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_123 vgnd vpwr scs8hd_decap_4
XFILLER_6_156 vgnd vpwr scs8hd_decap_12
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_23_80 vgnd vpwr scs8hd_decap_12
XFILLER_15_288 vgnd vpwr scs8hd_decap_8
XFILLER_21_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_9_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_262 vgnd vpwr scs8hd_decap_12
XFILLER_30_59 vpwr vgnd scs8hd_fill_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XFILLER_31_80 vgnd vpwr scs8hd_decap_12
XANTENNA__39__A chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_15_70 vpwr vgnd scs8hd_fill_2
XFILLER_1_268 vgnd vpwr scs8hd_decap_6
XFILLER_1_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_117 vgnd vpwr scs8hd_decap_12
XFILLER_9_154 vgnd vpwr scs8hd_decap_12
XFILLER_22_27 vgnd vpwr scs8hd_decap_12
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
X_11_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_18_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_168 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_190 vgnd vpwr scs8hd_decap_12
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_2_171 vgnd vpwr scs8hd_decap_12
XFILLER_28_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_281 vgnd vpwr scs8hd_decap_12
XFILLER_8_208 vgnd vpwr scs8hd_decap_12
XFILLER_7_274 vgnd vpwr scs8hd_fill_1
XFILLER_7_296 vgnd vpwr scs8hd_decap_3
XFILLER_30_27 vgnd vpwr scs8hd_decap_12
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XFILLER_29_91 vgnd vpwr scs8hd_fill_1
XFILLER_29_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_4
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_6_62 vgnd vpwr scs8hd_decap_12
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_17_137 vpwr vgnd scs8hd_fill_2
XFILLER_15_93 vgnd vpwr scs8hd_decap_12
XFILLER_23_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_280 vgnd vpwr scs8hd_decap_12
XFILLER_22_184 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0 mux_bottom_ipin_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_166 vgnd vpwr scs8hd_decap_12
XFILLER_22_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_276 vgnd vpwr scs8hd_decap_12
XFILLER_18_232 vgnd vpwr scs8hd_decap_12
XFILLER_10_110 vgnd vpwr scs8hd_decap_12
X_10_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_257 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S mux_bottom_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_117 vgnd vpwr scs8hd_decap_12
XFILLER_23_93 vgnd vpwr scs8hd_decap_12
XFILLER_21_227 vgnd vpwr scs8hd_decap_12
XFILLER_21_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_28_27 vgnd vpwr scs8hd_decap_12
XFILLER_20_293 vgnd vpwr scs8hd_decap_6
XFILLER_30_39 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1 mux_bottom_ipin_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_245 vgnd vpwr scs8hd_decap_12
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XFILLER_26_149 vgnd vpwr scs8hd_decap_12
XFILLER_19_190 vgnd vpwr scs8hd_decap_6
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_6_74 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XFILLER_34_171 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_17_105 vgnd vpwr scs8hd_decap_12
XFILLER_1_215 vgnd vpwr scs8hd_decap_12
XFILLER_31_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_93 vgnd vpwr scs8hd_decap_12
XFILLER_16_171 vgnd vpwr scs8hd_decap_12
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XFILLER_0_292 vgnd vpwr scs8hd_decap_6
XFILLER_22_196 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1 mux_bottom_ipin_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_19 vgnd vpwr scs8hd_decap_12
XFILLER_13_141 vgnd vpwr scs8hd_decap_12
XFILLER_9_178 vgnd vpwr scs8hd_decap_8
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_27_288 vgnd vpwr scs8hd_decap_8
XFILLER_12_62 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_269 vgnd vpwr scs8hd_decap_12
XFILLER_3_129 vgnd vpwr scs8hd_decap_12
XFILLER_30_239 vgnd vpwr scs8hd_decap_4
XFILLER_15_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_184 vgnd vpwr scs8hd_decap_12
XFILLER_28_39 vgnd vpwr scs8hd_decap_12
XFILLER_21_239 vgnd vpwr scs8hd_decap_8
XFILLER_18_83 vgnd vpwr scs8hd_decap_12
XFILLER_14_19 vgnd vpwr scs8hd_decap_12
XFILLER_7_276 vgnd vpwr scs8hd_decap_12
XFILLER_29_158 vpwr vgnd scs8hd_fill_2
XFILLER_20_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_117 vgnd vpwr scs8hd_fill_1
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_1_227 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_3_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_74 vgnd vpwr scs8hd_decap_12
XFILLER_10_123 vgnd vpwr scs8hd_decap_12
XFILLER_6_127 vgnd vpwr scs8hd_fill_1
XFILLER_33_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_281 vgnd vpwr scs8hd_decap_12
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_15_215 vgnd vpwr scs8hd_decap_12
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_11 vgnd vpwr scs8hd_decap_12
XFILLER_2_196 vgnd vpwr scs8hd_decap_12
XFILLER_14_281 vgnd vpwr scs8hd_decap_12
XFILLER_18_95 vgnd vpwr scs8hd_decap_12
XFILLER_18_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_288 vgnd vpwr scs8hd_decap_8
XFILLER_4_214 vgnd vpwr scs8hd_decap_12
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_83 vpwr vgnd scs8hd_fill_2
XFILLER_20_74 vgnd vpwr scs8hd_decap_12
XFILLER_4_269 vgnd vpwr scs8hd_decap_12
XFILLER_6_98 vgnd vpwr scs8hd_decap_12
XFILLER_34_184 vgnd vpwr scs8hd_decap_12
XFILLER_26_129 vgnd vpwr scs8hd_fill_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_1_239 vgnd vpwr scs8hd_decap_6
XFILLER_17_129 vpwr vgnd scs8hd_fill_2
XFILLER_31_154 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_184 vgnd vpwr scs8hd_decap_12
XFILLER_26_62 vgnd vpwr scs8hd_decap_12
XFILLER_26_51 vgnd vpwr scs8hd_decap_8
XFILLER_22_110 vgnd vpwr scs8hd_decap_12
XFILLER_13_154 vgnd vpwr scs8hd_decap_12
XFILLER_3_44 vgnd vpwr scs8hd_decap_12
XFILLER_27_213 vgnd vpwr scs8hd_fill_1
XFILLER_10_135 vgnd vpwr scs8hd_decap_12
XFILLER_33_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_86 vgnd vpwr scs8hd_decap_12
XFILLER_12_31 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_293 vgnd vpwr scs8hd_decap_6
XFILLER_30_208 vgnd vpwr scs8hd_decap_4
XFILLER_15_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_293 vgnd vpwr scs8hd_decap_6
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_0_23 vgnd vpwr scs8hd_decap_8
XFILLER_9_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_241 vgnd vpwr scs8hd_decap_3
XFILLER_12_208 vgnd vpwr scs8hd_decap_12
XFILLER_34_62 vgnd vpwr scs8hd_decap_12
XFILLER_34_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_296 vgnd vpwr scs8hd_decap_3
XFILLER_11_274 vgnd vpwr scs8hd_fill_1
XFILLER_11_252 vpwr vgnd scs8hd_fill_2
XFILLER_29_105 vgnd vpwr scs8hd_decap_12
XFILLER_28_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_86 vgnd vpwr scs8hd_decap_12
XFILLER_20_31 vgnd vpwr scs8hd_decap_12
XFILLER_4_226 vgnd vpwr scs8hd_decap_12
XFILLER_34_196 vgnd vpwr scs8hd_decap_12
XFILLER_25_152 vgnd vpwr scs8hd_fill_1
XFILLER_31_166 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_196 vgnd vpwr scs8hd_decap_12
.ends

